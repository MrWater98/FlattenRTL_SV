module RocketTile (
  input cov_store,
  input clock,
  input reset,
  output auto_broadcast_out_0_valid,
  output [39:0] auto_broadcast_out_0_iaddr,
  output [31:0] auto_broadcast_out_0_insn,
  output [2:0] auto_broadcast_out_0_priv,
  output auto_broadcast_out_0_exception,
  output auto_broadcast_out_0_interrupt,
  output [63:0] auto_broadcast_out_0_cause,
  output [39:0] auto_broadcast_out_0_tval,
  output auto_wfi_out_0,
  output auto_cease_out_0,
  output auto_halt_out_0,
  input auto_int_in_xing_in_2_sync_0,
  input auto_int_in_xing_in_1_sync_0,
  input auto_int_in_xing_in_0_sync_0,
  input auto_int_in_xing_in_0_sync_1,
  input auto_intsink_in_sync_0,
  output auto_trace_core_source_out_group_0_iretire,
  output [31:0] auto_trace_core_source_out_group_0_iaddr,
  output [3:0] auto_trace_core_source_out_group_0_itype,
  output auto_trace_core_source_out_group_0_ilastsize,
  output [3:0] auto_trace_core_source_out_priv,
  output [31:0] auto_trace_core_source_out_tval,
  output [31:0] auto_trace_core_source_out_cause,
  input auto_nmi_in_rnmi,
  input [31:0] auto_nmi_in_rnmi_interrupt_vector,
  input [31:0] auto_nmi_in_rnmi_exception_vector,
  input auto_nmi_in_unmi,
  input [31:0] auto_nmi_in_unmi_interrupt_vector,
  input [31:0] auto_nmi_in_unmi_exception_vector,
  input [31:0] auto_reset_vector_in,
  input auto_hartid_in,
  input auto_tl_master_xing_out_a_ready,
  output auto_tl_master_xing_out_a_valid,
  output [2:0] auto_tl_master_xing_out_a_bits_opcode,
  output [2:0] auto_tl_master_xing_out_a_bits_param,
  output [3:0] auto_tl_master_xing_out_a_bits_size,
  output [1:0] auto_tl_master_xing_out_a_bits_source,
  output [31:0] auto_tl_master_xing_out_a_bits_address,
  output [7:0] auto_tl_master_xing_out_a_bits_mask,
  output [63:0] auto_tl_master_xing_out_a_bits_data,
  output auto_tl_master_xing_out_a_bits_corrupt,
  output auto_tl_master_xing_out_b_ready,
  input auto_tl_master_xing_out_b_valid,
  input [2:0] auto_tl_master_xing_out_b_bits_opcode,
  input [1:0] auto_tl_master_xing_out_b_bits_param,
  input [3:0] auto_tl_master_xing_out_b_bits_size,
  input [1:0] auto_tl_master_xing_out_b_bits_source,
  input [31:0] auto_tl_master_xing_out_b_bits_address,
  input [7:0] auto_tl_master_xing_out_b_bits_mask,
  input [63:0] auto_tl_master_xing_out_b_bits_data,
  input auto_tl_master_xing_out_b_bits_corrupt,
  input auto_tl_master_xing_out_c_ready,
  output auto_tl_master_xing_out_c_valid,
  output [2:0] auto_tl_master_xing_out_c_bits_opcode,
  output [2:0] auto_tl_master_xing_out_c_bits_param,
  output [3:0] auto_tl_master_xing_out_c_bits_size,
  output [1:0] auto_tl_master_xing_out_c_bits_source,
  output [31:0] auto_tl_master_xing_out_c_bits_address,
  output [63:0] auto_tl_master_xing_out_c_bits_data,
  output auto_tl_master_xing_out_c_bits_corrupt,
  output auto_tl_master_xing_out_d_ready,
  input auto_tl_master_xing_out_d_valid,
  input [2:0] auto_tl_master_xing_out_d_bits_opcode,
  input [1:0] auto_tl_master_xing_out_d_bits_param,
  input [3:0] auto_tl_master_xing_out_d_bits_size,
  input [1:0] auto_tl_master_xing_out_d_bits_source,
  input [1:0] auto_tl_master_xing_out_d_bits_sink,
  input auto_tl_master_xing_out_d_bits_denied,
  input [63:0] auto_tl_master_xing_out_d_bits_data,
  input auto_tl_master_xing_out_d_bits_corrupt,
  input auto_tl_master_xing_out_e_ready,
  output auto_tl_master_xing_out_e_valid,
  output [1:0] auto_tl_master_xing_out_e_bits_sink,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input tlMasterXbar_halt,
  input intXbar_halt,
  input fpuOpt_halt,
  input dcacheArb_halt,
  input frontend_halt,
  input dcache_halt,
  input broadcast_3_halt,
  input core_halt,
  input broadcast_halt,
  input broadcast_1_halt,
  input ptw_halt,
  input eos,
  input cov_sr,
  output reg  eos_hs,
  output reg  cmt_instr) ; 
   reg debug_print ;  
   reg trace_en ;  
   integer fd ;  
   integer iteration ;  
   wire [63:0] mstatus_wire ;  
   wire tlMasterXbar_clock ;  
   wire tlMasterXbar_reset ;  
   wire tlMasterXbar_auto_in_1_a_ready ;  
   wire tlMasterXbar_auto_in_1_a_valid ;  
   wire [31:0] tlMasterXbar_auto_in_1_a_bits_address ;  
   wire tlMasterXbar_auto_in_1_d_valid ;  
   wire [2:0] tlMasterXbar_auto_in_1_d_bits_opcode ;  
   wire [3:0] tlMasterXbar_auto_in_1_d_bits_size ;  
   wire [63:0] tlMasterXbar_auto_in_1_d_bits_data ;  
   wire tlMasterXbar_auto_in_1_d_bits_corrupt ;  
   wire tlMasterXbar_auto_in_0_a_ready ;  
   wire tlMasterXbar_auto_in_0_a_valid ;  
   wire [2:0] tlMasterXbar_auto_in_0_a_bits_opcode ;  
   wire [2:0] tlMasterXbar_auto_in_0_a_bits_param ;  
   wire [3:0] tlMasterXbar_auto_in_0_a_bits_size ;  
   wire tlMasterXbar_auto_in_0_a_bits_source ;  
   wire [31:0] tlMasterXbar_auto_in_0_a_bits_address ;  
   wire [7:0] tlMasterXbar_auto_in_0_a_bits_mask ;  
   wire [63:0] tlMasterXbar_auto_in_0_a_bits_data ;  
   wire tlMasterXbar_auto_in_0_b_ready ;  
   wire tlMasterXbar_auto_in_0_b_valid ;  
   wire [1:0] tlMasterXbar_auto_in_0_b_bits_param ;  
   wire [3:0] tlMasterXbar_auto_in_0_b_bits_size ;  
   wire tlMasterXbar_auto_in_0_b_bits_source ;  
   wire [31:0] tlMasterXbar_auto_in_0_b_bits_address ;  
   wire tlMasterXbar_auto_in_0_c_ready ;  
   wire tlMasterXbar_auto_in_0_c_valid ;  
   wire [2:0] tlMasterXbar_auto_in_0_c_bits_opcode ;  
   wire [2:0] tlMasterXbar_auto_in_0_c_bits_param ;  
   wire [3:0] tlMasterXbar_auto_in_0_c_bits_size ;  
   wire tlMasterXbar_auto_in_0_c_bits_source ;  
   wire [31:0] tlMasterXbar_auto_in_0_c_bits_address ;  
   wire [63:0] tlMasterXbar_auto_in_0_c_bits_data ;  
   wire tlMasterXbar_auto_in_0_d_ready ;  
   wire tlMasterXbar_auto_in_0_d_valid ;  
   wire [2:0] tlMasterXbar_auto_in_0_d_bits_opcode ;  
   wire [1:0] tlMasterXbar_auto_in_0_d_bits_param ;  
   wire [3:0] tlMasterXbar_auto_in_0_d_bits_size ;  
   wire tlMasterXbar_auto_in_0_d_bits_source ;  
   wire [1:0] tlMasterXbar_auto_in_0_d_bits_sink ;  
   wire tlMasterXbar_auto_in_0_d_bits_denied ;  
   wire [63:0] tlMasterXbar_auto_in_0_d_bits_data ;  
   wire tlMasterXbar_auto_in_0_e_ready ;  
   wire tlMasterXbar_auto_in_0_e_valid ;  
   wire [1:0] tlMasterXbar_auto_in_0_e_bits_sink ;  
   wire tlMasterXbar_auto_out_a_ready ;  
   wire tlMasterXbar_auto_out_a_valid ;  
   wire [2:0] tlMasterXbar_auto_out_a_bits_opcode ;  
   wire [2:0] tlMasterXbar_auto_out_a_bits_param ;  
   wire [3:0] tlMasterXbar_auto_out_a_bits_size ;  
   wire [1:0] tlMasterXbar_auto_out_a_bits_source ;  
   wire [31:0] tlMasterXbar_auto_out_a_bits_address ;  
   wire [7:0] tlMasterXbar_auto_out_a_bits_mask ;  
   wire [63:0] tlMasterXbar_auto_out_a_bits_data ;  
   wire tlMasterXbar_auto_out_b_ready ;  
   wire tlMasterXbar_auto_out_b_valid ;  
   wire [2:0] tlMasterXbar_auto_out_b_bits_opcode ;  
   wire [1:0] tlMasterXbar_auto_out_b_bits_param ;  
   wire [3:0] tlMasterXbar_auto_out_b_bits_size ;  
   wire [1:0] tlMasterXbar_auto_out_b_bits_source ;  
   wire [31:0] tlMasterXbar_auto_out_b_bits_address ;  
   wire [7:0] tlMasterXbar_auto_out_b_bits_mask ;  
   wire tlMasterXbar_auto_out_b_bits_corrupt ;  
   wire tlMasterXbar_auto_out_c_ready ;  
   wire tlMasterXbar_auto_out_c_valid ;  
   wire [2:0] tlMasterXbar_auto_out_c_bits_opcode ;  
   wire [2:0] tlMasterXbar_auto_out_c_bits_param ;  
   wire [3:0] tlMasterXbar_auto_out_c_bits_size ;  
   wire [1:0] tlMasterXbar_auto_out_c_bits_source ;  
   wire [31:0] tlMasterXbar_auto_out_c_bits_address ;  
   wire [63:0] tlMasterXbar_auto_out_c_bits_data ;  
   wire tlMasterXbar_auto_out_d_ready ;  
   wire tlMasterXbar_auto_out_d_valid ;  
   wire [2:0] tlMasterXbar_auto_out_d_bits_opcode ;  
   wire [1:0] tlMasterXbar_auto_out_d_bits_param ;  
   wire [3:0] tlMasterXbar_auto_out_d_bits_size ;  
   wire [1:0] tlMasterXbar_auto_out_d_bits_source ;  
   wire [1:0] tlMasterXbar_auto_out_d_bits_sink ;  
   wire tlMasterXbar_auto_out_d_bits_denied ;  
   wire [63:0] tlMasterXbar_auto_out_d_bits_data ;  
   wire tlMasterXbar_auto_out_d_bits_corrupt ;  
   wire tlMasterXbar_auto_out_e_ready ;  
   wire tlMasterXbar_auto_out_e_valid ;  
   wire [1:0] tlMasterXbar_auto_out_e_bits_sink ;  
   wire [29:0] tlMasterXbar_io_covSum ;  
   wire tlMasterXbar_metaAssert ;  
   wire tlMasterXbar_metaReset ;  
   wire tlMasterXbar_monitor_halt ;  
   wire tlMasterXbar_monitor_1_halt ;  
   wire intXbar_auto_int_in_3_0 ;  
   wire intXbar_auto_int_in_2_0 ;  
   wire intXbar_auto_int_in_1_0 ;  
   wire intXbar_auto_int_in_1_1 ;  
   wire intXbar_auto_int_in_0_0 ;  
   wire intXbar_auto_int_out_0 ;  
   wire intXbar_auto_int_out_1 ;  
   wire intXbar_auto_int_out_2 ;  
   wire intXbar_auto_int_out_3 ;  
   wire intXbar_auto_int_out_4 ;  
   wire [29:0] intXbar_io_covSum ;  
   wire intXbar_metaAssert ;  
   wire broadcast_auto_in ;  
   wire broadcast_auto_out ;  
   wire [29:0] broadcast_io_covSum ;  
   wire broadcast_metaAssert ;  
   wire [31:0] broadcast_1_auto_in ;  
   wire [31:0] broadcast_1_auto_out_1 ;  
   wire [29:0] broadcast_1_io_covSum ;  
   wire broadcast_1_metaAssert ;  
   wire broadcast_3_auto_in_0_valid ;  
   wire [39:0] broadcast_3_auto_in_0_iaddr ;  
   wire [31:0] broadcast_3_auto_in_0_insn ;  
   wire [2:0] broadcast_3_auto_in_0_priv ;  
   wire broadcast_3_auto_in_0_exception ;  
   wire broadcast_3_auto_in_0_interrupt ;  
   wire [63:0] broadcast_3_auto_in_0_cause ;  
   wire [39:0] broadcast_3_auto_in_0_tval ;  
   wire broadcast_3_auto_out_0_valid ;  
   wire [39:0] broadcast_3_auto_out_0_iaddr ;  
   wire [31:0] broadcast_3_auto_out_0_insn ;  
   wire [2:0] broadcast_3_auto_out_0_priv ;  
   wire broadcast_3_auto_out_0_exception ;  
   wire broadcast_3_auto_out_0_interrupt ;  
   wire [63:0] broadcast_3_auto_out_0_cause ;  
   wire [39:0] broadcast_3_auto_out_0_tval ;  
   wire [29:0] broadcast_3_io_covSum ;  
   wire broadcast_3_metaAssert ;  
   wire dcache_gated_clock ;  
   wire dcache_reset ;  
   wire dcache_auto_out_a_ready ;  
   wire dcache_auto_out_a_valid ;  
   wire [2:0] dcache_auto_out_a_bits_opcode ;  
   wire [2:0] dcache_auto_out_a_bits_param ;  
   wire [3:0] dcache_auto_out_a_bits_size ;  
   wire dcache_auto_out_a_bits_source ;  
   wire [31:0] dcache_auto_out_a_bits_address ;  
   wire [7:0] dcache_auto_out_a_bits_mask ;  
   wire [63:0] dcache_auto_out_a_bits_data ;  
   wire dcache_auto_out_b_ready ;  
   wire dcache_auto_out_b_valid ;  
   wire [1:0] dcache_auto_out_b_bits_param ;  
   wire [3:0] dcache_auto_out_b_bits_size ;  
   wire dcache_auto_out_b_bits_source ;  
   wire [31:0] dcache_auto_out_b_bits_address ;  
   wire dcache_auto_out_c_ready ;  
   wire dcache_auto_out_c_valid ;  
   wire [2:0] dcache_auto_out_c_bits_opcode ;  
   wire [2:0] dcache_auto_out_c_bits_param ;  
   wire [3:0] dcache_auto_out_c_bits_size ;  
   wire dcache_auto_out_c_bits_source ;  
   wire [31:0] dcache_auto_out_c_bits_address ;  
   wire [63:0] dcache_auto_out_c_bits_data ;  
   wire dcache_auto_out_d_ready ;  
   wire dcache_auto_out_d_valid ;  
   wire [2:0] dcache_auto_out_d_bits_opcode ;  
   wire [1:0] dcache_auto_out_d_bits_param ;  
   wire [3:0] dcache_auto_out_d_bits_size ;  
   wire dcache_auto_out_d_bits_source ;  
   wire [1:0] dcache_auto_out_d_bits_sink ;  
   wire dcache_auto_out_d_bits_denied ;  
   wire [63:0] dcache_auto_out_d_bits_data ;  
   wire dcache_auto_out_e_ready ;  
   wire dcache_auto_out_e_valid ;  
   wire [1:0] dcache_auto_out_e_bits_sink ;  
   wire dcache_io_cpu_req_ready ;  
   wire dcache_io_cpu_req_valid ;  
   wire [39:0] dcache_io_cpu_req_bits_addr ;  
   wire [6:0] dcache_io_cpu_req_bits_tag ;  
   wire [4:0] dcache_io_cpu_req_bits_cmd ;  
   wire [1:0] dcache_io_cpu_req_bits_size ;  
   wire dcache_io_cpu_req_bits_signed ;  
   wire dcache_io_cpu_req_bits_phys ;  
   wire dcache_io_cpu_s1_kill ;  
   wire [63:0] dcache_io_cpu_s1_data_data ;  
   wire dcache_io_cpu_s2_nack ;  
   wire dcache_io_cpu_resp_valid ;  
   wire [6:0] dcache_io_cpu_resp_bits_tag ;  
   wire [1:0] dcache_io_cpu_resp_bits_size ;  
   wire [63:0] dcache_io_cpu_resp_bits_data ;  
   wire dcache_io_cpu_resp_bits_replay ;  
   wire dcache_io_cpu_resp_bits_has_data ;  
   wire [63:0] dcache_io_cpu_resp_bits_data_word_bypass ;  
   wire dcache_io_cpu_replay_next ;  
   wire dcache_io_cpu_s2_xcpt_ma_ld ;  
   wire dcache_io_cpu_s2_xcpt_ma_st ;  
   wire dcache_io_cpu_s2_xcpt_pf_ld ;  
   wire dcache_io_cpu_s2_xcpt_pf_st ;  
   wire dcache_io_cpu_s2_xcpt_ae_ld ;  
   wire dcache_io_cpu_s2_xcpt_ae_st ;  
   wire dcache_io_cpu_ordered ;  
   wire dcache_io_cpu_perf_release ;  
   wire dcache_io_cpu_perf_grant ;  
   wire dcache_io_ptw_req_ready ;  
   wire dcache_io_ptw_req_valid ;  
   wire [26:0] dcache_io_ptw_req_bits_bits_addr ;  
   wire dcache_io_ptw_resp_valid ;  
   wire dcache_io_ptw_resp_bits_ae ;  
   wire [53:0] dcache_io_ptw_resp_bits_pte_ppn ;  
   wire dcache_io_ptw_resp_bits_pte_d ;  
   wire dcache_io_ptw_resp_bits_pte_a ;  
   wire dcache_io_ptw_resp_bits_pte_g ;  
   wire dcache_io_ptw_resp_bits_pte_u ;  
   wire dcache_io_ptw_resp_bits_pte_x ;  
   wire dcache_io_ptw_resp_bits_pte_w ;  
   wire dcache_io_ptw_resp_bits_pte_r ;  
   wire dcache_io_ptw_resp_bits_pte_v ;  
   wire [1:0] dcache_io_ptw_resp_bits_level ;  
   wire dcache_io_ptw_resp_bits_homogeneous ;  
   wire [3:0] dcache_io_ptw_ptbr_mode ;  
   wire dcache_io_ptw_status_debug ;  
   wire [1:0] dcache_io_ptw_status_dprv ;  
   wire dcache_io_ptw_status_mxr ;  
   wire dcache_io_ptw_status_sum ;  
   wire dcache_io_ptw_pmp_0_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_0_cfg_a ;  
   wire dcache_io_ptw_pmp_0_cfg_x ;  
   wire dcache_io_ptw_pmp_0_cfg_w ;  
   wire dcache_io_ptw_pmp_0_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_0_addr ;  
   wire [31:0] dcache_io_ptw_pmp_0_mask ;  
   wire dcache_io_ptw_pmp_1_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_1_cfg_a ;  
   wire dcache_io_ptw_pmp_1_cfg_x ;  
   wire dcache_io_ptw_pmp_1_cfg_w ;  
   wire dcache_io_ptw_pmp_1_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_1_addr ;  
   wire [31:0] dcache_io_ptw_pmp_1_mask ;  
   wire dcache_io_ptw_pmp_2_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_2_cfg_a ;  
   wire dcache_io_ptw_pmp_2_cfg_x ;  
   wire dcache_io_ptw_pmp_2_cfg_w ;  
   wire dcache_io_ptw_pmp_2_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_2_addr ;  
   wire [31:0] dcache_io_ptw_pmp_2_mask ;  
   wire dcache_io_ptw_pmp_3_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_3_cfg_a ;  
   wire dcache_io_ptw_pmp_3_cfg_x ;  
   wire dcache_io_ptw_pmp_3_cfg_w ;  
   wire dcache_io_ptw_pmp_3_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_3_addr ;  
   wire [31:0] dcache_io_ptw_pmp_3_mask ;  
   wire dcache_io_ptw_pmp_4_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_4_cfg_a ;  
   wire dcache_io_ptw_pmp_4_cfg_x ;  
   wire dcache_io_ptw_pmp_4_cfg_w ;  
   wire dcache_io_ptw_pmp_4_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_4_addr ;  
   wire [31:0] dcache_io_ptw_pmp_4_mask ;  
   wire dcache_io_ptw_pmp_5_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_5_cfg_a ;  
   wire dcache_io_ptw_pmp_5_cfg_x ;  
   wire dcache_io_ptw_pmp_5_cfg_w ;  
   wire dcache_io_ptw_pmp_5_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_5_addr ;  
   wire [31:0] dcache_io_ptw_pmp_5_mask ;  
   wire dcache_io_ptw_pmp_6_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_6_cfg_a ;  
   wire dcache_io_ptw_pmp_6_cfg_x ;  
   wire dcache_io_ptw_pmp_6_cfg_w ;  
   wire dcache_io_ptw_pmp_6_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_6_addr ;  
   wire [31:0] dcache_io_ptw_pmp_6_mask ;  
   wire dcache_io_ptw_pmp_7_cfg_l ;  
   wire [1:0] dcache_io_ptw_pmp_7_cfg_a ;  
   wire dcache_io_ptw_pmp_7_cfg_x ;  
   wire dcache_io_ptw_pmp_7_cfg_w ;  
   wire dcache_io_ptw_pmp_7_cfg_r ;  
   wire [29:0] dcache_io_ptw_pmp_7_addr ;  
   wire [31:0] dcache_io_ptw_pmp_7_mask ;  
   wire [29:0] dcache_io_covSum ;  
   wire dcache_metaAssert ;  
   wire dcache_metaReset ;  
   wire dcache_data_halt ;  
   wire dcache_tlb_halt ;  
   wire dcache_pma_checker_halt ;  
   wire dcache_lfsr_prng_halt ;  
   wire frontend_gated_clock ;  
   wire frontend_reset ;  
   wire frontend_auto_icache_master_out_a_ready ;  
   wire frontend_auto_icache_master_out_a_valid ;  
   wire [31:0] frontend_auto_icache_master_out_a_bits_address ;  
   wire frontend_auto_icache_master_out_d_valid ;  
   wire [2:0] frontend_auto_icache_master_out_d_bits_opcode ;  
   wire [3:0] frontend_auto_icache_master_out_d_bits_size ;  
   wire [63:0] frontend_auto_icache_master_out_d_bits_data ;  
   wire frontend_auto_icache_master_out_d_bits_corrupt ;  
   wire [31:0] frontend_auto_reset_vector_sink_in ;  
   wire frontend_io_cpu_might_request ;  
   wire frontend_io_cpu_req_valid ;  
   wire [39:0] frontend_io_cpu_req_bits_pc ;  
   wire frontend_io_cpu_req_bits_speculative ;  
   wire frontend_io_cpu_sfence_valid ;  
   wire frontend_io_cpu_sfence_bits_rs1 ;  
   wire frontend_io_cpu_sfence_bits_rs2 ;  
   wire [38:0] frontend_io_cpu_sfence_bits_addr ;  
   wire frontend_io_cpu_resp_ready ;  
   wire frontend_io_cpu_resp_valid ;  
   wire frontend_io_cpu_resp_bits_btb_taken ;  
   wire frontend_io_cpu_resp_bits_btb_bridx ;  
   wire [4:0] frontend_io_cpu_resp_bits_btb_entry ;  
   wire [7:0] frontend_io_cpu_resp_bits_btb_bht_history ;  
   wire [39:0] frontend_io_cpu_resp_bits_pc ;  
   wire [31:0] frontend_io_cpu_resp_bits_data ;  
   wire frontend_io_cpu_resp_bits_xcpt_pf_inst ;  
   wire frontend_io_cpu_resp_bits_xcpt_ae_inst ;  
   wire frontend_io_cpu_resp_bits_replay ;  
   wire frontend_io_cpu_btb_update_valid ;  
   wire [4:0] frontend_io_cpu_btb_update_bits_prediction_entry ;  
   wire [38:0] frontend_io_cpu_btb_update_bits_pc ;  
   wire frontend_io_cpu_btb_update_bits_isValid ;  
   wire [38:0] frontend_io_cpu_btb_update_bits_br_pc ;  
   wire [1:0] frontend_io_cpu_btb_update_bits_cfiType ;  
   wire frontend_io_cpu_bht_update_valid ;  
   wire [7:0] frontend_io_cpu_bht_update_bits_prediction_history ;  
   wire [38:0] frontend_io_cpu_bht_update_bits_pc ;  
   wire frontend_io_cpu_bht_update_bits_branch ;  
   wire frontend_io_cpu_bht_update_bits_taken ;  
   wire frontend_io_cpu_bht_update_bits_mispredict ;  
   wire frontend_io_cpu_flush_icache ;  
   wire [39:0] frontend_io_cpu_npc ;  
   wire frontend_io_ptw_req_ready ;  
   wire frontend_io_ptw_req_valid ;  
   wire frontend_io_ptw_req_bits_valid ;  
   wire [26:0] frontend_io_ptw_req_bits_bits_addr ;  
   wire frontend_io_ptw_resp_valid ;  
   wire frontend_io_ptw_resp_bits_ae ;  
   wire [53:0] frontend_io_ptw_resp_bits_pte_ppn ;  
   wire frontend_io_ptw_resp_bits_pte_d ;  
   wire frontend_io_ptw_resp_bits_pte_a ;  
   wire frontend_io_ptw_resp_bits_pte_g ;  
   wire frontend_io_ptw_resp_bits_pte_u ;  
   wire frontend_io_ptw_resp_bits_pte_x ;  
   wire frontend_io_ptw_resp_bits_pte_w ;  
   wire frontend_io_ptw_resp_bits_pte_r ;  
   wire frontend_io_ptw_resp_bits_pte_v ;  
   wire [1:0] frontend_io_ptw_resp_bits_level ;  
   wire frontend_io_ptw_resp_bits_homogeneous ;  
   wire [3:0] frontend_io_ptw_ptbr_mode ;  
   wire frontend_io_ptw_status_debug ;  
   wire [1:0] frontend_io_ptw_status_prv ;  
   wire frontend_io_ptw_pmp_0_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_0_cfg_a ;  
   wire frontend_io_ptw_pmp_0_cfg_x ;  
   wire frontend_io_ptw_pmp_0_cfg_w ;  
   wire frontend_io_ptw_pmp_0_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_0_addr ;  
   wire [31:0] frontend_io_ptw_pmp_0_mask ;  
   wire frontend_io_ptw_pmp_1_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_1_cfg_a ;  
   wire frontend_io_ptw_pmp_1_cfg_x ;  
   wire frontend_io_ptw_pmp_1_cfg_w ;  
   wire frontend_io_ptw_pmp_1_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_1_addr ;  
   wire [31:0] frontend_io_ptw_pmp_1_mask ;  
   wire frontend_io_ptw_pmp_2_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_2_cfg_a ;  
   wire frontend_io_ptw_pmp_2_cfg_x ;  
   wire frontend_io_ptw_pmp_2_cfg_w ;  
   wire frontend_io_ptw_pmp_2_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_2_addr ;  
   wire [31:0] frontend_io_ptw_pmp_2_mask ;  
   wire frontend_io_ptw_pmp_3_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_3_cfg_a ;  
   wire frontend_io_ptw_pmp_3_cfg_x ;  
   wire frontend_io_ptw_pmp_3_cfg_w ;  
   wire frontend_io_ptw_pmp_3_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_3_addr ;  
   wire [31:0] frontend_io_ptw_pmp_3_mask ;  
   wire frontend_io_ptw_pmp_4_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_4_cfg_a ;  
   wire frontend_io_ptw_pmp_4_cfg_x ;  
   wire frontend_io_ptw_pmp_4_cfg_w ;  
   wire frontend_io_ptw_pmp_4_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_4_addr ;  
   wire [31:0] frontend_io_ptw_pmp_4_mask ;  
   wire frontend_io_ptw_pmp_5_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_5_cfg_a ;  
   wire frontend_io_ptw_pmp_5_cfg_x ;  
   wire frontend_io_ptw_pmp_5_cfg_w ;  
   wire frontend_io_ptw_pmp_5_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_5_addr ;  
   wire [31:0] frontend_io_ptw_pmp_5_mask ;  
   wire frontend_io_ptw_pmp_6_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_6_cfg_a ;  
   wire frontend_io_ptw_pmp_6_cfg_x ;  
   wire frontend_io_ptw_pmp_6_cfg_w ;  
   wire frontend_io_ptw_pmp_6_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_6_addr ;  
   wire [31:0] frontend_io_ptw_pmp_6_mask ;  
   wire frontend_io_ptw_pmp_7_cfg_l ;  
   wire [1:0] frontend_io_ptw_pmp_7_cfg_a ;  
   wire frontend_io_ptw_pmp_7_cfg_x ;  
   wire frontend_io_ptw_pmp_7_cfg_w ;  
   wire frontend_io_ptw_pmp_7_cfg_r ;  
   wire [29:0] frontend_io_ptw_pmp_7_addr ;  
   wire [31:0] frontend_io_ptw_pmp_7_mask ;  
   wire [63:0] frontend_io_ptw_customCSRs_csrs_0_value ;  
   wire [29:0] frontend_io_covSum ;  
   wire frontend_metaAssert ;  
   wire frontend_metaReset ;  
   wire frontend_icache_halt ;  
   wire frontend_fq_halt ;  
   wire frontend_tlb_halt ;  
   wire frontend_btb_halt ;  
   wire fpuOpt_clock ;  
   wire fpuOpt_reset ;  
   wire [31:0] fpuOpt_io_inst ;  
   wire [63:0] fpuOpt_io_fromint_data ;  
   wire [2:0] fpuOpt_io_fcsr_rm ;  
   wire fpuOpt_io_fcsr_flags_valid ;  
   wire [4:0] fpuOpt_io_fcsr_flags_bits ;  
   wire [63:0] fpuOpt_io_store_data ;  
   wire [63:0] fpuOpt_io_toint_data ;  
   wire fpuOpt_io_dmem_resp_val ;  
   wire [2:0] fpuOpt_io_dmem_resp_type ;  
   wire [4:0] fpuOpt_io_dmem_resp_tag ;  
   wire [63:0] fpuOpt_io_dmem_resp_data ;  
   wire fpuOpt_io_valid ;  
   wire fpuOpt_io_fcsr_rdy ;  
   wire fpuOpt_io_nack_mem ;  
   wire fpuOpt_io_illegal_rm ;  
   wire fpuOpt_io_killx ;  
   wire fpuOpt_io_killm ;  
   wire fpuOpt_io_dec_wen ;  
   wire fpuOpt_io_dec_ren1 ;  
   wire fpuOpt_io_dec_ren2 ;  
   wire fpuOpt_io_dec_ren3 ;  
   wire fpuOpt_io_sboard_set ;  
   wire fpuOpt_io_sboard_clr ;  
   wire [4:0] fpuOpt_io_sboard_clra ;  
   wire [29:0] fpuOpt_io_covSum ;  
   wire fpuOpt_metaAssert ;  
   wire fpuOpt_metaReset ;  
   wire fpuOpt_fpiu_halt ;  
   wire fpuOpt_ifpu_halt ;  
   wire fpuOpt_sfma_halt ;  
   wire fpuOpt_fpmu_halt ;  
   wire fpuOpt_divSqrt_1_halt ;  
   wire fpuOpt_dfma_halt ;  
   wire fpuOpt_divSqrt_halt ;  
   wire dcacheArb_clock ;  
   wire dcacheArb_io_requestor_0_req_ready ;  
   wire dcacheArb_io_requestor_0_req_valid ;  
   wire [39:0] dcacheArb_io_requestor_0_req_bits_addr ;  
   wire dcacheArb_io_requestor_0_s1_kill ;  
   wire dcacheArb_io_requestor_0_s2_nack ;  
   wire dcacheArb_io_requestor_0_resp_valid ;  
   wire [63:0] dcacheArb_io_requestor_0_resp_bits_data ;  
   wire dcacheArb_io_requestor_0_s2_xcpt_ae_ld ;  
   wire dcacheArb_io_requestor_1_req_ready ;  
   wire dcacheArb_io_requestor_1_req_valid ;  
   wire [39:0] dcacheArb_io_requestor_1_req_bits_addr ;  
   wire [6:0] dcacheArb_io_requestor_1_req_bits_tag ;  
   wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd ;  
   wire [1:0] dcacheArb_io_requestor_1_req_bits_size ;  
   wire dcacheArb_io_requestor_1_req_bits_signed ;  
   wire dcacheArb_io_requestor_1_s1_kill ;  
   wire [63:0] dcacheArb_io_requestor_1_s1_data_data ;  
   wire dcacheArb_io_requestor_1_s2_nack ;  
   wire dcacheArb_io_requestor_1_resp_valid ;  
   wire [6:0] dcacheArb_io_requestor_1_resp_bits_tag ;  
   wire [1:0] dcacheArb_io_requestor_1_resp_bits_size ;  
   wire [63:0] dcacheArb_io_requestor_1_resp_bits_data ;  
   wire dcacheArb_io_requestor_1_resp_bits_replay ;  
   wire dcacheArb_io_requestor_1_resp_bits_has_data ;  
   wire [63:0] dcacheArb_io_requestor_1_resp_bits_data_word_bypass ;  
   wire dcacheArb_io_requestor_1_replay_next ;  
   wire dcacheArb_io_requestor_1_s2_xcpt_ma_ld ;  
   wire dcacheArb_io_requestor_1_s2_xcpt_ma_st ;  
   wire dcacheArb_io_requestor_1_s2_xcpt_pf_ld ;  
   wire dcacheArb_io_requestor_1_s2_xcpt_pf_st ;  
   wire dcacheArb_io_requestor_1_s2_xcpt_ae_ld ;  
   wire dcacheArb_io_requestor_1_s2_xcpt_ae_st ;  
   wire dcacheArb_io_requestor_1_ordered ;  
   wire dcacheArb_io_requestor_1_perf_release ;  
   wire dcacheArb_io_requestor_1_perf_grant ;  
   wire dcacheArb_io_mem_req_ready ;  
   wire dcacheArb_io_mem_req_valid ;  
   wire [39:0] dcacheArb_io_mem_req_bits_addr ;  
   wire [6:0] dcacheArb_io_mem_req_bits_tag ;  
   wire [4:0] dcacheArb_io_mem_req_bits_cmd ;  
   wire [1:0] dcacheArb_io_mem_req_bits_size ;  
   wire dcacheArb_io_mem_req_bits_signed ;  
   wire dcacheArb_io_mem_req_bits_phys ;  
   wire dcacheArb_io_mem_s1_kill ;  
   wire [63:0] dcacheArb_io_mem_s1_data_data ;  
   wire dcacheArb_io_mem_s2_nack ;  
   wire dcacheArb_io_mem_resp_valid ;  
   wire [6:0] dcacheArb_io_mem_resp_bits_tag ;  
   wire [1:0] dcacheArb_io_mem_resp_bits_size ;  
   wire [63:0] dcacheArb_io_mem_resp_bits_data ;  
   wire dcacheArb_io_mem_resp_bits_replay ;  
   wire dcacheArb_io_mem_resp_bits_has_data ;  
   wire [63:0] dcacheArb_io_mem_resp_bits_data_word_bypass ;  
   wire dcacheArb_io_mem_replay_next ;  
   wire dcacheArb_io_mem_s2_xcpt_ma_ld ;  
   wire dcacheArb_io_mem_s2_xcpt_ma_st ;  
   wire dcacheArb_io_mem_s2_xcpt_pf_ld ;  
   wire dcacheArb_io_mem_s2_xcpt_pf_st ;  
   wire dcacheArb_io_mem_s2_xcpt_ae_ld ;  
   wire dcacheArb_io_mem_s2_xcpt_ae_st ;  
   wire dcacheArb_io_mem_ordered ;  
   wire dcacheArb_io_mem_perf_release ;  
   wire dcacheArb_io_mem_perf_grant ;  
   wire [29:0] dcacheArb_io_covSum ;  
   wire dcacheArb_metaAssert ;  
   wire dcacheArb_metaReset ;  
   wire ptw_clock ;  
   wire ptw_reset ;  
   wire ptw_io_requestor_0_req_ready ;  
   wire ptw_io_requestor_0_req_valid ;  
   wire [26:0] ptw_io_requestor_0_req_bits_bits_addr ;  
   wire ptw_io_requestor_0_resp_valid ;  
   wire ptw_io_requestor_0_resp_bits_ae ;  
   wire [53:0] ptw_io_requestor_0_resp_bits_pte_ppn ;  
   wire ptw_io_requestor_0_resp_bits_pte_d ;  
   wire ptw_io_requestor_0_resp_bits_pte_a ;  
   wire ptw_io_requestor_0_resp_bits_pte_g ;  
   wire ptw_io_requestor_0_resp_bits_pte_u ;  
   wire ptw_io_requestor_0_resp_bits_pte_x ;  
   wire ptw_io_requestor_0_resp_bits_pte_w ;  
   wire ptw_io_requestor_0_resp_bits_pte_r ;  
   wire ptw_io_requestor_0_resp_bits_pte_v ;  
   wire [1:0] ptw_io_requestor_0_resp_bits_level ;  
   wire ptw_io_requestor_0_resp_bits_homogeneous ;  
   wire [3:0] ptw_io_requestor_0_ptbr_mode ;  
   wire ptw_io_requestor_0_status_debug ;  
   wire [1:0] ptw_io_requestor_0_status_dprv ;  
   wire ptw_io_requestor_0_status_mxr ;  
   wire ptw_io_requestor_0_status_sum ;  
   wire ptw_io_requestor_0_pmp_0_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_0_cfg_a ;  
   wire ptw_io_requestor_0_pmp_0_cfg_x ;  
   wire ptw_io_requestor_0_pmp_0_cfg_w ;  
   wire ptw_io_requestor_0_pmp_0_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_0_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_0_mask ;  
   wire ptw_io_requestor_0_pmp_1_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_1_cfg_a ;  
   wire ptw_io_requestor_0_pmp_1_cfg_x ;  
   wire ptw_io_requestor_0_pmp_1_cfg_w ;  
   wire ptw_io_requestor_0_pmp_1_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_1_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_1_mask ;  
   wire ptw_io_requestor_0_pmp_2_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_2_cfg_a ;  
   wire ptw_io_requestor_0_pmp_2_cfg_x ;  
   wire ptw_io_requestor_0_pmp_2_cfg_w ;  
   wire ptw_io_requestor_0_pmp_2_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_2_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_2_mask ;  
   wire ptw_io_requestor_0_pmp_3_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_3_cfg_a ;  
   wire ptw_io_requestor_0_pmp_3_cfg_x ;  
   wire ptw_io_requestor_0_pmp_3_cfg_w ;  
   wire ptw_io_requestor_0_pmp_3_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_3_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_3_mask ;  
   wire ptw_io_requestor_0_pmp_4_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_4_cfg_a ;  
   wire ptw_io_requestor_0_pmp_4_cfg_x ;  
   wire ptw_io_requestor_0_pmp_4_cfg_w ;  
   wire ptw_io_requestor_0_pmp_4_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_4_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_4_mask ;  
   wire ptw_io_requestor_0_pmp_5_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_5_cfg_a ;  
   wire ptw_io_requestor_0_pmp_5_cfg_x ;  
   wire ptw_io_requestor_0_pmp_5_cfg_w ;  
   wire ptw_io_requestor_0_pmp_5_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_5_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_5_mask ;  
   wire ptw_io_requestor_0_pmp_6_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_6_cfg_a ;  
   wire ptw_io_requestor_0_pmp_6_cfg_x ;  
   wire ptw_io_requestor_0_pmp_6_cfg_w ;  
   wire ptw_io_requestor_0_pmp_6_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_6_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_6_mask ;  
   wire ptw_io_requestor_0_pmp_7_cfg_l ;  
   wire [1:0] ptw_io_requestor_0_pmp_7_cfg_a ;  
   wire ptw_io_requestor_0_pmp_7_cfg_x ;  
   wire ptw_io_requestor_0_pmp_7_cfg_w ;  
   wire ptw_io_requestor_0_pmp_7_cfg_r ;  
   wire [29:0] ptw_io_requestor_0_pmp_7_addr ;  
   wire [31:0] ptw_io_requestor_0_pmp_7_mask ;  
   wire ptw_io_requestor_1_req_ready ;  
   wire ptw_io_requestor_1_req_valid ;  
   wire ptw_io_requestor_1_req_bits_valid ;  
   wire [26:0] ptw_io_requestor_1_req_bits_bits_addr ;  
   wire ptw_io_requestor_1_resp_valid ;  
   wire ptw_io_requestor_1_resp_bits_ae ;  
   wire [53:0] ptw_io_requestor_1_resp_bits_pte_ppn ;  
   wire ptw_io_requestor_1_resp_bits_pte_d ;  
   wire ptw_io_requestor_1_resp_bits_pte_a ;  
   wire ptw_io_requestor_1_resp_bits_pte_g ;  
   wire ptw_io_requestor_1_resp_bits_pte_u ;  
   wire ptw_io_requestor_1_resp_bits_pte_x ;  
   wire ptw_io_requestor_1_resp_bits_pte_w ;  
   wire ptw_io_requestor_1_resp_bits_pte_r ;  
   wire ptw_io_requestor_1_resp_bits_pte_v ;  
   wire [1:0] ptw_io_requestor_1_resp_bits_level ;  
   wire ptw_io_requestor_1_resp_bits_homogeneous ;  
   wire [3:0] ptw_io_requestor_1_ptbr_mode ;  
   wire ptw_io_requestor_1_status_debug ;  
   wire [1:0] ptw_io_requestor_1_status_prv ;  
   wire ptw_io_requestor_1_pmp_0_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_0_cfg_a ;  
   wire ptw_io_requestor_1_pmp_0_cfg_x ;  
   wire ptw_io_requestor_1_pmp_0_cfg_w ;  
   wire ptw_io_requestor_1_pmp_0_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_0_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_0_mask ;  
   wire ptw_io_requestor_1_pmp_1_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_1_cfg_a ;  
   wire ptw_io_requestor_1_pmp_1_cfg_x ;  
   wire ptw_io_requestor_1_pmp_1_cfg_w ;  
   wire ptw_io_requestor_1_pmp_1_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_1_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_1_mask ;  
   wire ptw_io_requestor_1_pmp_2_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_2_cfg_a ;  
   wire ptw_io_requestor_1_pmp_2_cfg_x ;  
   wire ptw_io_requestor_1_pmp_2_cfg_w ;  
   wire ptw_io_requestor_1_pmp_2_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_2_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_2_mask ;  
   wire ptw_io_requestor_1_pmp_3_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_3_cfg_a ;  
   wire ptw_io_requestor_1_pmp_3_cfg_x ;  
   wire ptw_io_requestor_1_pmp_3_cfg_w ;  
   wire ptw_io_requestor_1_pmp_3_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_3_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_3_mask ;  
   wire ptw_io_requestor_1_pmp_4_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_4_cfg_a ;  
   wire ptw_io_requestor_1_pmp_4_cfg_x ;  
   wire ptw_io_requestor_1_pmp_4_cfg_w ;  
   wire ptw_io_requestor_1_pmp_4_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_4_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_4_mask ;  
   wire ptw_io_requestor_1_pmp_5_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_5_cfg_a ;  
   wire ptw_io_requestor_1_pmp_5_cfg_x ;  
   wire ptw_io_requestor_1_pmp_5_cfg_w ;  
   wire ptw_io_requestor_1_pmp_5_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_5_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_5_mask ;  
   wire ptw_io_requestor_1_pmp_6_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_6_cfg_a ;  
   wire ptw_io_requestor_1_pmp_6_cfg_x ;  
   wire ptw_io_requestor_1_pmp_6_cfg_w ;  
   wire ptw_io_requestor_1_pmp_6_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_6_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_6_mask ;  
   wire ptw_io_requestor_1_pmp_7_cfg_l ;  
   wire [1:0] ptw_io_requestor_1_pmp_7_cfg_a ;  
   wire ptw_io_requestor_1_pmp_7_cfg_x ;  
   wire ptw_io_requestor_1_pmp_7_cfg_w ;  
   wire ptw_io_requestor_1_pmp_7_cfg_r ;  
   wire [29:0] ptw_io_requestor_1_pmp_7_addr ;  
   wire [31:0] ptw_io_requestor_1_pmp_7_mask ;  
   wire [63:0] ptw_io_requestor_1_customCSRs_csrs_0_value ;  
   wire ptw_io_mem_req_ready ;  
   wire ptw_io_mem_req_valid ;  
   wire [39:0] ptw_io_mem_req_bits_addr ;  
   wire ptw_io_mem_s1_kill ;  
   wire ptw_io_mem_s2_nack ;  
   wire ptw_io_mem_resp_valid ;  
   wire [63:0] ptw_io_mem_resp_bits_data ;  
   wire ptw_io_mem_s2_xcpt_ae_ld ;  
   wire [3:0] ptw_io_dpath_ptbr_mode ;  
   wire [43:0] ptw_io_dpath_ptbr_ppn ;  
   wire ptw_io_dpath_sfence_valid ;  
   wire ptw_io_dpath_sfence_bits_rs1 ;  
   wire ptw_io_dpath_status_debug ;  
   wire [1:0] ptw_io_dpath_status_dprv ;  
   wire [1:0] ptw_io_dpath_status_prv ;  
   wire ptw_io_dpath_status_mxr ;  
   wire ptw_io_dpath_status_sum ;  
   wire ptw_io_dpath_pmp_0_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_0_cfg_a ;  
   wire ptw_io_dpath_pmp_0_cfg_x ;  
   wire ptw_io_dpath_pmp_0_cfg_w ;  
   wire ptw_io_dpath_pmp_0_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_0_addr ;  
   wire [31:0] ptw_io_dpath_pmp_0_mask ;  
   wire ptw_io_dpath_pmp_1_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_1_cfg_a ;  
   wire ptw_io_dpath_pmp_1_cfg_x ;  
   wire ptw_io_dpath_pmp_1_cfg_w ;  
   wire ptw_io_dpath_pmp_1_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_1_addr ;  
   wire [31:0] ptw_io_dpath_pmp_1_mask ;  
   wire ptw_io_dpath_pmp_2_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_2_cfg_a ;  
   wire ptw_io_dpath_pmp_2_cfg_x ;  
   wire ptw_io_dpath_pmp_2_cfg_w ;  
   wire ptw_io_dpath_pmp_2_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_2_addr ;  
   wire [31:0] ptw_io_dpath_pmp_2_mask ;  
   wire ptw_io_dpath_pmp_3_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_3_cfg_a ;  
   wire ptw_io_dpath_pmp_3_cfg_x ;  
   wire ptw_io_dpath_pmp_3_cfg_w ;  
   wire ptw_io_dpath_pmp_3_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_3_addr ;  
   wire [31:0] ptw_io_dpath_pmp_3_mask ;  
   wire ptw_io_dpath_pmp_4_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_4_cfg_a ;  
   wire ptw_io_dpath_pmp_4_cfg_x ;  
   wire ptw_io_dpath_pmp_4_cfg_w ;  
   wire ptw_io_dpath_pmp_4_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_4_addr ;  
   wire [31:0] ptw_io_dpath_pmp_4_mask ;  
   wire ptw_io_dpath_pmp_5_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_5_cfg_a ;  
   wire ptw_io_dpath_pmp_5_cfg_x ;  
   wire ptw_io_dpath_pmp_5_cfg_w ;  
   wire ptw_io_dpath_pmp_5_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_5_addr ;  
   wire [31:0] ptw_io_dpath_pmp_5_mask ;  
   wire ptw_io_dpath_pmp_6_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_6_cfg_a ;  
   wire ptw_io_dpath_pmp_6_cfg_x ;  
   wire ptw_io_dpath_pmp_6_cfg_w ;  
   wire ptw_io_dpath_pmp_6_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_6_addr ;  
   wire [31:0] ptw_io_dpath_pmp_6_mask ;  
   wire ptw_io_dpath_pmp_7_cfg_l ;  
   wire [1:0] ptw_io_dpath_pmp_7_cfg_a ;  
   wire ptw_io_dpath_pmp_7_cfg_x ;  
   wire ptw_io_dpath_pmp_7_cfg_w ;  
   wire ptw_io_dpath_pmp_7_cfg_r ;  
   wire [29:0] ptw_io_dpath_pmp_7_addr ;  
   wire [31:0] ptw_io_dpath_pmp_7_mask ;  
   wire ptw_io_dpath_perf_l2hit ;  
   wire ptw_io_dpath_perf_pte_miss ;  
   wire ptw_io_dpath_perf_pte_hit ;  
   wire [63:0] ptw_io_dpath_customCSRs_csrs_0_value ;  
   wire [29:0] ptw_io_covSum ;  
   wire ptw_metaAssert ;  
   wire ptw_metaReset ;  
   wire core_clock ;  
   wire core_reset ;  
   wire core_io_hartid ;  
   wire core_io_interrupts_debug ;  
   wire core_io_interrupts_mtip ;  
   wire core_io_interrupts_msip ;  
   wire core_io_interrupts_meip ;  
   wire core_io_interrupts_seip ;  
   wire core_io_imem_might_request ;  
   wire core_io_imem_req_valid ;  
   wire [39:0] core_io_imem_req_bits_pc ;  
   wire core_io_imem_req_bits_speculative ;  
   wire core_io_imem_sfence_valid ;  
   wire core_io_imem_sfence_bits_rs1 ;  
   wire core_io_imem_sfence_bits_rs2 ;  
   wire [38:0] core_io_imem_sfence_bits_addr ;  
   wire core_io_imem_resp_ready ;  
   wire core_io_imem_resp_valid ;  
   wire core_io_imem_resp_bits_btb_taken ;  
   wire core_io_imem_resp_bits_btb_bridx ;  
   wire [4:0] core_io_imem_resp_bits_btb_entry ;  
   wire [7:0] core_io_imem_resp_bits_btb_bht_history ;  
   wire [39:0] core_io_imem_resp_bits_pc ;  
   wire [31:0] core_io_imem_resp_bits_data ;  
   wire core_io_imem_resp_bits_xcpt_pf_inst ;  
   wire core_io_imem_resp_bits_xcpt_ae_inst ;  
   wire core_io_imem_resp_bits_replay ;  
   wire core_io_imem_btb_update_valid ;  
   wire [4:0] core_io_imem_btb_update_bits_prediction_entry ;  
   wire [38:0] core_io_imem_btb_update_bits_pc ;  
   wire core_io_imem_btb_update_bits_isValid ;  
   wire [38:0] core_io_imem_btb_update_bits_br_pc ;  
   wire [1:0] core_io_imem_btb_update_bits_cfiType ;  
   wire core_io_imem_bht_update_valid ;  
   wire [7:0] core_io_imem_bht_update_bits_prediction_history ;  
   wire [38:0] core_io_imem_bht_update_bits_pc ;  
   wire core_io_imem_bht_update_bits_branch ;  
   wire core_io_imem_bht_update_bits_taken ;  
   wire core_io_imem_bht_update_bits_mispredict ;  
   wire core_io_imem_flush_icache ;  
   wire core_io_dmem_req_ready ;  
   wire core_io_dmem_req_valid ;  
   wire [39:0] core_io_dmem_req_bits_addr ;  
   wire [6:0] core_io_dmem_req_bits_tag ;  
   wire [4:0] core_io_dmem_req_bits_cmd ;  
   wire [1:0] core_io_dmem_req_bits_size ;  
   wire core_io_dmem_req_bits_signed ;  
   wire core_io_dmem_s1_kill ;  
   wire [63:0] core_io_dmem_s1_data_data ;  
   wire core_io_dmem_s2_nack ;  
   wire core_io_dmem_resp_valid ;  
   wire [6:0] core_io_dmem_resp_bits_tag ;  
   wire [1:0] core_io_dmem_resp_bits_size ;  
   wire [63:0] core_io_dmem_resp_bits_data ;  
   wire core_io_dmem_resp_bits_replay ;  
   wire core_io_dmem_resp_bits_has_data ;  
   wire [63:0] core_io_dmem_resp_bits_data_word_bypass ;  
   wire core_io_dmem_replay_next ;  
   wire core_io_dmem_s2_xcpt_ma_ld ;  
   wire core_io_dmem_s2_xcpt_ma_st ;  
   wire core_io_dmem_s2_xcpt_pf_ld ;  
   wire core_io_dmem_s2_xcpt_pf_st ;  
   wire core_io_dmem_s2_xcpt_ae_ld ;  
   wire core_io_dmem_s2_xcpt_ae_st ;  
   wire core_io_dmem_ordered ;  
   wire core_io_dmem_perf_release ;  
   wire core_io_dmem_perf_grant ;  
   wire [3:0] core_io_ptw_ptbr_mode ;  
   wire [43:0] core_io_ptw_ptbr_ppn ;  
   wire core_io_ptw_sfence_valid ;  
   wire core_io_ptw_sfence_bits_rs1 ;  
   wire core_io_ptw_status_debug ;  
   wire [1:0] core_io_ptw_status_dprv ;  
   wire [1:0] core_io_ptw_status_prv ;  
   wire core_io_ptw_status_mxr ;  
   wire core_io_ptw_status_sum ;  
   wire core_io_ptw_pmp_0_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_0_cfg_a ;  
   wire core_io_ptw_pmp_0_cfg_x ;  
   wire core_io_ptw_pmp_0_cfg_w ;  
   wire core_io_ptw_pmp_0_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_0_addr ;  
   wire [31:0] core_io_ptw_pmp_0_mask ;  
   wire core_io_ptw_pmp_1_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_1_cfg_a ;  
   wire core_io_ptw_pmp_1_cfg_x ;  
   wire core_io_ptw_pmp_1_cfg_w ;  
   wire core_io_ptw_pmp_1_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_1_addr ;  
   wire [31:0] core_io_ptw_pmp_1_mask ;  
   wire core_io_ptw_pmp_2_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_2_cfg_a ;  
   wire core_io_ptw_pmp_2_cfg_x ;  
   wire core_io_ptw_pmp_2_cfg_w ;  
   wire core_io_ptw_pmp_2_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_2_addr ;  
   wire [31:0] core_io_ptw_pmp_2_mask ;  
   wire core_io_ptw_pmp_3_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_3_cfg_a ;  
   wire core_io_ptw_pmp_3_cfg_x ;  
   wire core_io_ptw_pmp_3_cfg_w ;  
   wire core_io_ptw_pmp_3_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_3_addr ;  
   wire [31:0] core_io_ptw_pmp_3_mask ;  
   wire core_io_ptw_pmp_4_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_4_cfg_a ;  
   wire core_io_ptw_pmp_4_cfg_x ;  
   wire core_io_ptw_pmp_4_cfg_w ;  
   wire core_io_ptw_pmp_4_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_4_addr ;  
   wire [31:0] core_io_ptw_pmp_4_mask ;  
   wire core_io_ptw_pmp_5_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_5_cfg_a ;  
   wire core_io_ptw_pmp_5_cfg_x ;  
   wire core_io_ptw_pmp_5_cfg_w ;  
   wire core_io_ptw_pmp_5_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_5_addr ;  
   wire [31:0] core_io_ptw_pmp_5_mask ;  
   wire core_io_ptw_pmp_6_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_6_cfg_a ;  
   wire core_io_ptw_pmp_6_cfg_x ;  
   wire core_io_ptw_pmp_6_cfg_w ;  
   wire core_io_ptw_pmp_6_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_6_addr ;  
   wire [31:0] core_io_ptw_pmp_6_mask ;  
   wire core_io_ptw_pmp_7_cfg_l ;  
   wire [1:0] core_io_ptw_pmp_7_cfg_a ;  
   wire core_io_ptw_pmp_7_cfg_x ;  
   wire core_io_ptw_pmp_7_cfg_w ;  
   wire core_io_ptw_pmp_7_cfg_r ;  
   wire [29:0] core_io_ptw_pmp_7_addr ;  
   wire [31:0] core_io_ptw_pmp_7_mask ;  
   wire [63:0] core_io_ptw_customCSRs_csrs_0_value ;  
   wire [31:0] core_io_fpu_inst ;  
   wire [63:0] core_io_fpu_fromint_data ;  
   wire [2:0] core_io_fpu_fcsr_rm ;  
   wire core_io_fpu_fcsr_flags_valid ;  
   wire [4:0] core_io_fpu_fcsr_flags_bits ;  
   wire [63:0] core_io_fpu_store_data ;  
   wire [63:0] core_io_fpu_toint_data ;  
   wire core_io_fpu_dmem_resp_val ;  
   wire [2:0] core_io_fpu_dmem_resp_type ;  
   wire [4:0] core_io_fpu_dmem_resp_tag ;  
   wire [63:0] core_io_fpu_dmem_resp_data ;  
   wire core_io_fpu_valid ;  
   wire core_io_fpu_fcsr_rdy ;  
   wire core_io_fpu_nack_mem ;  
   wire core_io_fpu_illegal_rm ;  
   wire core_io_fpu_killx ;  
   wire core_io_fpu_killm ;  
   wire core_io_fpu_dec_wen ;  
   wire core_io_fpu_dec_ren1 ;  
   wire core_io_fpu_dec_ren2 ;  
   wire core_io_fpu_dec_ren3 ;  
   wire core_io_fpu_sboard_set ;  
   wire core_io_fpu_sboard_clr ;  
   wire [4:0] core_io_fpu_sboard_clra ;  
   wire core_io_trace_0_valid ;  
   wire [39:0] core_io_trace_0_iaddr ;  
   wire [31:0] core_io_trace_0_insn ;  
   wire [2:0] core_io_trace_0_priv ;  
   wire core_io_trace_0_exception ;  
   wire core_io_trace_0_interrupt ;  
   wire [63:0] core_io_trace_0_cause ;  
   wire [39:0] core_io_trace_0_tval ;  
   wire core_io_wfi ;  
   wire [29:0] core_io_covSum ;  
   wire core_metaAssert ;  
   wire core_metaReset ;  
   wire core_PlusArgTimeout_halt ;  
   wire core_csr_halt ;  
   wire core_ibuf_halt ;  
   wire core_div_halt ;  
   reg bundleOut_0_0_REG ;  
   reg [31:0] _RAND_0 ;  
   wire [29:0] RocketTile_covSum ;  
   wire [29:0] tlMasterXbar_sum ;  
   wire [29:0] intXbar_sum ;  
   wire [29:0] fpuOpt_sum ;  
   wire [29:0] dcacheArb_sum ;  
   wire [29:0] frontend_sum ;  
   wire [29:0] dcache_sum ;  
   wire [29:0] broadcast_3_sum ;  
   wire [29:0] core_sum ;  
   wire [29:0] broadcast_sum ;  
   wire [29:0] broadcast_1_sum ;  
   wire [29:0] ptw_sum ;  
   wire ptw_metaAssert_wire ;  
   wire fpuOpt_metaAssert_wire ;  
   wire frontend_metaAssert_wire ;  
   wire dcacheArb_metaAssert_wire ;  
   wire broadcast_1_metaAssert_wire ;  
   wire broadcast_3_metaAssert_wire ;  
   wire intXbar_metaAssert_wire ;  
   wire core_metaAssert_wire ;  
   wire tlMasterXbar_metaAssert_wire ;  
   wire dcache_metaAssert_wire ;  
   wire broadcast_metaAssert_wire ;  
   wire RocketTile_or3 ;  
   wire RocketTile_or10 ;  
   wire RocketTile_or4 ;  
   wire RocketTile_or1 ;  
   wire RocketTile_or12 ;  
   wire RocketTile_or5 ;  
   wire RocketTile_or14 ;  
   wire RocketTile_or6 ;  
   wire RocketTile_or2 ;  
   wire RocketTile_or0 ;  
   reg RocketTile_metaAssert ;  
   reg [31:0] _RAND_1 ;  
  
wire  tlMasterXbar__clock;
wire  tlMasterXbar__reset;
wire  tlMasterXbar__auto_in_1_a_ready;
wire  tlMasterXbar__auto_in_1_a_valid;
wire [31:0] tlMasterXbar__auto_in_1_a_bits_address;
wire  tlMasterXbar__auto_in_1_d_valid;
wire [2:0] tlMasterXbar__auto_in_1_d_bits_opcode;
wire [3:0] tlMasterXbar__auto_in_1_d_bits_size;
wire [63:0] tlMasterXbar__auto_in_1_d_bits_data;
wire  tlMasterXbar__auto_in_1_d_bits_corrupt;
wire  tlMasterXbar__auto_in_0_a_ready;
wire  tlMasterXbar__auto_in_0_a_valid;
wire [2:0] tlMasterXbar__auto_in_0_a_bits_opcode;
wire [2:0] tlMasterXbar__auto_in_0_a_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_a_bits_size;
wire  tlMasterXbar__auto_in_0_a_bits_source;
wire [31:0] tlMasterXbar__auto_in_0_a_bits_address;
wire [7:0] tlMasterXbar__auto_in_0_a_bits_mask;
wire [63:0] tlMasterXbar__auto_in_0_a_bits_data;
wire  tlMasterXbar__auto_in_0_b_ready;
wire  tlMasterXbar__auto_in_0_b_valid;
wire [1:0] tlMasterXbar__auto_in_0_b_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_b_bits_size;
wire  tlMasterXbar__auto_in_0_b_bits_source;
wire [31:0] tlMasterXbar__auto_in_0_b_bits_address;
wire  tlMasterXbar__auto_in_0_c_ready;
wire  tlMasterXbar__auto_in_0_c_valid;
wire [2:0] tlMasterXbar__auto_in_0_c_bits_opcode;
wire [2:0] tlMasterXbar__auto_in_0_c_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_c_bits_size;
wire  tlMasterXbar__auto_in_0_c_bits_source;
wire [31:0] tlMasterXbar__auto_in_0_c_bits_address;
wire [63:0] tlMasterXbar__auto_in_0_c_bits_data;
wire  tlMasterXbar__auto_in_0_d_ready;
wire  tlMasterXbar__auto_in_0_d_valid;
wire [2:0] tlMasterXbar__auto_in_0_d_bits_opcode;
wire [1:0] tlMasterXbar__auto_in_0_d_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_d_bits_size;
wire  tlMasterXbar__auto_in_0_d_bits_source;
wire [1:0] tlMasterXbar__auto_in_0_d_bits_sink;
wire  tlMasterXbar__auto_in_0_d_bits_denied;
wire [63:0] tlMasterXbar__auto_in_0_d_bits_data;
wire  tlMasterXbar__auto_in_0_e_ready;
wire  tlMasterXbar__auto_in_0_e_valid;
wire [1:0] tlMasterXbar__auto_in_0_e_bits_sink;
wire  tlMasterXbar__auto_out_a_ready;
wire  tlMasterXbar__auto_out_a_valid;
wire [2:0] tlMasterXbar__auto_out_a_bits_opcode;
wire [2:0] tlMasterXbar__auto_out_a_bits_param;
wire [3:0] tlMasterXbar__auto_out_a_bits_size;
wire [1:0] tlMasterXbar__auto_out_a_bits_source;
wire [31:0] tlMasterXbar__auto_out_a_bits_address;
wire [7:0] tlMasterXbar__auto_out_a_bits_mask;
wire [63:0] tlMasterXbar__auto_out_a_bits_data;
wire  tlMasterXbar__auto_out_b_ready;
wire  tlMasterXbar__auto_out_b_valid;
wire [2:0] tlMasterXbar__auto_out_b_bits_opcode;
wire [1:0] tlMasterXbar__auto_out_b_bits_param;
wire [3:0] tlMasterXbar__auto_out_b_bits_size;
wire [1:0] tlMasterXbar__auto_out_b_bits_source;
wire [31:0] tlMasterXbar__auto_out_b_bits_address;
wire [7:0] tlMasterXbar__auto_out_b_bits_mask;
wire  tlMasterXbar__auto_out_b_bits_corrupt;
wire  tlMasterXbar__auto_out_c_ready;
wire  tlMasterXbar__auto_out_c_valid;
wire [2:0] tlMasterXbar__auto_out_c_bits_opcode;
wire [2:0] tlMasterXbar__auto_out_c_bits_param;
wire [3:0] tlMasterXbar__auto_out_c_bits_size;
wire [1:0] tlMasterXbar__auto_out_c_bits_source;
wire [31:0] tlMasterXbar__auto_out_c_bits_address;
wire [63:0] tlMasterXbar__auto_out_c_bits_data;
wire  tlMasterXbar__auto_out_d_ready;
wire  tlMasterXbar__auto_out_d_valid;
wire [2:0] tlMasterXbar__auto_out_d_bits_opcode;
wire [1:0] tlMasterXbar__auto_out_d_bits_param;
wire [3:0] tlMasterXbar__auto_out_d_bits_size;
wire [1:0] tlMasterXbar__auto_out_d_bits_source;
wire [1:0] tlMasterXbar__auto_out_d_bits_sink;
wire  tlMasterXbar__auto_out_d_bits_denied;
wire [63:0] tlMasterXbar__auto_out_d_bits_data;
wire  tlMasterXbar__auto_out_d_bits_corrupt;
wire  tlMasterXbar__auto_out_e_ready;
wire  tlMasterXbar__auto_out_e_valid;
wire [1:0] tlMasterXbar__auto_out_e_bits_sink;
wire [29:0] tlMasterXbar__io_covSum;
wire  tlMasterXbar__metaAssert;
wire  tlMasterXbar__metaReset;
wire  tlMasterXbar__monitor_halt;
wire  tlMasterXbar__monitor_1_halt;
 
   wire  tlMasterXbar__monitor_clock  ; 
   wire  tlMasterXbar__monitor_reset  ; 
   wire  tlMasterXbar__monitor_io_in_a_ready  ; 
   wire  tlMasterXbar__monitor_io_in_a_valid  ; 
   wire[2:0]  tlMasterXbar__monitor_io_in_a_bits_opcode  ; 
   wire[2:0]  tlMasterXbar__monitor_io_in_a_bits_param  ; 
   wire[3:0]  tlMasterXbar__monitor_io_in_a_bits_size  ; 
   wire  tlMasterXbar__monitor_io_in_a_bits_source  ; 
   wire[31:0]  tlMasterXbar__monitor_io_in_a_bits_address  ; 
   wire[7:0]  tlMasterXbar__monitor_io_in_a_bits_mask  ; 
   wire  tlMasterXbar__monitor_io_in_b_ready  ; 
   wire  tlMasterXbar__monitor_io_in_b_valid  ; 
   wire[2:0]  tlMasterXbar__monitor_io_in_b_bits_opcode  ; 
   wire[1:0]  tlMasterXbar__monitor_io_in_b_bits_param  ; 
   wire[3:0]  tlMasterXbar__monitor_io_in_b_bits_size  ; 
   wire  tlMasterXbar__monitor_io_in_b_bits_source  ; 
   wire[31:0]  tlMasterXbar__monitor_io_in_b_bits_address  ; 
   wire[7:0]  tlMasterXbar__monitor_io_in_b_bits_mask  ; 
   wire  tlMasterXbar__monitor_io_in_b_bits_corrupt  ; 
   wire  tlMasterXbar__monitor_io_in_c_ready  ; 
   wire  tlMasterXbar__monitor_io_in_c_valid  ; 
   wire[2:0]  tlMasterXbar__monitor_io_in_c_bits_opcode  ; 
   wire[2:0]  tlMasterXbar__monitor_io_in_c_bits_param  ; 
   wire[3:0]  tlMasterXbar__monitor_io_in_c_bits_size  ; 
   wire  tlMasterXbar__monitor_io_in_c_bits_source  ; 
   wire[31:0]  tlMasterXbar__monitor_io_in_c_bits_address  ; 
   wire  tlMasterXbar__monitor_io_in_d_ready  ; 
   wire  tlMasterXbar__monitor_io_in_d_valid  ; 
   wire[2:0]  tlMasterXbar__monitor_io_in_d_bits_opcode  ; 
   wire[1:0]  tlMasterXbar__monitor_io_in_d_bits_param  ; 
   wire[3:0]  tlMasterXbar__monitor_io_in_d_bits_size  ; 
   wire  tlMasterXbar__monitor_io_in_d_bits_source  ; 
   wire[1:0]  tlMasterXbar__monitor_io_in_d_bits_sink  ; 
   wire  tlMasterXbar__monitor_io_in_d_bits_denied  ; 
   wire  tlMasterXbar__monitor_io_in_d_bits_corrupt  ; 
   wire  tlMasterXbar__monitor_io_in_e_ready  ; 
   wire  tlMasterXbar__monitor_io_in_e_valid  ; 
   wire[1:0]  tlMasterXbar__monitor_io_in_e_bits_sink  ; 
   wire[29:0]  tlMasterXbar__monitor_io_covSum  ; 
   wire  tlMasterXbar__monitor_metaAssert  ; 
   wire  tlMasterXbar__monitor_metaReset  ; 
   wire  tlMasterXbar__monitor_1_clock  ; 
   wire  tlMasterXbar__monitor_1_reset  ; 
   wire  tlMasterXbar__monitor_1_io_in_a_ready  ; 
   wire  tlMasterXbar__monitor_1_io_in_a_valid  ; 
   wire[31:0]  tlMasterXbar__monitor_1_io_in_a_bits_address  ; 
   wire  tlMasterXbar__monitor_1_io_in_d_valid  ; 
   wire[2:0]  tlMasterXbar__monitor_1_io_in_d_bits_opcode  ; 
   wire[1:0]  tlMasterXbar__monitor_1_io_in_d_bits_param  ; 
   wire[3:0]  tlMasterXbar__monitor_1_io_in_d_bits_size  ; 
   wire[1:0]  tlMasterXbar__monitor_1_io_in_d_bits_sink  ; 
   wire  tlMasterXbar__monitor_1_io_in_d_bits_denied  ; 
   wire  tlMasterXbar__monitor_1_io_in_d_bits_corrupt  ; 
   wire[29:0]  tlMasterXbar__monitor_1_io_covSum  ; 
   wire  tlMasterXbar__monitor_1_metaAssert  ; 
   wire  tlMasterXbar__monitor_1_metaReset  ; 
   wire  tlMasterXbar__requestBOI_0_0  ; 
   wire  tlMasterXbar__requestDOI_0_0  ; 
   wire  tlMasterXbar__requestDOI_0_1  ; 
   wire[26:0]  tlMasterXbar___beatsAI_decode_T_1  ; 
   wire[8:0]  tlMasterXbar__beatsAI_decode  ; 
   wire  tlMasterXbar__beatsAI_opdata  ; 
   wire  tlMasterXbar___portsDIO_out_0_d_ready_T  ; 
   reg[8:0]  tlMasterXbar__beatsLeft  ; 
   reg[31:0]  tlMasterXbar___RAND_0  ; 
   wire  tlMasterXbar__idle  ; 
   wire  tlMasterXbar__latch  ; 
   wire[1:0]  tlMasterXbar__readys_filter_lo  ; 
   wire  tlMasterXbar___readys_T_1  ; 
   wire  tlMasterXbar___readys_T_3  ; 
   reg[1:0]  tlMasterXbar__readys_mask  ; 
   reg[31:0]  tlMasterXbar___RAND_1  ; 
   wire[1:0]  tlMasterXbar__readys_filter_hi  ; 
   wire[3:0]  tlMasterXbar__readys_filter  ; 
   wire[3:0]  tlMasterXbar___GEN_1  ; 
   wire[3:0]  tlMasterXbar___readys_unready_T_1  ; 
   wire[3:0]  tlMasterXbar___readys_unready_T_4  ; 
   wire[3:0]  tlMasterXbar___GEN_2  ; 
   wire[3:0]  tlMasterXbar__readys_unready  ; 
   wire[1:0]  tlMasterXbar___readys_readys_T_2  ; 
   wire[1:0]  tlMasterXbar__readys_readys  ; 
   wire  tlMasterXbar___readys_T_5  ; 
   wire  tlMasterXbar___readys_T_6  ; 
   wire[1:0]  tlMasterXbar___readys_mask_T  ; 
   wire[2:0]  tlMasterXbar___readys_mask_T_1  ; 
   wire[1:0]  tlMasterXbar___readys_mask_T_3  ; 
   wire  tlMasterXbar__readys_0  ; 
   wire  tlMasterXbar__readys_1  ; 
   wire  tlMasterXbar__earlyWinner_0  ; 
   wire  tlMasterXbar__earlyWinner_1  ; 
   wire  tlMasterXbar___prefixOR_T  ; 
   wire  tlMasterXbar___T_6  ; 
   wire  tlMasterXbar___T_9  ; 
   wire  tlMasterXbar___T_11  ; 
   wire  tlMasterXbar___T_14  ; 
   wire  tlMasterXbar___T_16  ; 
   wire  tlMasterXbar___T_21  ; 
   wire  tlMasterXbar___T_23  ; 
   reg  tlMasterXbar__state_0  ; 
   reg[31:0]  tlMasterXbar___RAND_2  ; 
   wire  tlMasterXbar__muxStateEarly_0  ; 
   reg  tlMasterXbar__state_1  ; 
   reg[31:0]  tlMasterXbar___RAND_3  ; 
   wire  tlMasterXbar__muxStateEarly_1  ; 
   wire  tlMasterXbar___out_0_a_earlyValid_T_1  ; 
   wire  tlMasterXbar___out_0_a_earlyValid_T_2  ; 
   wire  tlMasterXbar___out_0_a_earlyValid_T_3  ; 
   wire  tlMasterXbar__out_2_0_a_earlyValid  ; 
   wire  tlMasterXbar___beatsLeft_T_2  ; 
   wire[8:0]  tlMasterXbar___GEN_3  ; 
   wire[8:0]  tlMasterXbar___beatsLeft_T_4  ; 
   wire  tlMasterXbar__allowed_0  ; 
   wire  tlMasterXbar__allowed_1  ; 
   wire[7:0]  tlMasterXbar___T_31  ; 
   wire[7:0]  tlMasterXbar___T_32  ; 
   wire[31:0]  tlMasterXbar___T_34  ; 
   wire[31:0]  tlMasterXbar___T_35  ; 
   wire[1:0]  tlMasterXbar__in_0_a_bits_source  ; 
   wire[1:0]  tlMasterXbar___T_37  ; 
   wire[1:0]  tlMasterXbar___T_38  ; 
   wire[3:0]  tlMasterXbar___T_40  ; 
   wire[3:0]  tlMasterXbar___T_41  ; 
   wire[2:0]  tlMasterXbar___T_46  ; 
   wire[2:0]  tlMasterXbar___T_47  ; 
   reg[2:0]  tlMasterXbar__TLXbar_7_state  ; 
   reg[31:0]  tlMasterXbar___RAND_4  ; 
   reg  tlMasterXbar__TLXbar_7_cov  [0:7]; 
   reg[31:0]  tlMasterXbar___RAND_5  ; 
   wire  tlMasterXbar__TLXbar_7_cov_read_data  ; 
   wire[2:0]  tlMasterXbar__TLXbar_7_cov_read_addr  ; 
   wire  tlMasterXbar__TLXbar_7_cov_write_data  ; 
   wire[2:0]  tlMasterXbar__TLXbar_7_cov_write_addr  ; 
   wire  tlMasterXbar__TLXbar_7_cov_write_mask  ; 
   wire  tlMasterXbar__TLXbar_7_cov_write_en  ; 
   reg[29:0]  tlMasterXbar__TLXbar_7_covSum  ; 
   reg[31:0]  tlMasterXbar___RAND_6  ; 
   wire[1:0]  tlMasterXbar__readys_mask_shl  ; 
   wire[2:0]  tlMasterXbar__readys_mask_pad  ; 
   wire[2:0]  tlMasterXbar__state_0_shl  ; 
   wire[2:0]  tlMasterXbar__state_0_pad  ; 
   wire[2:0]  tlMasterXbar__state_1_shl  ; 
   wire[2:0]  tlMasterXbar__state_1_pad  ; 
   wire[2:0]  tlMasterXbar__TLXbar_7_xor2  ; 
   wire[2:0]  tlMasterXbar__TLXbar_7_xor0  ; 
   wire[29:0]  tlMasterXbar__monitor_sum  ; 
   wire[29:0]  tlMasterXbar__monitor_1_sum  ; 
   wire  tlMasterXbar__stopEn0  ; 
   wire  tlMasterXbar__stopEn1  ; 
   wire  tlMasterXbar__stopEn2  ; 
   wire  tlMasterXbar__stopEn3  ; 
   wire  tlMasterXbar__monitor_metaAssert_wire  ; 
   wire  tlMasterXbar__monitor_1_metaAssert_wire  ; 
   wire  tlMasterXbar__TLXbar_7_or4  ; 
   wire  tlMasterXbar__TLXbar_7_or1  ; 
   wire  tlMasterXbar__TLXbar_7_or6  ; 
   wire  tlMasterXbar__TLXbar_7_or2  ; 
   wire  tlMasterXbar__TLXbar_7_or0  ; 
   reg  tlMasterXbar__TLXbar_7_metaAssert  ; 
   reg[31:0]  tlMasterXbar___RAND_7  ;  
  
wire  tlMasterXbar__monitor__clock;
wire  tlMasterXbar__monitor__reset;
wire  tlMasterXbar__monitor__io_in_a_ready;
wire  tlMasterXbar__monitor__io_in_a_valid;
wire [2:0] tlMasterXbar__monitor__io_in_a_bits_opcode;
wire [2:0] tlMasterXbar__monitor__io_in_a_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_a_bits_size;
wire  tlMasterXbar__monitor__io_in_a_bits_source;
wire [31:0] tlMasterXbar__monitor__io_in_a_bits_address;
wire [7:0] tlMasterXbar__monitor__io_in_a_bits_mask;
wire  tlMasterXbar__monitor__io_in_b_ready;
wire  tlMasterXbar__monitor__io_in_b_valid;
wire [2:0] tlMasterXbar__monitor__io_in_b_bits_opcode;
wire [1:0] tlMasterXbar__monitor__io_in_b_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_b_bits_size;
wire  tlMasterXbar__monitor__io_in_b_bits_source;
wire [31:0] tlMasterXbar__monitor__io_in_b_bits_address;
wire [7:0] tlMasterXbar__monitor__io_in_b_bits_mask;
wire  tlMasterXbar__monitor__io_in_b_bits_corrupt;
wire  tlMasterXbar__monitor__io_in_c_ready;
wire  tlMasterXbar__monitor__io_in_c_valid;
wire [2:0] tlMasterXbar__monitor__io_in_c_bits_opcode;
wire [2:0] tlMasterXbar__monitor__io_in_c_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_c_bits_size;
wire  tlMasterXbar__monitor__io_in_c_bits_source;
wire [31:0] tlMasterXbar__monitor__io_in_c_bits_address;
wire  tlMasterXbar__monitor__io_in_d_ready;
wire  tlMasterXbar__monitor__io_in_d_valid;
wire [2:0] tlMasterXbar__monitor__io_in_d_bits_opcode;
wire [1:0] tlMasterXbar__monitor__io_in_d_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_d_bits_size;
wire  tlMasterXbar__monitor__io_in_d_bits_source;
wire [1:0] tlMasterXbar__monitor__io_in_d_bits_sink;
wire  tlMasterXbar__monitor__io_in_d_bits_denied;
wire  tlMasterXbar__monitor__io_in_d_bits_corrupt;
wire  tlMasterXbar__monitor__io_in_e_ready;
wire  tlMasterXbar__monitor__io_in_e_valid;
wire [1:0] tlMasterXbar__monitor__io_in_e_bits_sink;
wire [29:0] tlMasterXbar__monitor__io_covSum;
wire  tlMasterXbar__monitor__metaAssert;
wire  tlMasterXbar__monitor__metaReset;
 
   wire[31:0]  tlMasterXbar__monitor__plusarg_reader_out  ; 
   wire[31:0]  tlMasterXbar__monitor__plusarg_reader_1_out  ; 
   wire  tlMasterXbar__monitor__source_ok  ; 
   wire[26:0]  tlMasterXbar__monitor___is_aligned_mask_T_1  ; 
   wire[11:0]  tlMasterXbar__monitor__is_aligned_mask  ; 
   wire[31:0]  tlMasterXbar__monitor___GEN_86  ; 
   wire[31:0]  tlMasterXbar__monitor___is_aligned_T  ; 
   wire  tlMasterXbar__monitor__is_aligned  ; 
   wire[1:0]  tlMasterXbar__monitor__mask_sizeOH_shiftAmount  ; 
   wire[3:0]  tlMasterXbar__monitor___mask_sizeOH_T_1  ; 
   wire[2:0]  tlMasterXbar__monitor__mask_sizeOH  ; 
   wire  tlMasterXbar__monitor___mask_T  ; 
   wire  tlMasterXbar__monitor__mask_size  ; 
   wire  tlMasterXbar__monitor__mask_bit  ; 
   wire  tlMasterXbar__monitor__mask_nbit  ; 
   wire  tlMasterXbar__monitor___mask_acc_T  ; 
   wire  tlMasterXbar__monitor__mask_acc  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_1  ; 
   wire  tlMasterXbar__monitor__mask_acc_1  ; 
   wire  tlMasterXbar__monitor__mask_size_1  ; 
   wire  tlMasterXbar__monitor__mask_bit_1  ; 
   wire  tlMasterXbar__monitor__mask_nbit_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_2  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_2  ; 
   wire  tlMasterXbar__monitor__mask_acc_2  ; 
   wire  tlMasterXbar__monitor__mask_eq_3  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_3  ; 
   wire  tlMasterXbar__monitor__mask_acc_3  ; 
   wire  tlMasterXbar__monitor__mask_eq_4  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_4  ; 
   wire  tlMasterXbar__monitor__mask_acc_4  ; 
   wire  tlMasterXbar__monitor__mask_eq_5  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_5  ; 
   wire  tlMasterXbar__monitor__mask_acc_5  ; 
   wire  tlMasterXbar__monitor__mask_size_2  ; 
   wire  tlMasterXbar__monitor__mask_bit_2  ; 
   wire  tlMasterXbar__monitor__mask_nbit_2  ; 
   wire  tlMasterXbar__monitor__mask_eq_6  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_6  ; 
   wire  tlMasterXbar__monitor__mask_lo_lo_lo  ; 
   wire  tlMasterXbar__monitor__mask_eq_7  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_7  ; 
   wire  tlMasterXbar__monitor__mask_lo_lo_hi  ; 
   wire  tlMasterXbar__monitor__mask_eq_8  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_8  ; 
   wire  tlMasterXbar__monitor__mask_lo_hi_lo  ; 
   wire  tlMasterXbar__monitor__mask_eq_9  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_9  ; 
   wire  tlMasterXbar__monitor__mask_lo_hi_hi  ; 
   wire  tlMasterXbar__monitor__mask_eq_10  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_10  ; 
   wire  tlMasterXbar__monitor__mask_hi_lo_lo  ; 
   wire  tlMasterXbar__monitor__mask_eq_11  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_11  ; 
   wire  tlMasterXbar__monitor__mask_hi_lo_hi  ; 
   wire  tlMasterXbar__monitor__mask_eq_12  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_12  ; 
   wire  tlMasterXbar__monitor__mask_hi_hi_lo  ; 
   wire  tlMasterXbar__monitor__mask_eq_13  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_13  ; 
   wire  tlMasterXbar__monitor__mask_hi_hi_hi  ; 
   wire[7:0]  tlMasterXbar__monitor__mask  ; 
   wire[32:0]  tlMasterXbar__monitor___T_7  ; 
   wire  tlMasterXbar__monitor___T_24  ; 
   wire  tlMasterXbar__monitor___T_26  ; 
   wire  tlMasterXbar__monitor___T_31  ; 
   wire[32:0]  tlMasterXbar__monitor___T_37  ; 
   wire  tlMasterXbar__monitor___T_38  ; 
   wire[31:0]  tlMasterXbar__monitor___T_39  ; 
   wire[32:0]  tlMasterXbar__monitor___T_40  ; 
   wire[32:0]  tlMasterXbar__monitor___T_42  ; 
   wire  tlMasterXbar__monitor___T_43  ; 
   wire[31:0]  tlMasterXbar__monitor___T_44  ; 
   wire[32:0]  tlMasterXbar__monitor___T_45  ; 
   wire[32:0]  tlMasterXbar__monitor___T_47  ; 
   wire  tlMasterXbar__monitor___T_48  ; 
   wire[31:0]  tlMasterXbar__monitor___T_49  ; 
   wire[32:0]  tlMasterXbar__monitor___T_50  ; 
   wire[32:0]  tlMasterXbar__monitor___T_52  ; 
   wire  tlMasterXbar__monitor___T_53  ; 
   wire[31:0]  tlMasterXbar__monitor___T_54  ; 
   wire[32:0]  tlMasterXbar__monitor___T_55  ; 
   wire[32:0]  tlMasterXbar__monitor___T_57  ; 
   wire  tlMasterXbar__monitor___T_58  ; 
   wire[31:0]  tlMasterXbar__monitor___T_59  ; 
   wire[32:0]  tlMasterXbar__monitor___T_60  ; 
   wire[32:0]  tlMasterXbar__monitor___T_62  ; 
   wire  tlMasterXbar__monitor___T_63  ; 
   wire  tlMasterXbar__monitor___T_64  ; 
   wire  tlMasterXbar__monitor___T_65  ; 
   wire  tlMasterXbar__monitor___T_66  ; 
   wire  tlMasterXbar__monitor___T_67  ; 
   wire  tlMasterXbar__monitor___T_68  ; 
   wire  tlMasterXbar__monitor___T_71  ; 
   wire[31:0]  tlMasterXbar__monitor___T_74  ; 
   wire[32:0]  tlMasterXbar__monitor___T_75  ; 
   wire[32:0]  tlMasterXbar__monitor___T_77  ; 
   wire  tlMasterXbar__monitor___T_78  ; 
   wire  tlMasterXbar__monitor___T_79  ; 
   wire  tlMasterXbar__monitor___T_82  ; 
   wire  tlMasterXbar__monitor___T_84  ; 
   wire  tlMasterXbar__monitor___T_88  ; 
   wire  tlMasterXbar__monitor___T_89  ; 
   wire  tlMasterXbar__monitor___T_136  ; 
   wire  tlMasterXbar__monitor___T_137  ; 
   wire  tlMasterXbar__monitor___T_139  ; 
   wire  tlMasterXbar__monitor___T_141  ; 
   wire  tlMasterXbar__monitor___T_144  ; 
   wire  tlMasterXbar__monitor___T_148  ; 
   wire  tlMasterXbar__monitor___T_151  ; 
   wire  tlMasterXbar__monitor___T_153  ; 
   wire  tlMasterXbar__monitor___T_155  ; 
   wire  tlMasterXbar__monitor___T_158  ; 
   wire  tlMasterXbar__monitor___T_160  ; 
   wire  tlMasterXbar__monitor___T_166  ; 
   wire  tlMasterXbar__monitor___T_299  ; 
   wire  tlMasterXbar__monitor___T_301  ; 
   wire  tlMasterXbar__monitor___T_312  ; 
   wire  tlMasterXbar__monitor___T_322  ; 
   wire  tlMasterXbar__monitor___T_333  ; 
   wire  tlMasterXbar__monitor___T_368  ; 
   wire  tlMasterXbar__monitor___T_369  ; 
   wire  tlMasterXbar__monitor___T_370  ; 
   wire  tlMasterXbar__monitor___T_371  ; 
   wire  tlMasterXbar__monitor___T_372  ; 
   wire  tlMasterXbar__monitor___T_373  ; 
   wire  tlMasterXbar__monitor___T_375  ; 
   wire  tlMasterXbar__monitor___T_377  ; 
   wire  tlMasterXbar__monitor___T_385  ; 
   wire  tlMasterXbar__monitor___T_387  ; 
   wire  tlMasterXbar__monitor___T_389  ; 
   wire  tlMasterXbar__monitor___T_391  ; 
   wire  tlMasterXbar__monitor___T_397  ; 
   wire  tlMasterXbar__monitor___T_440  ; 
   wire  tlMasterXbar__monitor___T_441  ; 
   wire  tlMasterXbar__monitor___T_442  ; 
   wire  tlMasterXbar__monitor___T_443  ; 
   wire  tlMasterXbar__monitor___T_452  ; 
   wire  tlMasterXbar__monitor___T_460  ; 
   wire  tlMasterXbar__monitor___T_462  ; 
   wire  tlMasterXbar__monitor___T_464  ; 
   wire  tlMasterXbar__monitor___T_465  ; 
   wire  tlMasterXbar__monitor___T_467  ; 
   wire  tlMasterXbar__monitor___T_483  ; 
   wire[7:0]  tlMasterXbar__monitor___T_566  ; 
   wire  tlMasterXbar__monitor___T_567  ; 
   wire  tlMasterXbar__monitor___T_569  ; 
   wire  tlMasterXbar__monitor___T_571  ; 
   wire  tlMasterXbar__monitor___T_581  ; 
   wire  tlMasterXbar__monitor___T_605  ; 
   wire  tlMasterXbar__monitor___T_606  ; 
   wire  tlMasterXbar__monitor___T_607  ; 
   wire  tlMasterXbar__monitor___T_629  ; 
   wire  tlMasterXbar__monitor___T_631  ; 
   wire  tlMasterXbar__monitor___T_639  ; 
   wire  tlMasterXbar__monitor___T_641  ; 
   wire  tlMasterXbar__monitor___T_647  ; 
   wire  tlMasterXbar__monitor___T_715  ; 
   wire  tlMasterXbar__monitor___T_717  ; 
   wire  tlMasterXbar__monitor___T_723  ; 
   wire  tlMasterXbar__monitor___T_781  ; 
   wire  tlMasterXbar__monitor___T_783  ; 
   wire  tlMasterXbar__monitor___T_791  ; 
   wire  tlMasterXbar__monitor___T_793  ; 
   wire  tlMasterXbar__monitor___T_803  ; 
   wire  tlMasterXbar__monitor___T_805  ; 
   wire  tlMasterXbar__monitor__source_ok_1  ; 
   wire  tlMasterXbar__monitor___T_807  ; 
   wire  tlMasterXbar__monitor___T_809  ; 
   wire  tlMasterXbar__monitor___T_811  ; 
   wire  tlMasterXbar__monitor___T_813  ; 
   wire  tlMasterXbar__monitor___T_815  ; 
   wire  tlMasterXbar__monitor___T_817  ; 
   wire  tlMasterXbar__monitor___T_821  ; 
   wire  tlMasterXbar__monitor___T_825  ; 
   wire  tlMasterXbar__monitor___T_827  ; 
   wire  tlMasterXbar__monitor___T_838  ; 
   wire  tlMasterXbar__monitor___T_840  ; 
   wire  tlMasterXbar__monitor___T_842  ; 
   wire  tlMasterXbar__monitor___T_844  ; 
   wire  tlMasterXbar__monitor___T_855  ; 
   wire  tlMasterXbar__monitor___T_875  ; 
   wire  tlMasterXbar__monitor___T_877  ; 
   wire  tlMasterXbar__monitor___T_884  ; 
   wire  tlMasterXbar__monitor___T_901  ; 
   wire  tlMasterXbar__monitor___T_919  ; 
   wire  tlMasterXbar__monitor___T_936  ; 
   wire  tlMasterXbar__monitor___T_938  ; 
   wire[32:0]  tlMasterXbar__monitor___T_943  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_1  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_3  ; 
   wire  tlMasterXbar__monitor___address_ok_T_4  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_5  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_6  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_8  ; 
   wire  tlMasterXbar__monitor___address_ok_T_9  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_10  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_11  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_13  ; 
   wire  tlMasterXbar__monitor___address_ok_T_14  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_18  ; 
   wire  tlMasterXbar__monitor___address_ok_T_19  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_20  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_21  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_23  ; 
   wire  tlMasterXbar__monitor___address_ok_T_24  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_25  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_26  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_28  ; 
   wire  tlMasterXbar__monitor___address_ok_T_29  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_30  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_31  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_33  ; 
   wire  tlMasterXbar__monitor___address_ok_T_34  ; 
   wire  tlMasterXbar__monitor___address_ok_T_35  ; 
   wire  tlMasterXbar__monitor___address_ok_T_36  ; 
   wire  tlMasterXbar__monitor___address_ok_T_37  ; 
   wire  tlMasterXbar__monitor___address_ok_T_38  ; 
   wire  tlMasterXbar__monitor___address_ok_T_39  ; 
   wire  tlMasterXbar__monitor__address_ok  ; 
   wire[26:0]  tlMasterXbar__monitor___is_aligned_mask_T_4  ; 
   wire[11:0]  tlMasterXbar__monitor__is_aligned_mask_1  ; 
   wire[31:0]  tlMasterXbar__monitor___GEN_87  ; 
   wire[31:0]  tlMasterXbar__monitor___is_aligned_T_1  ; 
   wire  tlMasterXbar__monitor__is_aligned_1  ; 
   wire[1:0]  tlMasterXbar__monitor__mask_sizeOH_shiftAmount_1  ; 
   wire[3:0]  tlMasterXbar__monitor___mask_sizeOH_T_4  ; 
   wire[2:0]  tlMasterXbar__monitor__mask_sizeOH_1  ; 
   wire  tlMasterXbar__monitor___mask_T_1  ; 
   wire  tlMasterXbar__monitor__mask_size_3  ; 
   wire  tlMasterXbar__monitor__mask_bit_3  ; 
   wire  tlMasterXbar__monitor__mask_nbit_3  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_14  ; 
   wire  tlMasterXbar__monitor__mask_acc_6  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_15  ; 
   wire  tlMasterXbar__monitor__mask_acc_7  ; 
   wire  tlMasterXbar__monitor__mask_size_4  ; 
   wire  tlMasterXbar__monitor__mask_bit_4  ; 
   wire  tlMasterXbar__monitor__mask_nbit_4  ; 
   wire  tlMasterXbar__monitor__mask_eq_16  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_16  ; 
   wire  tlMasterXbar__monitor__mask_acc_8  ; 
   wire  tlMasterXbar__monitor__mask_eq_17  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_17  ; 
   wire  tlMasterXbar__monitor__mask_acc_9  ; 
   wire  tlMasterXbar__monitor__mask_eq_18  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_18  ; 
   wire  tlMasterXbar__monitor__mask_acc_10  ; 
   wire  tlMasterXbar__monitor__mask_eq_19  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_19  ; 
   wire  tlMasterXbar__monitor__mask_acc_11  ; 
   wire  tlMasterXbar__monitor__mask_size_5  ; 
   wire  tlMasterXbar__monitor__mask_bit_5  ; 
   wire  tlMasterXbar__monitor__mask_nbit_5  ; 
   wire  tlMasterXbar__monitor__mask_eq_20  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_20  ; 
   wire  tlMasterXbar__monitor__mask_lo_lo_lo_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_21  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_21  ; 
   wire  tlMasterXbar__monitor__mask_lo_lo_hi_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_22  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_22  ; 
   wire  tlMasterXbar__monitor__mask_lo_hi_lo_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_23  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_23  ; 
   wire  tlMasterXbar__monitor__mask_lo_hi_hi_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_24  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_24  ; 
   wire  tlMasterXbar__monitor__mask_hi_lo_lo_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_25  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_25  ; 
   wire  tlMasterXbar__monitor__mask_hi_lo_hi_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_26  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_26  ; 
   wire  tlMasterXbar__monitor__mask_hi_hi_lo_1  ; 
   wire  tlMasterXbar__monitor__mask_eq_27  ; 
   wire  tlMasterXbar__monitor___mask_acc_T_27  ; 
   wire  tlMasterXbar__monitor__mask_hi_hi_hi_1  ; 
   wire[7:0]  tlMasterXbar__monitor__mask_1  ; 
   wire  tlMasterXbar__monitor__legal_source  ; 
   wire  tlMasterXbar__monitor___T_960  ; 
   wire  tlMasterXbar__monitor___T_963  ; 
   wire  tlMasterXbar__monitor___T_964  ; 
   wire  tlMasterXbar__monitor___T_968  ; 
   wire  tlMasterXbar__monitor___T_1006  ; 
   wire  tlMasterXbar__monitor___T_1007  ; 
   wire  tlMasterXbar__monitor___T_1008  ; 
   wire  tlMasterXbar__monitor___T_1009  ; 
   wire  tlMasterXbar__monitor___T_1010  ; 
   wire  tlMasterXbar__monitor___T_1011  ; 
   wire  tlMasterXbar__monitor___T_1012  ; 
   wire  tlMasterXbar__monitor___T_1014  ; 
   wire  tlMasterXbar__monitor___T_1016  ; 
   wire  tlMasterXbar__monitor___T_1019  ; 
   wire  tlMasterXbar__monitor___T_1022  ; 
   wire  tlMasterXbar__monitor___T_1025  ; 
   wire  tlMasterXbar__monitor___T_1027  ; 
   wire  tlMasterXbar__monitor___T_1029  ; 
   wire  tlMasterXbar__monitor___T_1031  ; 
   wire  tlMasterXbar__monitor___T_1033  ; 
   wire  tlMasterXbar__monitor___T_1037  ; 
   wire  tlMasterXbar__monitor___T_1039  ; 
   wire  tlMasterXbar__monitor___T_1100  ; 
   wire  tlMasterXbar__monitor___T_1102  ; 
   wire  tlMasterXbar__monitor___T_1112  ; 
   wire  tlMasterXbar__monitor___T_1181  ; 
   wire[7:0]  tlMasterXbar__monitor___T_1247  ; 
   wire  tlMasterXbar__monitor___T_1248  ; 
   wire  tlMasterXbar__monitor___T_1250  ; 
   wire  tlMasterXbar__monitor___T_1252  ; 
   wire  tlMasterXbar__monitor___T_1321  ; 
   wire  tlMasterXbar__monitor___T_1390  ; 
   wire  tlMasterXbar__monitor__source_ok_2  ; 
   wire[26:0]  tlMasterXbar__monitor___is_aligned_mask_T_7  ; 
   wire[11:0]  tlMasterXbar__monitor__is_aligned_mask_2  ; 
   wire[31:0]  tlMasterXbar__monitor___GEN_88  ; 
   wire[31:0]  tlMasterXbar__monitor___is_aligned_T_2  ; 
   wire  tlMasterXbar__monitor__is_aligned_2  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_40  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_41  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_43  ; 
   wire  tlMasterXbar__monitor___address_ok_T_44  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_45  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_46  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_48  ; 
   wire  tlMasterXbar__monitor___address_ok_T_49  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_50  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_51  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_53  ; 
   wire  tlMasterXbar__monitor___address_ok_T_54  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_56  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_58  ; 
   wire  tlMasterXbar__monitor___address_ok_T_59  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_60  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_61  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_63  ; 
   wire  tlMasterXbar__monitor___address_ok_T_64  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_65  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_66  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_68  ; 
   wire  tlMasterXbar__monitor___address_ok_T_69  ; 
   wire[31:0]  tlMasterXbar__monitor___address_ok_T_70  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_71  ; 
   wire[32:0]  tlMasterXbar__monitor___address_ok_T_73  ; 
   wire  tlMasterXbar__monitor___address_ok_T_74  ; 
   wire  tlMasterXbar__monitor___address_ok_T_75  ; 
   wire  tlMasterXbar__monitor___address_ok_T_76  ; 
   wire  tlMasterXbar__monitor___address_ok_T_77  ; 
   wire  tlMasterXbar__monitor___address_ok_T_78  ; 
   wire  tlMasterXbar__monitor___address_ok_T_79  ; 
   wire  tlMasterXbar__monitor__address_ok_1  ; 
   wire  tlMasterXbar__monitor___T_1483  ; 
   wire  tlMasterXbar__monitor___T_1485  ; 
   wire  tlMasterXbar__monitor___T_1488  ; 
   wire  tlMasterXbar__monitor___T_1490  ; 
   wire  tlMasterXbar__monitor___T_1492  ; 
   wire  tlMasterXbar__monitor___T_1495  ; 
   wire  tlMasterXbar__monitor___T_1497  ; 
   wire  tlMasterXbar__monitor___T_1499  ; 
   wire  tlMasterXbar__monitor___T_1505  ; 
   wire  tlMasterXbar__monitor___T_1523  ; 
   wire  tlMasterXbar__monitor___T_1525  ; 
   wire  tlMasterXbar__monitor___T_1530  ; 
   wire  tlMasterXbar__monitor___T_1563  ; 
   wire  tlMasterXbar__monitor___T_1564  ; 
   wire  tlMasterXbar__monitor___T_1565  ; 
   wire  tlMasterXbar__monitor___T_1566  ; 
   wire  tlMasterXbar__monitor___T_1567  ; 
   wire  tlMasterXbar__monitor___T_1570  ; 
   wire  tlMasterXbar__monitor___T_1578  ; 
   wire  tlMasterXbar__monitor___T_1581  ; 
   wire  tlMasterXbar__monitor___T_1583  ; 
   wire  tlMasterXbar__monitor___T_1587  ; 
   wire  tlMasterXbar__monitor___T_1588  ; 
   wire  tlMasterXbar__monitor___T_1635  ; 
   wire  tlMasterXbar__monitor___T_1636  ; 
   wire  tlMasterXbar__monitor___T_1638  ; 
   wire  tlMasterXbar__monitor___T_1640  ; 
   wire  tlMasterXbar__monitor___T_1660  ; 
   wire  tlMasterXbar__monitor___T_1793  ; 
   wire  tlMasterXbar__monitor___T_1803  ; 
   wire  tlMasterXbar__monitor___T_1805  ; 
   wire  tlMasterXbar__monitor___T_1811  ; 
   wire  tlMasterXbar__monitor___T_1825  ; 
   wire  tlMasterXbar__monitor___a_first_T  ; 
   wire[8:0]  tlMasterXbar__monitor__a_first_beats1_decode  ; 
   wire  tlMasterXbar__monitor__a_first_beats1_opdata  ; 
   reg[8:0]  tlMasterXbar__monitor__a_first_counter  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_0  ; 
   wire[8:0]  tlMasterXbar__monitor__a_first_counter1  ; 
   wire  tlMasterXbar__monitor__a_first  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_1  ; 
   reg[2:0]  tlMasterXbar__monitor__param  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_2  ; 
   reg[3:0]  tlMasterXbar__monitor__size  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_3  ; 
   reg  tlMasterXbar__monitor__source  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_4  ; 
   reg[31:0]  tlMasterXbar__monitor__address  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_5  ; 
   wire  tlMasterXbar__monitor___T_1847  ; 
   wire  tlMasterXbar__monitor___T_1848  ; 
   wire  tlMasterXbar__monitor___T_1850  ; 
   wire  tlMasterXbar__monitor___T_1852  ; 
   wire  tlMasterXbar__monitor___T_1854  ; 
   wire  tlMasterXbar__monitor___T_1856  ; 
   wire  tlMasterXbar__monitor___T_1858  ; 
   wire  tlMasterXbar__monitor___T_1860  ; 
   wire  tlMasterXbar__monitor___T_1862  ; 
   wire  tlMasterXbar__monitor___T_1864  ; 
   wire  tlMasterXbar__monitor___T_1866  ; 
   wire  tlMasterXbar__monitor___T_1869  ; 
   wire  tlMasterXbar__monitor___d_first_T  ; 
   wire[26:0]  tlMasterXbar__monitor___d_first_beats1_decode_T_1  ; 
   wire[8:0]  tlMasterXbar__monitor__d_first_beats1_decode  ; 
   wire  tlMasterXbar__monitor__d_first_beats1_opdata  ; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_6  ; 
   wire[8:0]  tlMasterXbar__monitor__d_first_counter1  ; 
   wire  tlMasterXbar__monitor__d_first  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_7  ; 
   reg[1:0]  tlMasterXbar__monitor__param_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_8  ; 
   reg[3:0]  tlMasterXbar__monitor__size_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_9  ; 
   reg  tlMasterXbar__monitor__source_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_10  ; 
   reg[1:0]  tlMasterXbar__monitor__sink  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_11  ; 
   reg  tlMasterXbar__monitor__denied  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_12  ; 
   wire  tlMasterXbar__monitor___T_1871  ; 
   wire  tlMasterXbar__monitor___T_1872  ; 
   wire  tlMasterXbar__monitor___T_1874  ; 
   wire  tlMasterXbar__monitor___T_1876  ; 
   wire  tlMasterXbar__monitor___T_1878  ; 
   wire  tlMasterXbar__monitor___T_1880  ; 
   wire  tlMasterXbar__monitor___T_1882  ; 
   wire  tlMasterXbar__monitor___T_1884  ; 
   wire  tlMasterXbar__monitor___T_1886  ; 
   wire  tlMasterXbar__monitor___T_1888  ; 
   wire  tlMasterXbar__monitor___T_1890  ; 
   wire  tlMasterXbar__monitor___T_1892  ; 
   wire  tlMasterXbar__monitor___T_1894  ; 
   wire  tlMasterXbar__monitor___T_1897  ; 
   wire  tlMasterXbar__monitor__b_first_done  ; 
   reg[8:0]  tlMasterXbar__monitor__b_first_counter  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_13  ; 
   wire[8:0]  tlMasterXbar__monitor__b_first_counter1  ; 
   wire  tlMasterXbar__monitor__b_first  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode_2  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_14  ; 
   reg[1:0]  tlMasterXbar__monitor__param_2  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_15  ; 
   reg[3:0]  tlMasterXbar__monitor__size_2  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_16  ; 
   reg  tlMasterXbar__monitor__source_2  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_17  ; 
   reg[31:0]  tlMasterXbar__monitor__address_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_18  ; 
   wire  tlMasterXbar__monitor___T_1899  ; 
   wire  tlMasterXbar__monitor___T_1900  ; 
   wire  tlMasterXbar__monitor___T_1902  ; 
   wire  tlMasterXbar__monitor___T_1904  ; 
   wire  tlMasterXbar__monitor___T_1906  ; 
   wire  tlMasterXbar__monitor___T_1908  ; 
   wire  tlMasterXbar__monitor___T_1910  ; 
   wire  tlMasterXbar__monitor___T_1912  ; 
   wire  tlMasterXbar__monitor___T_1914  ; 
   wire  tlMasterXbar__monitor___T_1916  ; 
   wire  tlMasterXbar__monitor___T_1918  ; 
   wire  tlMasterXbar__monitor___T_1921  ; 
   wire  tlMasterXbar__monitor___c_first_T  ; 
   wire[8:0]  tlMasterXbar__monitor__c_first_beats1_decode  ; 
   wire  tlMasterXbar__monitor__c_first_beats1_opdata  ; 
   reg[8:0]  tlMasterXbar__monitor__c_first_counter  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_19  ; 
   wire[8:0]  tlMasterXbar__monitor__c_first_counter1  ; 
   wire  tlMasterXbar__monitor__c_first  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode_3  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_20  ; 
   reg[2:0]  tlMasterXbar__monitor__param_3  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_21  ; 
   reg[3:0]  tlMasterXbar__monitor__size_3  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_22  ; 
   reg  tlMasterXbar__monitor__source_3  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_23  ; 
   reg[31:0]  tlMasterXbar__monitor__address_2  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_24  ; 
   wire  tlMasterXbar__monitor___T_1923  ; 
   wire  tlMasterXbar__monitor___T_1924  ; 
   wire  tlMasterXbar__monitor___T_1926  ; 
   wire  tlMasterXbar__monitor___T_1928  ; 
   wire  tlMasterXbar__monitor___T_1930  ; 
   wire  tlMasterXbar__monitor___T_1932  ; 
   wire  tlMasterXbar__monitor___T_1934  ; 
   wire  tlMasterXbar__monitor___T_1936  ; 
   wire  tlMasterXbar__monitor___T_1938  ; 
   wire  tlMasterXbar__monitor___T_1940  ; 
   wire  tlMasterXbar__monitor___T_1942  ; 
   wire  tlMasterXbar__monitor___T_1945  ; 
   reg[1:0]  tlMasterXbar__monitor__inflight  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_25  ; 
   reg[7:0]  tlMasterXbar__monitor__inflight_opcodes  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_26  ; 
   reg[15:0]  tlMasterXbar__monitor__inflight_sizes  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_27  ; 
   reg[8:0]  tlMasterXbar__monitor__a_first_counter_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_28  ; 
   wire[8:0]  tlMasterXbar__monitor__a_first_counter1_1  ; 
   wire  tlMasterXbar__monitor__a_first_1  ; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_29  ; 
   wire[8:0]  tlMasterXbar__monitor__d_first_counter1_1  ; 
   wire  tlMasterXbar__monitor__d_first_1  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_89  ; 
   wire[3:0]  tlMasterXbar__monitor___a_opcode_lookup_T  ; 
   wire[7:0]  tlMasterXbar__monitor___a_opcode_lookup_T_1  ; 
   wire[15:0]  tlMasterXbar__monitor___a_opcode_lookup_T_5  ; 
   wire[15:0]  tlMasterXbar__monitor___GEN_90  ; 
   wire[15:0]  tlMasterXbar__monitor___a_opcode_lookup_T_6  ; 
   wire[15:0]  tlMasterXbar__monitor___a_opcode_lookup_T_7  ; 
   wire[3:0]  tlMasterXbar__monitor___a_size_lookup_T  ; 
   wire[15:0]  tlMasterXbar__monitor___a_size_lookup_T_1  ; 
   wire[15:0]  tlMasterXbar__monitor___a_size_lookup_T_5  ; 
   wire[15:0]  tlMasterXbar__monitor___a_size_lookup_T_6  ; 
   wire[15:0]  tlMasterXbar__monitor___a_size_lookup_T_7  ; 
   wire  tlMasterXbar__monitor___T_1946  ; 
   wire[1:0]  tlMasterXbar__monitor___a_set_wo_ready_T  ; 
   wire[1:0]  tlMasterXbar__monitor__a_set_wo_ready  ; 
   wire  tlMasterXbar__monitor___T_1949  ; 
   wire[3:0]  tlMasterXbar__monitor___a_opcodes_set_interm_T  ; 
   wire[3:0]  tlMasterXbar__monitor___a_opcodes_set_interm_T_1  ; 
   wire[4:0]  tlMasterXbar__monitor___a_sizes_set_interm_T  ; 
   wire[4:0]  tlMasterXbar__monitor___a_sizes_set_interm_T_1  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_93  ; 
   wire[3:0]  tlMasterXbar__monitor___a_opcodes_set_T  ; 
   wire[3:0]  tlMasterXbar__monitor__a_opcodes_set_interm  ; 
   wire[18:0]  tlMasterXbar__monitor___GEN_94  ; 
   wire[18:0]  tlMasterXbar__monitor___a_opcodes_set_T_1  ; 
   wire[3:0]  tlMasterXbar__monitor___a_sizes_set_T  ; 
   wire[4:0]  tlMasterXbar__monitor__a_sizes_set_interm  ; 
   wire[19:0]  tlMasterXbar__monitor___GEN_95  ; 
   wire[19:0]  tlMasterXbar__monitor___a_sizes_set_T_1  ; 
   wire[1:0]  tlMasterXbar__monitor___T_1951  ; 
   wire  tlMasterXbar__monitor___T_1955  ; 
   wire[1:0]  tlMasterXbar__monitor__a_set  ; 
   wire[18:0]  tlMasterXbar__monitor___GEN_31  ; 
   wire[19:0]  tlMasterXbar__monitor___GEN_32  ; 
   wire  tlMasterXbar__monitor___T_1957  ; 
   wire  tlMasterXbar__monitor___T_1960  ; 
   wire[1:0]  tlMasterXbar__monitor___d_clr_wo_ready_T  ; 
   wire[1:0]  tlMasterXbar__monitor__d_clr_wo_ready  ; 
   wire  tlMasterXbar__monitor___T_1962  ; 
   wire  tlMasterXbar__monitor___T_1965  ; 
   wire[30:0]  tlMasterXbar__monitor___GEN_97  ; 
   wire[30:0]  tlMasterXbar__monitor___d_opcodes_clr_T_5  ; 
   wire[30:0]  tlMasterXbar__monitor___GEN_98  ; 
   wire[30:0]  tlMasterXbar__monitor___d_sizes_clr_T_5  ; 
   wire[1:0]  tlMasterXbar__monitor__d_clr  ; 
   wire[30:0]  tlMasterXbar__monitor___GEN_35  ; 
   wire[30:0]  tlMasterXbar__monitor___GEN_36  ; 
   wire  tlMasterXbar__monitor___same_cycle_resp_T_2  ; 
   wire  tlMasterXbar__monitor__same_cycle_resp  ; 
   wire[1:0]  tlMasterXbar__monitor___T_1970  ; 
   wire  tlMasterXbar__monitor___T_1972  ; 
   wire  tlMasterXbar__monitor___T_1974  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_39  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_40  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_41  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_42  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_43  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_44  ; 
   wire  tlMasterXbar__monitor___T_1976  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_51  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_52  ; 
   wire  tlMasterXbar__monitor___T_1977  ; 
   wire  tlMasterXbar__monitor___T_1978  ; 
   wire  tlMasterXbar__monitor___T_1980  ; 
   wire  tlMasterXbar__monitor___T_1982  ; 
   wire  tlMasterXbar__monitor___T_1984  ; 
   wire[3:0]  tlMasterXbar__monitor__a_opcode_lookup  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_55  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_56  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_57  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_58  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_59  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_60  ; 
   wire  tlMasterXbar__monitor___T_1987  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_67  ; 
   wire[2:0]  tlMasterXbar__monitor___GEN_68  ; 
   wire  tlMasterXbar__monitor___T_1989  ; 
   wire  tlMasterXbar__monitor___T_1990  ; 
   wire  tlMasterXbar__monitor___T_1992  ; 
   wire[7:0]  tlMasterXbar__monitor__a_size_lookup  ; 
   wire[7:0]  tlMasterXbar__monitor___GEN_99  ; 
   wire  tlMasterXbar__monitor___T_1994  ; 
   wire  tlMasterXbar__monitor___T_1996  ; 
   wire  tlMasterXbar__monitor___T_1999  ; 
   wire  tlMasterXbar__monitor___T_2000  ; 
   wire  tlMasterXbar__monitor___T_2002  ; 
   wire  tlMasterXbar__monitor___T_2004  ; 
   wire  tlMasterXbar__monitor___T_2006  ; 
   wire  tlMasterXbar__monitor___T_2008  ; 
   wire  tlMasterXbar__monitor___T_2010  ; 
   wire  tlMasterXbar__monitor___T_2011  ; 
   wire  tlMasterXbar__monitor___T_2013  ; 
   wire  tlMasterXbar__monitor___T_2015  ; 
   wire[1:0]  tlMasterXbar__monitor___inflight_T  ; 
   wire[1:0]  tlMasterXbar__monitor___inflight_T_2  ; 
   wire[7:0]  tlMasterXbar__monitor__a_opcodes_set  ; 
   wire[7:0]  tlMasterXbar__monitor___inflight_opcodes_T  ; 
   wire[7:0]  tlMasterXbar__monitor__d_opcodes_clr  ; 
   wire[7:0]  tlMasterXbar__monitor___inflight_opcodes_T_2  ; 
   wire[15:0]  tlMasterXbar__monitor__a_sizes_set  ; 
   wire[15:0]  tlMasterXbar__monitor___inflight_sizes_T  ; 
   wire[15:0]  tlMasterXbar__monitor__d_sizes_clr  ; 
   wire[15:0]  tlMasterXbar__monitor___inflight_sizes_T_2  ; 
   reg[31:0]  tlMasterXbar__monitor__watchdog  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_30  ; 
   wire  tlMasterXbar__monitor___T_2017  ; 
   wire  tlMasterXbar__monitor___T_2019  ; 
   wire  tlMasterXbar__monitor___T_2020  ; 
   wire  tlMasterXbar__monitor___T_2021  ; 
   wire  tlMasterXbar__monitor___T_2022  ; 
   wire  tlMasterXbar__monitor___T_2024  ; 
   wire[31:0]  tlMasterXbar__monitor___watchdog_T_1  ; 
   wire  tlMasterXbar__monitor___T_2028  ; 
   reg[1:0]  tlMasterXbar__monitor__inflight_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_31  ; 
   reg[15:0]  tlMasterXbar__monitor__inflight_sizes_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_32  ; 
   reg[8:0]  tlMasterXbar__monitor__c_first_counter_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_33  ; 
   wire[8:0]  tlMasterXbar__monitor__c_first_counter1_1  ; 
   wire  tlMasterXbar__monitor__c_first_1  ; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter_2  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_34  ; 
   wire[8:0]  tlMasterXbar__monitor__d_first_counter1_2  ; 
   wire  tlMasterXbar__monitor__d_first_2  ; 
   wire[15:0]  tlMasterXbar__monitor___c_size_lookup_T_1  ; 
   wire[15:0]  tlMasterXbar__monitor___c_size_lookup_T_6  ; 
   wire[15:0]  tlMasterXbar__monitor___c_size_lookup_T_7  ; 
   wire  tlMasterXbar__monitor___T_2029  ; 
   wire  tlMasterXbar__monitor___T_2032  ; 
   wire  tlMasterXbar__monitor___T_2033  ; 
   wire[1:0]  tlMasterXbar__monitor___c_set_wo_ready_T  ; 
   wire[1:0]  tlMasterXbar__monitor__c_set_wo_ready  ; 
   wire  tlMasterXbar__monitor___T_2035  ; 
   wire  tlMasterXbar__monitor___T_2039  ; 
   wire[4:0]  tlMasterXbar__monitor___c_sizes_set_interm_T  ; 
   wire[4:0]  tlMasterXbar__monitor___c_sizes_set_interm_T_1  ; 
   wire[3:0]  tlMasterXbar__monitor___c_sizes_set_T  ; 
   wire[4:0]  tlMasterXbar__monitor__c_sizes_set_interm  ; 
   wire[19:0]  tlMasterXbar__monitor___GEN_106  ; 
   wire[19:0]  tlMasterXbar__monitor___c_sizes_set_T_1  ; 
   wire[1:0]  tlMasterXbar__monitor___T_2040  ; 
   wire  tlMasterXbar__monitor___T_2044  ; 
   wire[1:0]  tlMasterXbar__monitor__c_set  ; 
   wire[19:0]  tlMasterXbar__monitor___GEN_77  ; 
   wire  tlMasterXbar__monitor___T_2046  ; 
   wire  tlMasterXbar__monitor___T_2048  ; 
   wire[1:0]  tlMasterXbar__monitor__d_clr_wo_ready_1  ; 
   wire  tlMasterXbar__monitor___T_2050  ; 
   wire  tlMasterXbar__monitor___T_2052  ; 
   wire[1:0]  tlMasterXbar__monitor__d_clr_1  ; 
   wire[30:0]  tlMasterXbar__monitor___GEN_81  ; 
   wire  tlMasterXbar__monitor___same_cycle_resp_T_8  ; 
   wire  tlMasterXbar__monitor__same_cycle_resp_1  ; 
   wire[1:0]  tlMasterXbar__monitor___T_2056  ; 
   wire  tlMasterXbar__monitor___T_2058  ; 
   wire  tlMasterXbar__monitor___T_2060  ; 
   wire  tlMasterXbar__monitor___T_2062  ; 
   wire  tlMasterXbar__monitor___T_2064  ; 
   wire[7:0]  tlMasterXbar__monitor__c_size_lookup  ; 
   wire  tlMasterXbar__monitor___T_2066  ; 
   wire  tlMasterXbar__monitor___T_2068  ; 
   wire  tlMasterXbar__monitor___T_2071  ; 
   wire  tlMasterXbar__monitor___T_2072  ; 
   wire  tlMasterXbar__monitor___T_2074  ; 
   wire  tlMasterXbar__monitor___T_2075  ; 
   wire  tlMasterXbar__monitor___T_2077  ; 
   wire  tlMasterXbar__monitor___T_2079  ; 
   wire  tlMasterXbar__monitor___T_2081  ; 
   wire  tlMasterXbar__monitor___T_2082  ; 
   wire  tlMasterXbar__monitor___T_2084  ; 
   wire[1:0]  tlMasterXbar__monitor___inflight_T_3  ; 
   wire[1:0]  tlMasterXbar__monitor___inflight_T_5  ; 
   wire[15:0]  tlMasterXbar__monitor__c_sizes_set  ; 
   wire[15:0]  tlMasterXbar__monitor___inflight_sizes_T_3  ; 
   wire[15:0]  tlMasterXbar__monitor__d_sizes_clr_1  ; 
   wire[15:0]  tlMasterXbar__monitor___inflight_sizes_T_5  ; 
   reg[31:0]  tlMasterXbar__monitor__watchdog_1  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_35  ; 
   wire  tlMasterXbar__monitor___T_2086  ; 
   wire  tlMasterXbar__monitor___T_2088  ; 
   wire  tlMasterXbar__monitor___T_2089  ; 
   wire  tlMasterXbar__monitor___T_2090  ; 
   wire  tlMasterXbar__monitor___T_2091  ; 
   wire  tlMasterXbar__monitor___T_2093  ; 
   wire[31:0]  tlMasterXbar__monitor___watchdog_T_3  ; 
   wire  tlMasterXbar__monitor___T_2097  ; 
   reg[3:0]  tlMasterXbar__monitor__inflight_2  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_36  ; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter_3  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_37  ; 
   wire[8:0]  tlMasterXbar__monitor__d_first_counter1_3  ; 
   wire  tlMasterXbar__monitor__d_first_3  ; 
   wire  tlMasterXbar__monitor___T_2099  ; 
   wire  tlMasterXbar__monitor___T_2103  ; 
   wire  tlMasterXbar__monitor___T_2104  ; 
   wire[3:0]  tlMasterXbar__monitor___d_set_T  ; 
   wire[3:0]  tlMasterXbar__monitor___T_2105  ; 
   wire  tlMasterXbar__monitor___T_2109  ; 
   wire[3:0]  tlMasterXbar__monitor__d_set  ; 
   wire  tlMasterXbar__monitor___T_2111  ; 
   wire[3:0]  tlMasterXbar__monitor___e_clr_T  ; 
   wire[3:0]  tlMasterXbar__monitor___T_2114  ; 
   wire[3:0]  tlMasterXbar__monitor___T_2115  ; 
   wire  tlMasterXbar__monitor___T_2118  ; 
   wire[3:0]  tlMasterXbar__monitor__e_clr  ; 
   wire[3:0]  tlMasterXbar__monitor___inflight_T_6  ; 
   wire[3:0]  tlMasterXbar__monitor___inflight_T_8  ; 
   wire  tlMasterXbar__monitor___GEN_111  ; 
   wire  tlMasterXbar__monitor___GEN_125  ; 
   wire  tlMasterXbar__monitor___GEN_141  ; 
   wire  tlMasterXbar__monitor___GEN_153  ; 
   wire  tlMasterXbar__monitor___GEN_163  ; 
   wire  tlMasterXbar__monitor___GEN_173  ; 
   wire  tlMasterXbar__monitor___GEN_183  ; 
   wire  tlMasterXbar__monitor___GEN_193  ; 
   wire  tlMasterXbar__monitor___GEN_203  ; 
   wire  tlMasterXbar__monitor___GEN_213  ; 
   wire  tlMasterXbar__monitor___GEN_223  ; 
   wire  tlMasterXbar__monitor___GEN_233  ; 
   wire  tlMasterXbar__monitor___GEN_239  ; 
   wire  tlMasterXbar__monitor___GEN_245  ; 
   wire  tlMasterXbar__monitor___GEN_251  ; 
   wire  tlMasterXbar__monitor___GEN_265  ; 
   wire  tlMasterXbar__monitor___GEN_279  ; 
   wire  tlMasterXbar__monitor___GEN_291  ; 
   wire  tlMasterXbar__monitor___GEN_303  ; 
   wire  tlMasterXbar__monitor___GEN_313  ; 
   wire  tlMasterXbar__monitor___GEN_323  ; 
   wire  tlMasterXbar__monitor___GEN_335  ; 
   wire  tlMasterXbar__monitor___GEN_345  ; 
   wire  tlMasterXbar__monitor___GEN_355  ; 
   wire  tlMasterXbar__monitor___GEN_367  ; 
   wire  tlMasterXbar__monitor___GEN_379  ; 
   wire  tlMasterXbar__monitor___GEN_387  ; 
   wire  tlMasterXbar__monitor___GEN_395  ; 
   wire  tlMasterXbar__monitor___GEN_403  ; 
   wire  tlMasterXbar__monitor___GEN_408  ; 
   wire  tlMasterXbar__monitor___GEN_415  ; 
   wire  tlMasterXbar__monitor___GEN_418  ; 
   wire[29:0]  tlMasterXbar__monitor__TLMonitor_23_covSum  ; 
   wire  tlMasterXbar__monitor__stopEn0  ; 
   wire  tlMasterXbar__monitor__stopEn1  ; 
   wire  tlMasterXbar__monitor__stopEn2  ; 
   wire  tlMasterXbar__monitor__stopEn3  ; 
   wire  tlMasterXbar__monitor__stopEn4  ; 
   wire  tlMasterXbar__monitor__stopEn5  ; 
   wire  tlMasterXbar__monitor__stopEn6  ; 
   wire  tlMasterXbar__monitor__stopEn7  ; 
   wire  tlMasterXbar__monitor__stopEn8  ; 
   wire  tlMasterXbar__monitor__stopEn9  ; 
   wire  tlMasterXbar__monitor__stopEn10  ; 
   wire  tlMasterXbar__monitor__stopEn11  ; 
   wire  tlMasterXbar__monitor__stopEn12  ; 
   wire  tlMasterXbar__monitor__stopEn13  ; 
   wire  tlMasterXbar__monitor__stopEn14  ; 
   wire  tlMasterXbar__monitor__stopEn15  ; 
   wire  tlMasterXbar__monitor__stopEn16  ; 
   wire  tlMasterXbar__monitor__stopEn17  ; 
   wire  tlMasterXbar__monitor__stopEn18  ; 
   wire  tlMasterXbar__monitor__stopEn19  ; 
   wire  tlMasterXbar__monitor__stopEn20  ; 
   wire  tlMasterXbar__monitor__stopEn21  ; 
   wire  tlMasterXbar__monitor__stopEn22  ; 
   wire  tlMasterXbar__monitor__stopEn23  ; 
   wire  tlMasterXbar__monitor__stopEn24  ; 
   wire  tlMasterXbar__monitor__stopEn25  ; 
   wire  tlMasterXbar__monitor__stopEn26  ; 
   wire  tlMasterXbar__monitor__stopEn27  ; 
   wire  tlMasterXbar__monitor__stopEn28  ; 
   wire  tlMasterXbar__monitor__stopEn29  ; 
   wire  tlMasterXbar__monitor__stopEn30  ; 
   wire  tlMasterXbar__monitor__stopEn31  ; 
   wire  tlMasterXbar__monitor__stopEn32  ; 
   wire  tlMasterXbar__monitor__stopEn33  ; 
   wire  tlMasterXbar__monitor__stopEn34  ; 
   wire  tlMasterXbar__monitor__stopEn35  ; 
   wire  tlMasterXbar__monitor__stopEn36  ; 
   wire  tlMasterXbar__monitor__stopEn37  ; 
   wire  tlMasterXbar__monitor__stopEn38  ; 
   wire  tlMasterXbar__monitor__stopEn39  ; 
   wire  tlMasterXbar__monitor__stopEn40  ; 
   wire  tlMasterXbar__monitor__stopEn41  ; 
   wire  tlMasterXbar__monitor__stopEn42  ; 
   wire  tlMasterXbar__monitor__stopEn43  ; 
   wire  tlMasterXbar__monitor__stopEn44  ; 
   wire  tlMasterXbar__monitor__stopEn45  ; 
   wire  tlMasterXbar__monitor__stopEn46  ; 
   wire  tlMasterXbar__monitor__stopEn47  ; 
   wire  tlMasterXbar__monitor__stopEn48  ; 
   wire  tlMasterXbar__monitor__stopEn49  ; 
   wire  tlMasterXbar__monitor__stopEn50  ; 
   wire  tlMasterXbar__monitor__stopEn51  ; 
   wire  tlMasterXbar__monitor__stopEn52  ; 
   wire  tlMasterXbar__monitor__stopEn53  ; 
   wire  tlMasterXbar__monitor__stopEn54  ; 
   wire  tlMasterXbar__monitor__stopEn55  ; 
   wire  tlMasterXbar__monitor__stopEn56  ; 
   wire  tlMasterXbar__monitor__stopEn57  ; 
   wire  tlMasterXbar__monitor__stopEn58  ; 
   wire  tlMasterXbar__monitor__stopEn59  ; 
   wire  tlMasterXbar__monitor__stopEn60  ; 
   wire  tlMasterXbar__monitor__stopEn61  ; 
   wire  tlMasterXbar__monitor__stopEn62  ; 
   wire  tlMasterXbar__monitor__stopEn63  ; 
   wire  tlMasterXbar__monitor__stopEn64  ; 
   wire  tlMasterXbar__monitor__stopEn65  ; 
   wire  tlMasterXbar__monitor__stopEn66  ; 
   wire  tlMasterXbar__monitor__stopEn67  ; 
   wire  tlMasterXbar__monitor__stopEn68  ; 
   wire  tlMasterXbar__monitor__stopEn69  ; 
   wire  tlMasterXbar__monitor__stopEn70  ; 
   wire  tlMasterXbar__monitor__stopEn71  ; 
   wire  tlMasterXbar__monitor__stopEn72  ; 
   wire  tlMasterXbar__monitor__stopEn73  ; 
   wire  tlMasterXbar__monitor__stopEn74  ; 
   wire  tlMasterXbar__monitor__stopEn75  ; 
   wire  tlMasterXbar__monitor__stopEn76  ; 
   wire  tlMasterXbar__monitor__stopEn77  ; 
   wire  tlMasterXbar__monitor__stopEn78  ; 
   wire  tlMasterXbar__monitor__stopEn79  ; 
   wire  tlMasterXbar__monitor__stopEn80  ; 
   wire  tlMasterXbar__monitor__stopEn81  ; 
   wire  tlMasterXbar__monitor__stopEn82  ; 
   wire  tlMasterXbar__monitor__stopEn83  ; 
   wire  tlMasterXbar__monitor__stopEn84  ; 
   wire  tlMasterXbar__monitor__stopEn85  ; 
   wire  tlMasterXbar__monitor__stopEn86  ; 
   wire  tlMasterXbar__monitor__stopEn87  ; 
   wire  tlMasterXbar__monitor__stopEn88  ; 
   wire  tlMasterXbar__monitor__stopEn89  ; 
   wire  tlMasterXbar__monitor__stopEn90  ; 
   wire  tlMasterXbar__monitor__stopEn91  ; 
   wire  tlMasterXbar__monitor__stopEn92  ; 
   wire  tlMasterXbar__monitor__stopEn93  ; 
   wire  tlMasterXbar__monitor__stopEn94  ; 
   wire  tlMasterXbar__monitor__stopEn95  ; 
   wire  tlMasterXbar__monitor__stopEn96  ; 
   wire  tlMasterXbar__monitor__stopEn97  ; 
   wire  tlMasterXbar__monitor__stopEn98  ; 
   wire  tlMasterXbar__monitor__stopEn99  ; 
   wire  tlMasterXbar__monitor__stopEn100  ; 
   wire  tlMasterXbar__monitor__stopEn101  ; 
   wire  tlMasterXbar__monitor__stopEn102  ; 
   wire  tlMasterXbar__monitor__stopEn103  ; 
   wire  tlMasterXbar__monitor__stopEn104  ; 
   wire  tlMasterXbar__monitor__stopEn105  ; 
   wire  tlMasterXbar__monitor__stopEn106  ; 
   wire  tlMasterXbar__monitor__stopEn107  ; 
   wire  tlMasterXbar__monitor__stopEn108  ; 
   wire  tlMasterXbar__monitor__stopEn109  ; 
   wire  tlMasterXbar__monitor__stopEn110  ; 
   wire  tlMasterXbar__monitor__stopEn111  ; 
   wire  tlMasterXbar__monitor__stopEn112  ; 
   wire  tlMasterXbar__monitor__stopEn113  ; 
   wire  tlMasterXbar__monitor__stopEn114  ; 
   wire  tlMasterXbar__monitor__stopEn115  ; 
   wire  tlMasterXbar__monitor__stopEn116  ; 
   wire  tlMasterXbar__monitor__stopEn117  ; 
   wire  tlMasterXbar__monitor__stopEn118  ; 
   wire  tlMasterXbar__monitor__stopEn119  ; 
   wire  tlMasterXbar__monitor__stopEn120  ; 
   wire  tlMasterXbar__monitor__stopEn121  ; 
   wire  tlMasterXbar__monitor__stopEn122  ; 
   wire  tlMasterXbar__monitor__stopEn123  ; 
   wire  tlMasterXbar__monitor__stopEn124  ; 
   wire  tlMasterXbar__monitor__stopEn125  ; 
   wire  tlMasterXbar__monitor__stopEn126  ; 
   wire  tlMasterXbar__monitor__stopEn127  ; 
   wire  tlMasterXbar__monitor__stopEn128  ; 
   wire  tlMasterXbar__monitor__stopEn129  ; 
   wire  tlMasterXbar__monitor__stopEn130  ; 
   wire  tlMasterXbar__monitor__stopEn131  ; 
   wire  tlMasterXbar__monitor__stopEn132  ; 
   wire  tlMasterXbar__monitor__stopEn133  ; 
   wire  tlMasterXbar__monitor__stopEn134  ; 
   wire  tlMasterXbar__monitor__stopEn135  ; 
   wire  tlMasterXbar__monitor__stopEn136  ; 
   wire  tlMasterXbar__monitor__stopEn137  ; 
   wire  tlMasterXbar__monitor__stopEn138  ; 
   wire  tlMasterXbar__monitor__stopEn139  ; 
   wire  tlMasterXbar__monitor__stopEn140  ; 
   wire  tlMasterXbar__monitor__stopEn141  ; 
   wire  tlMasterXbar__monitor__stopEn142  ; 
   wire  tlMasterXbar__monitor__stopEn143  ; 
   wire  tlMasterXbar__monitor__stopEn144  ; 
   wire  tlMasterXbar__monitor__stopEn145  ; 
   wire  tlMasterXbar__monitor__stopEn146  ; 
   wire  tlMasterXbar__monitor__stopEn147  ; 
   wire  tlMasterXbar__monitor__stopEn148  ; 
   wire  tlMasterXbar__monitor__stopEn149  ; 
   wire  tlMasterXbar__monitor__stopEn150  ; 
   wire  tlMasterXbar__monitor__stopEn151  ; 
   wire  tlMasterXbar__monitor__stopEn152  ; 
   wire  tlMasterXbar__monitor__stopEn153  ; 
   wire  tlMasterXbar__monitor__stopEn154  ; 
   wire  tlMasterXbar__monitor__stopEn155  ; 
   wire  tlMasterXbar__monitor__stopEn156  ; 
   wire  tlMasterXbar__monitor__stopEn157  ; 
   wire  tlMasterXbar__monitor__stopEn158  ; 
   wire  tlMasterXbar__monitor__stopEn159  ; 
   wire  tlMasterXbar__monitor__stopEn160  ; 
   wire  tlMasterXbar__monitor__stopEn161  ; 
   wire  tlMasterXbar__monitor__stopEn162  ; 
   wire  tlMasterXbar__monitor__stopEn163  ; 
   wire  tlMasterXbar__monitor__stopEn164  ; 
   wire  tlMasterXbar__monitor__stopEn165  ; 
   wire  tlMasterXbar__monitor__stopEn166  ; 
   wire  tlMasterXbar__monitor__stopEn167  ; 
   wire  tlMasterXbar__monitor__stopEn168  ; 
   wire  tlMasterXbar__monitor__stopEn169  ; 
   wire  tlMasterXbar__monitor__stopEn170  ; 
   wire  tlMasterXbar__monitor__stopEn171  ; 
   wire  tlMasterXbar__monitor__stopEn172  ; 
   wire  tlMasterXbar__monitor__stopEn173  ; 
   wire  tlMasterXbar__monitor__stopEn174  ; 
   wire  tlMasterXbar__monitor__stopEn175  ; 
   wire  tlMasterXbar__monitor__stopEn176  ; 
   wire  tlMasterXbar__monitor__stopEn177  ; 
   wire  tlMasterXbar__monitor__stopEn178  ; 
   wire  tlMasterXbar__monitor__stopEn179  ; 
   wire  tlMasterXbar__monitor__stopEn180  ; 
   wire  tlMasterXbar__monitor__stopEn181  ; 
   wire  tlMasterXbar__monitor__stopEn182  ; 
   wire  tlMasterXbar__monitor__stopEn183  ; 
   wire  tlMasterXbar__monitor__stopEn184  ; 
   wire  tlMasterXbar__monitor__stopEn185  ; 
   wire  tlMasterXbar__monitor__stopEn186  ; 
   wire  tlMasterXbar__monitor__plusarg_reader_metaAssert_wire  ; 
   wire  tlMasterXbar__monitor__plusarg_reader_1_metaAssert_wire  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or63  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or130  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or64  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or31  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or132  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or65  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or134  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or66  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or32  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or15  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or136  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or67  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or138  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or68  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or33  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or140  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or69  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or142  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or70  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or34  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or16  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or7  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or144  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or71  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or146  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or72  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or35  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or148  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or73  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or150  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or74  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or36  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or17  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or152  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or75  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or154  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or76  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or37  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or156  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or77  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or158  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or78  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or38  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or18  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or8  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or3  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or79  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or162  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or80  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or39  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or164  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or81  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or166  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or82  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or40  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or19  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or168  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or83  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or170  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or84  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or41  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or172  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or85  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or174  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or86  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or42  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or20  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or9  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or176  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or87  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or178  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or88  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or43  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or180  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or89  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or182  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or90  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or44  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or21  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or184  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or91  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or186  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or92  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or45  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or188  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or93  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or190  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or94  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or46  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or22  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or10  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or4  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or1  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or95  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or194  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or96  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or47  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or196  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or97  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or198  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or98  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or48  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or23  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or200  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or99  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or202  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or100  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or49  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or204  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or101  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or206  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or102  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or50  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or24  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or11  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or208  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or103  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or210  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or104  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or51  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or212  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or105  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or214  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or106  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or52  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or25  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or216  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or107  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or218  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or108  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or53  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or220  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or109  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or222  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or110  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or54  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or26  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or12  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or5  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or224  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or111  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or226  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or112  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or55  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or228  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or113  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or230  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or114  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or56  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or27  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or232  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or115  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or234  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or116  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or57  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or236  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or117  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or238  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or118  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or58  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or28  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or13  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or240  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or119  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or242  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or120  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or59  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or244  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or121  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or246  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or122  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or60  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or29  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or248  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or123  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or250  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or124  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or61  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or252  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or125  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or254  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or126  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or62  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or30  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or14  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or6  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or2  ; 
   wire  tlMasterXbar__monitor__TLMonitor_23_or0  ; 
   reg  tlMasterXbar__monitor__TLMonitor_23_metaAssert  ; 
   reg[31:0]  tlMasterXbar__monitor___RAND_38  ; 
  assign   tlMasterXbar__monitor__source_ok  =~  tlMasterXbar__monitor__io_in_a_bits_source  |  tlMasterXbar__monitor__io_in_a_bits_source  ; 
  assign   tlMasterXbar__monitor___is_aligned_mask_T_1  =27'hfff<<  tlMasterXbar__monitor__io_in_a_bits_size  ; 
  assign   tlMasterXbar__monitor__is_aligned_mask  =~  tlMasterXbar__monitor___is_aligned_mask_T_1  [11:0]; 
  assign   tlMasterXbar__monitor___GEN_86  ={20'b0,  tlMasterXbar__monitor__is_aligned_mask  }; 
  assign   tlMasterXbar__monitor___is_aligned_T  =  tlMasterXbar__monitor__io_in_a_bits_address  &  tlMasterXbar__monitor___GEN_86  ; 
  assign   tlMasterXbar__monitor__is_aligned  =  tlMasterXbar__monitor___is_aligned_T  ==32'h0; 
  assign   tlMasterXbar__monitor__mask_sizeOH_shiftAmount  =  tlMasterXbar__monitor__io_in_a_bits_size  [1:0]; 
  assign   tlMasterXbar__monitor___mask_sizeOH_T_1  =4'h1<<  tlMasterXbar__monitor__mask_sizeOH_shiftAmount  ; 
  assign   tlMasterXbar__monitor__mask_sizeOH  =  tlMasterXbar__monitor___mask_sizeOH_T_1  [2:0]|3'h1; 
  assign   tlMasterXbar__monitor___mask_T  =  tlMasterXbar__monitor__io_in_a_bits_size  >=4'h3; 
  assign   tlMasterXbar__monitor__mask_size  =  tlMasterXbar__monitor__mask_sizeOH  [2]; 
  assign   tlMasterXbar__monitor__mask_bit  =  tlMasterXbar__monitor__io_in_a_bits_address  [2]; 
  assign   tlMasterXbar__monitor__mask_nbit  =~  tlMasterXbar__monitor__mask_bit  ; 
  assign   tlMasterXbar__monitor___mask_acc_T  =  tlMasterXbar__monitor__mask_size  &  tlMasterXbar__monitor__mask_nbit  ; 
  assign   tlMasterXbar__monitor__mask_acc  =  tlMasterXbar__monitor___mask_T  |  tlMasterXbar__monitor___mask_acc_T  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_1  =  tlMasterXbar__monitor__mask_size  &  tlMasterXbar__monitor__mask_bit  ; 
  assign   tlMasterXbar__monitor__mask_acc_1  =  tlMasterXbar__monitor___mask_T  |  tlMasterXbar__monitor___mask_acc_T_1  ; 
  assign   tlMasterXbar__monitor__mask_size_1  =  tlMasterXbar__monitor__mask_sizeOH  [1]; 
  assign   tlMasterXbar__monitor__mask_bit_1  =  tlMasterXbar__monitor__io_in_a_bits_address  [1]; 
  assign   tlMasterXbar__monitor__mask_nbit_1  =~  tlMasterXbar__monitor__mask_bit_1  ; 
  assign   tlMasterXbar__monitor__mask_eq_2  =  tlMasterXbar__monitor__mask_nbit  &  tlMasterXbar__monitor__mask_nbit_1  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_2  =  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_2  ; 
  assign   tlMasterXbar__monitor__mask_acc_2  =  tlMasterXbar__monitor__mask_acc  |  tlMasterXbar__monitor___mask_acc_T_2  ; 
  assign   tlMasterXbar__monitor__mask_eq_3  =  tlMasterXbar__monitor__mask_nbit  &  tlMasterXbar__monitor__mask_bit_1  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_3  =  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_3  ; 
  assign   tlMasterXbar__monitor__mask_acc_3  =  tlMasterXbar__monitor__mask_acc  |  tlMasterXbar__monitor___mask_acc_T_3  ; 
  assign   tlMasterXbar__monitor__mask_eq_4  =  tlMasterXbar__monitor__mask_bit  &  tlMasterXbar__monitor__mask_nbit_1  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_4  =  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_4  ; 
  assign   tlMasterXbar__monitor__mask_acc_4  =  tlMasterXbar__monitor__mask_acc_1  |  tlMasterXbar__monitor___mask_acc_T_4  ; 
  assign   tlMasterXbar__monitor__mask_eq_5  =  tlMasterXbar__monitor__mask_bit  &  tlMasterXbar__monitor__mask_bit_1  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_5  =  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_5  ; 
  assign   tlMasterXbar__monitor__mask_acc_5  =  tlMasterXbar__monitor__mask_acc_1  |  tlMasterXbar__monitor___mask_acc_T_5  ; 
  assign   tlMasterXbar__monitor__mask_size_2  =  tlMasterXbar__monitor__mask_sizeOH  [0]; 
  assign   tlMasterXbar__monitor__mask_bit_2  =  tlMasterXbar__monitor__io_in_a_bits_address  [0]; 
  assign   tlMasterXbar__monitor__mask_nbit_2  =~  tlMasterXbar__monitor__mask_bit_2  ; 
  assign   tlMasterXbar__monitor__mask_eq_6  =  tlMasterXbar__monitor__mask_eq_2  &  tlMasterXbar__monitor__mask_nbit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_6  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_6  ; 
  assign   tlMasterXbar__monitor__mask_lo_lo_lo  =  tlMasterXbar__monitor__mask_acc_2  |  tlMasterXbar__monitor___mask_acc_T_6  ; 
  assign   tlMasterXbar__monitor__mask_eq_7  =  tlMasterXbar__monitor__mask_eq_2  &  tlMasterXbar__monitor__mask_bit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_7  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_7  ; 
  assign   tlMasterXbar__monitor__mask_lo_lo_hi  =  tlMasterXbar__monitor__mask_acc_2  |  tlMasterXbar__monitor___mask_acc_T_7  ; 
  assign   tlMasterXbar__monitor__mask_eq_8  =  tlMasterXbar__monitor__mask_eq_3  &  tlMasterXbar__monitor__mask_nbit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_8  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_8  ; 
  assign   tlMasterXbar__monitor__mask_lo_hi_lo  =  tlMasterXbar__monitor__mask_acc_3  |  tlMasterXbar__monitor___mask_acc_T_8  ; 
  assign   tlMasterXbar__monitor__mask_eq_9  =  tlMasterXbar__monitor__mask_eq_3  &  tlMasterXbar__monitor__mask_bit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_9  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_9  ; 
  assign   tlMasterXbar__monitor__mask_lo_hi_hi  =  tlMasterXbar__monitor__mask_acc_3  |  tlMasterXbar__monitor___mask_acc_T_9  ; 
  assign   tlMasterXbar__monitor__mask_eq_10  =  tlMasterXbar__monitor__mask_eq_4  &  tlMasterXbar__monitor__mask_nbit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_10  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_10  ; 
  assign   tlMasterXbar__monitor__mask_hi_lo_lo  =  tlMasterXbar__monitor__mask_acc_4  |  tlMasterXbar__monitor___mask_acc_T_10  ; 
  assign   tlMasterXbar__monitor__mask_eq_11  =  tlMasterXbar__monitor__mask_eq_4  &  tlMasterXbar__monitor__mask_bit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_11  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_11  ; 
  assign   tlMasterXbar__monitor__mask_hi_lo_hi  =  tlMasterXbar__monitor__mask_acc_4  |  tlMasterXbar__monitor___mask_acc_T_11  ; 
  assign   tlMasterXbar__monitor__mask_eq_12  =  tlMasterXbar__monitor__mask_eq_5  &  tlMasterXbar__monitor__mask_nbit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_12  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_12  ; 
  assign   tlMasterXbar__monitor__mask_hi_hi_lo  =  tlMasterXbar__monitor__mask_acc_5  |  tlMasterXbar__monitor___mask_acc_T_12  ; 
  assign   tlMasterXbar__monitor__mask_eq_13  =  tlMasterXbar__monitor__mask_eq_5  &  tlMasterXbar__monitor__mask_bit_2  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_13  =  tlMasterXbar__monitor__mask_size_2  &  tlMasterXbar__monitor__mask_eq_13  ; 
  assign   tlMasterXbar__monitor__mask_hi_hi_hi  =  tlMasterXbar__monitor__mask_acc_5  |  tlMasterXbar__monitor___mask_acc_T_13  ; 
  assign   tlMasterXbar__monitor__mask  ={  tlMasterXbar__monitor__mask_hi_hi_hi  ,  tlMasterXbar__monitor__mask_hi_hi_lo  ,  tlMasterXbar__monitor__mask_hi_lo_hi  ,  tlMasterXbar__monitor__mask_hi_lo_lo  ,  tlMasterXbar__monitor__mask_lo_hi_hi  ,  tlMasterXbar__monitor__mask_lo_hi_lo  ,  tlMasterXbar__monitor__mask_lo_lo_hi  ,  tlMasterXbar__monitor__mask_lo_lo_lo  }; 
  assign   tlMasterXbar__monitor___T_7  ={1'b0,$signed(  tlMasterXbar__monitor__io_in_a_bits_address  )}; 
  assign   tlMasterXbar__monitor___T_24  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h6; 
  assign   tlMasterXbar__monitor___T_26  =  tlMasterXbar__monitor__io_in_a_bits_size  <=4'hc; 
  assign   tlMasterXbar__monitor___T_31  =  tlMasterXbar__monitor___T_26  &  tlMasterXbar__monitor__source_ok  ; 
  assign   tlMasterXbar__monitor___T_37  =$signed(  tlMasterXbar__monitor___T_7  )&-33'sh1000; 
  assign   tlMasterXbar__monitor___T_38  =$signed(  tlMasterXbar__monitor___T_37  )==33'sh0; 
  assign   tlMasterXbar__monitor___T_39  =  tlMasterXbar__monitor__io_in_a_bits_address  ^32'h3000; 
  assign   tlMasterXbar__monitor___T_40  ={1'b0,$signed(  tlMasterXbar__monitor___T_39  )}; 
  assign   tlMasterXbar__monitor___T_42  =$signed(  tlMasterXbar__monitor___T_40  )&-33'sh1000; 
  assign   tlMasterXbar__monitor___T_43  =$signed(  tlMasterXbar__monitor___T_42  )==33'sh0; 
  assign   tlMasterXbar__monitor___T_44  =  tlMasterXbar__monitor__io_in_a_bits_address  ^32'h10000; 
  assign   tlMasterXbar__monitor___T_45  ={1'b0,$signed(  tlMasterXbar__monitor___T_44  )}; 
  assign   tlMasterXbar__monitor___T_47  =$signed(  tlMasterXbar__monitor___T_45  )&-33'sh10000; 
  assign   tlMasterXbar__monitor___T_48  =$signed(  tlMasterXbar__monitor___T_47  )==33'sh0; 
  assign   tlMasterXbar__monitor___T_49  =  tlMasterXbar__monitor__io_in_a_bits_address  ^32'h2000000; 
  assign   tlMasterXbar__monitor___T_50  ={1'b0,$signed(  tlMasterXbar__monitor___T_49  )}; 
  assign   tlMasterXbar__monitor___T_52  =$signed(  tlMasterXbar__monitor___T_50  )&-33'sh10000; 
  assign   tlMasterXbar__monitor___T_53  =$signed(  tlMasterXbar__monitor___T_52  )==33'sh0; 
  assign   tlMasterXbar__monitor___T_54  =  tlMasterXbar__monitor__io_in_a_bits_address  ^32'hc000000; 
  assign   tlMasterXbar__monitor___T_55  ={1'b0,$signed(  tlMasterXbar__monitor___T_54  )}; 
  assign   tlMasterXbar__monitor___T_57  =$signed(  tlMasterXbar__monitor___T_55  )&-33'sh4000000; 
  assign   tlMasterXbar__monitor___T_58  =$signed(  tlMasterXbar__monitor___T_57  )==33'sh0; 
  assign   tlMasterXbar__monitor___T_59  =  tlMasterXbar__monitor__io_in_a_bits_address  ^32'h60000000; 
  assign   tlMasterXbar__monitor___T_60  ={1'b0,$signed(  tlMasterXbar__monitor___T_59  )}; 
  assign   tlMasterXbar__monitor___T_62  =$signed(  tlMasterXbar__monitor___T_60  )&-33'sh20000000; 
  assign   tlMasterXbar__monitor___T_63  =$signed(  tlMasterXbar__monitor___T_62  )==33'sh0; 
  assign   tlMasterXbar__monitor___T_64  =  tlMasterXbar__monitor___T_38  |  tlMasterXbar__monitor___T_43  ; 
  assign   tlMasterXbar__monitor___T_65  =  tlMasterXbar__monitor___T_64  |  tlMasterXbar__monitor___T_48  ; 
  assign   tlMasterXbar__monitor___T_66  =  tlMasterXbar__monitor___T_65  |  tlMasterXbar__monitor___T_53  ; 
  assign   tlMasterXbar__monitor___T_67  =  tlMasterXbar__monitor___T_66  |  tlMasterXbar__monitor___T_58  ; 
  assign   tlMasterXbar__monitor___T_68  =  tlMasterXbar__monitor___T_67  |  tlMasterXbar__monitor___T_63  ; 
  assign   tlMasterXbar__monitor___T_71  =  tlMasterXbar__monitor__io_in_a_bits_size  <=4'h6; 
  assign   tlMasterXbar__monitor___T_74  =  tlMasterXbar__monitor__io_in_a_bits_address  ^32'h80000000; 
  assign   tlMasterXbar__monitor___T_75  ={1'b0,$signed(  tlMasterXbar__monitor___T_74  )}; 
  assign   tlMasterXbar__monitor___T_77  =$signed(  tlMasterXbar__monitor___T_75  )&-33'sh10000000; 
  assign   tlMasterXbar__monitor___T_78  =$signed(  tlMasterXbar__monitor___T_77  )==33'sh0; 
  assign   tlMasterXbar__monitor___T_79  =  tlMasterXbar__monitor___T_71  &  tlMasterXbar__monitor___T_78  ; 
  assign   tlMasterXbar__monitor___T_82  =  tlMasterXbar__monitor___T_31  &  tlMasterXbar__monitor___T_79  ; 
  assign   tlMasterXbar__monitor___T_84  =  tlMasterXbar__monitor___T_82  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_88  =4'h6==  tlMasterXbar__monitor__io_in_a_bits_size  ; 
  assign   tlMasterXbar__monitor___T_89  =~  tlMasterXbar__monitor__io_in_a_bits_source  &  tlMasterXbar__monitor___T_88  ; 
  assign   tlMasterXbar__monitor___T_136  =  tlMasterXbar__monitor___T_68  |  tlMasterXbar__monitor___T_78  ; 
  assign   tlMasterXbar__monitor___T_137  =  tlMasterXbar__monitor___T_26  &  tlMasterXbar__monitor___T_136  ; 
  assign   tlMasterXbar__monitor___T_139  =  tlMasterXbar__monitor___T_89  &  tlMasterXbar__monitor___T_137  ; 
  assign   tlMasterXbar__monitor___T_141  =  tlMasterXbar__monitor___T_139  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_144  =  tlMasterXbar__monitor__source_ok  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_148  =  tlMasterXbar__monitor___mask_T  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_151  =  tlMasterXbar__monitor__is_aligned  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_153  =  tlMasterXbar__monitor__io_in_a_bits_param  <=3'h2; 
  assign   tlMasterXbar__monitor___T_155  =  tlMasterXbar__monitor___T_153  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_158  =~  tlMasterXbar__monitor__io_in_a_bits_mask  ==8'h0; 
  assign   tlMasterXbar__monitor___T_160  =  tlMasterXbar__monitor___T_158  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_166  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h7; 
  assign   tlMasterXbar__monitor___T_299  =  tlMasterXbar__monitor__io_in_a_bits_param  !=3'h0; 
  assign   tlMasterXbar__monitor___T_301  =  tlMasterXbar__monitor___T_299  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_312  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h4; 
  assign   tlMasterXbar__monitor___T_322  =  tlMasterXbar__monitor___T_31  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_333  =  tlMasterXbar__monitor___T_26  &  tlMasterXbar__monitor___T_43  ; 
  assign   tlMasterXbar__monitor___T_368  =  tlMasterXbar__monitor___T_38  |  tlMasterXbar__monitor___T_48  ; 
  assign   tlMasterXbar__monitor___T_369  =  tlMasterXbar__monitor___T_368  |  tlMasterXbar__monitor___T_53  ; 
  assign   tlMasterXbar__monitor___T_370  =  tlMasterXbar__monitor___T_369  |  tlMasterXbar__monitor___T_58  ; 
  assign   tlMasterXbar__monitor___T_371  =  tlMasterXbar__monitor___T_370  |  tlMasterXbar__monitor___T_63  ; 
  assign   tlMasterXbar__monitor___T_372  =  tlMasterXbar__monitor___T_371  |  tlMasterXbar__monitor___T_78  ; 
  assign   tlMasterXbar__monitor___T_373  =  tlMasterXbar__monitor___T_71  &  tlMasterXbar__monitor___T_372  ; 
  assign   tlMasterXbar__monitor___T_375  =  tlMasterXbar__monitor___T_333  |  tlMasterXbar__monitor___T_373  ; 
  assign   tlMasterXbar__monitor___T_377  =  tlMasterXbar__monitor___T_375  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_385  =  tlMasterXbar__monitor__io_in_a_bits_param  ==3'h0; 
  assign   tlMasterXbar__monitor___T_387  =  tlMasterXbar__monitor___T_385  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_389  =  tlMasterXbar__monitor__io_in_a_bits_mask  ==  tlMasterXbar__monitor__mask  ; 
  assign   tlMasterXbar__monitor___T_391  =  tlMasterXbar__monitor___T_389  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_397  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h0; 
  assign   tlMasterXbar__monitor___T_440  =  tlMasterXbar__monitor___T_38  |  tlMasterXbar__monitor___T_53  ; 
  assign   tlMasterXbar__monitor___T_441  =  tlMasterXbar__monitor___T_440  |  tlMasterXbar__monitor___T_58  ; 
  assign   tlMasterXbar__monitor___T_442  =  tlMasterXbar__monitor___T_441  |  tlMasterXbar__monitor___T_78  ; 
  assign   tlMasterXbar__monitor___T_443  =  tlMasterXbar__monitor___T_71  &  tlMasterXbar__monitor___T_442  ; 
  assign   tlMasterXbar__monitor___T_452  =  tlMasterXbar__monitor__io_in_a_bits_size  <=4'h8; 
  assign   tlMasterXbar__monitor___T_460  =  tlMasterXbar__monitor___T_452  &  tlMasterXbar__monitor___T_63  ; 
  assign   tlMasterXbar__monitor___T_462  =  tlMasterXbar__monitor___T_333  |  tlMasterXbar__monitor___T_443  ; 
  assign   tlMasterXbar__monitor___T_464  =  tlMasterXbar__monitor___T_462  |  tlMasterXbar__monitor___T_460  ; 
  assign   tlMasterXbar__monitor___T_465  =  tlMasterXbar__monitor___T_31  &  tlMasterXbar__monitor___T_464  ; 
  assign   tlMasterXbar__monitor___T_467  =  tlMasterXbar__monitor___T_465  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_483  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h1; 
  assign   tlMasterXbar__monitor___T_566  =  tlMasterXbar__monitor__io_in_a_bits_mask  &~  tlMasterXbar__monitor__mask  ; 
  assign   tlMasterXbar__monitor___T_567  =  tlMasterXbar__monitor___T_566  ==8'h0; 
  assign   tlMasterXbar__monitor___T_569  =  tlMasterXbar__monitor___T_567  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_571  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h2; 
  assign   tlMasterXbar__monitor___T_581  =  tlMasterXbar__monitor__io_in_a_bits_size  <=4'h3; 
  assign   tlMasterXbar__monitor___T_605  =  tlMasterXbar__monitor___T_64  |  tlMasterXbar__monitor___T_53  ; 
  assign   tlMasterXbar__monitor___T_606  =  tlMasterXbar__monitor___T_605  |  tlMasterXbar__monitor___T_58  ; 
  assign   tlMasterXbar__monitor___T_607  =  tlMasterXbar__monitor___T_581  &  tlMasterXbar__monitor___T_606  ; 
  assign   tlMasterXbar__monitor___T_629  =  tlMasterXbar__monitor___T_31  &  tlMasterXbar__monitor___T_607  ; 
  assign   tlMasterXbar__monitor___T_631  =  tlMasterXbar__monitor___T_629  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_639  =  tlMasterXbar__monitor__io_in_a_bits_param  <=3'h4; 
  assign   tlMasterXbar__monitor___T_641  =  tlMasterXbar__monitor___T_639  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_647  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h3; 
  assign   tlMasterXbar__monitor___T_715  =  tlMasterXbar__monitor__io_in_a_bits_param  <=3'h3; 
  assign   tlMasterXbar__monitor___T_717  =  tlMasterXbar__monitor___T_715  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_723  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h5; 
  assign   tlMasterXbar__monitor___T_781  =  tlMasterXbar__monitor___T_31  &  tlMasterXbar__monitor___T_333  ; 
  assign   tlMasterXbar__monitor___T_783  =  tlMasterXbar__monitor___T_781  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_791  =  tlMasterXbar__monitor__io_in_a_bits_param  <=3'h1; 
  assign   tlMasterXbar__monitor___T_793  =  tlMasterXbar__monitor___T_791  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_803  =  tlMasterXbar__monitor__io_in_d_bits_opcode  <=3'h6; 
  assign   tlMasterXbar__monitor___T_805  =  tlMasterXbar__monitor___T_803  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__source_ok_1  =~  tlMasterXbar__monitor__io_in_d_bits_source  |  tlMasterXbar__monitor__io_in_d_bits_source  ; 
  assign   tlMasterXbar__monitor___T_807  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h6; 
  assign   tlMasterXbar__monitor___T_809  =  tlMasterXbar__monitor__source_ok_1  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_811  =  tlMasterXbar__monitor__io_in_d_bits_size  >=4'h3; 
  assign   tlMasterXbar__monitor___T_813  =  tlMasterXbar__monitor___T_811  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_815  =  tlMasterXbar__monitor__io_in_d_bits_param  ==2'h0; 
  assign   tlMasterXbar__monitor___T_817  =  tlMasterXbar__monitor___T_815  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_821  =~  tlMasterXbar__monitor__io_in_d_bits_corrupt  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_825  =~  tlMasterXbar__monitor__io_in_d_bits_denied  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_827  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h4; 
  assign   tlMasterXbar__monitor___T_838  =  tlMasterXbar__monitor__io_in_d_bits_param  <=2'h2; 
  assign   tlMasterXbar__monitor___T_840  =  tlMasterXbar__monitor___T_838  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_842  =  tlMasterXbar__monitor__io_in_d_bits_param  !=2'h2; 
  assign   tlMasterXbar__monitor___T_844  =  tlMasterXbar__monitor___T_842  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_855  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h5; 
  assign   tlMasterXbar__monitor___T_875  =~  tlMasterXbar__monitor__io_in_d_bits_denied  |  tlMasterXbar__monitor__io_in_d_bits_corrupt  ; 
  assign   tlMasterXbar__monitor___T_877  =  tlMasterXbar__monitor___T_875  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_884  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h0; 
  assign   tlMasterXbar__monitor___T_901  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h1; 
  assign   tlMasterXbar__monitor___T_919  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h2; 
  assign   tlMasterXbar__monitor___T_936  =  tlMasterXbar__monitor__io_in_b_bits_opcode  <=3'h6; 
  assign   tlMasterXbar__monitor___T_938  =  tlMasterXbar__monitor___T_936  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_943  ={1'b0,$signed(  tlMasterXbar__monitor__io_in_b_bits_address  )}; 
  assign   tlMasterXbar__monitor___address_ok_T  =  tlMasterXbar__monitor__io_in_b_bits_address  ^32'h3000; 
  assign   tlMasterXbar__monitor___address_ok_T_1  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_3  =$signed(  tlMasterXbar__monitor___address_ok_T_1  )&-33'sh1000; 
  assign   tlMasterXbar__monitor___address_ok_T_4  =$signed(  tlMasterXbar__monitor___address_ok_T_3  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_5  =  tlMasterXbar__monitor__io_in_b_bits_address  ^32'hc000000; 
  assign   tlMasterXbar__monitor___address_ok_T_6  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_5  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_8  =$signed(  tlMasterXbar__monitor___address_ok_T_6  )&-33'sh4000000; 
  assign   tlMasterXbar__monitor___address_ok_T_9  =$signed(  tlMasterXbar__monitor___address_ok_T_8  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_10  =  tlMasterXbar__monitor__io_in_b_bits_address  ^32'h2000000; 
  assign   tlMasterXbar__monitor___address_ok_T_11  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_10  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_13  =$signed(  tlMasterXbar__monitor___address_ok_T_11  )&-33'sh10000; 
  assign   tlMasterXbar__monitor___address_ok_T_14  =$signed(  tlMasterXbar__monitor___address_ok_T_13  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_18  =$signed(  tlMasterXbar__monitor___T_943  )&-33'sh1000; 
  assign   tlMasterXbar__monitor___address_ok_T_19  =$signed(  tlMasterXbar__monitor___address_ok_T_18  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_20  =  tlMasterXbar__monitor__io_in_b_bits_address  ^32'h10000; 
  assign   tlMasterXbar__monitor___address_ok_T_21  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_20  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_23  =$signed(  tlMasterXbar__monitor___address_ok_T_21  )&-33'sh10000; 
  assign   tlMasterXbar__monitor___address_ok_T_24  =$signed(  tlMasterXbar__monitor___address_ok_T_23  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_25  =  tlMasterXbar__monitor__io_in_b_bits_address  ^32'h80000000; 
  assign   tlMasterXbar__monitor___address_ok_T_26  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_25  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_28  =$signed(  tlMasterXbar__monitor___address_ok_T_26  )&-33'sh10000000; 
  assign   tlMasterXbar__monitor___address_ok_T_29  =$signed(  tlMasterXbar__monitor___address_ok_T_28  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_30  =  tlMasterXbar__monitor__io_in_b_bits_address  ^32'h60000000; 
  assign   tlMasterXbar__monitor___address_ok_T_31  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_30  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_33  =$signed(  tlMasterXbar__monitor___address_ok_T_31  )&-33'sh20000000; 
  assign   tlMasterXbar__monitor___address_ok_T_34  =$signed(  tlMasterXbar__monitor___address_ok_T_33  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_35  =  tlMasterXbar__monitor___address_ok_T_4  |  tlMasterXbar__monitor___address_ok_T_9  ; 
  assign   tlMasterXbar__monitor___address_ok_T_36  =  tlMasterXbar__monitor___address_ok_T_35  |  tlMasterXbar__monitor___address_ok_T_14  ; 
  assign   tlMasterXbar__monitor___address_ok_T_37  =  tlMasterXbar__monitor___address_ok_T_36  |  tlMasterXbar__monitor___address_ok_T_19  ; 
  assign   tlMasterXbar__monitor___address_ok_T_38  =  tlMasterXbar__monitor___address_ok_T_37  |  tlMasterXbar__monitor___address_ok_T_24  ; 
  assign   tlMasterXbar__monitor___address_ok_T_39  =  tlMasterXbar__monitor___address_ok_T_38  |  tlMasterXbar__monitor___address_ok_T_29  ; 
  assign   tlMasterXbar__monitor__address_ok  =  tlMasterXbar__monitor___address_ok_T_39  |  tlMasterXbar__monitor___address_ok_T_34  ; 
  assign   tlMasterXbar__monitor___is_aligned_mask_T_4  =27'hfff<<  tlMasterXbar__monitor__io_in_b_bits_size  ; 
  assign   tlMasterXbar__monitor__is_aligned_mask_1  =~  tlMasterXbar__monitor___is_aligned_mask_T_4  [11:0]; 
  assign   tlMasterXbar__monitor___GEN_87  ={20'b0,  tlMasterXbar__monitor__is_aligned_mask_1  }; 
  assign   tlMasterXbar__monitor___is_aligned_T_1  =  tlMasterXbar__monitor__io_in_b_bits_address  &  tlMasterXbar__monitor___GEN_87  ; 
  assign   tlMasterXbar__monitor__is_aligned_1  =  tlMasterXbar__monitor___is_aligned_T_1  ==32'h0; 
  assign   tlMasterXbar__monitor__mask_sizeOH_shiftAmount_1  =  tlMasterXbar__monitor__io_in_b_bits_size  [1:0]; 
  assign   tlMasterXbar__monitor___mask_sizeOH_T_4  =4'h1<<  tlMasterXbar__monitor__mask_sizeOH_shiftAmount_1  ; 
  assign   tlMasterXbar__monitor__mask_sizeOH_1  =  tlMasterXbar__monitor___mask_sizeOH_T_4  [2:0]|3'h1; 
  assign   tlMasterXbar__monitor___mask_T_1  =  tlMasterXbar__monitor__io_in_b_bits_size  >=4'h3; 
  assign   tlMasterXbar__monitor__mask_size_3  =  tlMasterXbar__monitor__mask_sizeOH_1  [2]; 
  assign   tlMasterXbar__monitor__mask_bit_3  =  tlMasterXbar__monitor__io_in_b_bits_address  [2]; 
  assign   tlMasterXbar__monitor__mask_nbit_3  =~  tlMasterXbar__monitor__mask_bit_3  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_14  =  tlMasterXbar__monitor__mask_size_3  &  tlMasterXbar__monitor__mask_nbit_3  ; 
  assign   tlMasterXbar__monitor__mask_acc_6  =  tlMasterXbar__monitor___mask_T_1  |  tlMasterXbar__monitor___mask_acc_T_14  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_15  =  tlMasterXbar__monitor__mask_size_3  &  tlMasterXbar__monitor__mask_bit_3  ; 
  assign   tlMasterXbar__monitor__mask_acc_7  =  tlMasterXbar__monitor___mask_T_1  |  tlMasterXbar__monitor___mask_acc_T_15  ; 
  assign   tlMasterXbar__monitor__mask_size_4  =  tlMasterXbar__monitor__mask_sizeOH_1  [1]; 
  assign   tlMasterXbar__monitor__mask_bit_4  =  tlMasterXbar__monitor__io_in_b_bits_address  [1]; 
  assign   tlMasterXbar__monitor__mask_nbit_4  =~  tlMasterXbar__monitor__mask_bit_4  ; 
  assign   tlMasterXbar__monitor__mask_eq_16  =  tlMasterXbar__monitor__mask_nbit_3  &  tlMasterXbar__monitor__mask_nbit_4  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_16  =  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_16  ; 
  assign   tlMasterXbar__monitor__mask_acc_8  =  tlMasterXbar__monitor__mask_acc_6  |  tlMasterXbar__monitor___mask_acc_T_16  ; 
  assign   tlMasterXbar__monitor__mask_eq_17  =  tlMasterXbar__monitor__mask_nbit_3  &  tlMasterXbar__monitor__mask_bit_4  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_17  =  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_17  ; 
  assign   tlMasterXbar__monitor__mask_acc_9  =  tlMasterXbar__monitor__mask_acc_6  |  tlMasterXbar__monitor___mask_acc_T_17  ; 
  assign   tlMasterXbar__monitor__mask_eq_18  =  tlMasterXbar__monitor__mask_bit_3  &  tlMasterXbar__monitor__mask_nbit_4  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_18  =  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_18  ; 
  assign   tlMasterXbar__monitor__mask_acc_10  =  tlMasterXbar__monitor__mask_acc_7  |  tlMasterXbar__monitor___mask_acc_T_18  ; 
  assign   tlMasterXbar__monitor__mask_eq_19  =  tlMasterXbar__monitor__mask_bit_3  &  tlMasterXbar__monitor__mask_bit_4  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_19  =  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_19  ; 
  assign   tlMasterXbar__monitor__mask_acc_11  =  tlMasterXbar__monitor__mask_acc_7  |  tlMasterXbar__monitor___mask_acc_T_19  ; 
  assign   tlMasterXbar__monitor__mask_size_5  =  tlMasterXbar__monitor__mask_sizeOH_1  [0]; 
  assign   tlMasterXbar__monitor__mask_bit_5  =  tlMasterXbar__monitor__io_in_b_bits_address  [0]; 
  assign   tlMasterXbar__monitor__mask_nbit_5  =~  tlMasterXbar__monitor__mask_bit_5  ; 
  assign   tlMasterXbar__monitor__mask_eq_20  =  tlMasterXbar__monitor__mask_eq_16  &  tlMasterXbar__monitor__mask_nbit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_20  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_20  ; 
  assign   tlMasterXbar__monitor__mask_lo_lo_lo_1  =  tlMasterXbar__monitor__mask_acc_8  |  tlMasterXbar__monitor___mask_acc_T_20  ; 
  assign   tlMasterXbar__monitor__mask_eq_21  =  tlMasterXbar__monitor__mask_eq_16  &  tlMasterXbar__monitor__mask_bit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_21  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_21  ; 
  assign   tlMasterXbar__monitor__mask_lo_lo_hi_1  =  tlMasterXbar__monitor__mask_acc_8  |  tlMasterXbar__monitor___mask_acc_T_21  ; 
  assign   tlMasterXbar__monitor__mask_eq_22  =  tlMasterXbar__monitor__mask_eq_17  &  tlMasterXbar__monitor__mask_nbit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_22  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_22  ; 
  assign   tlMasterXbar__monitor__mask_lo_hi_lo_1  =  tlMasterXbar__monitor__mask_acc_9  |  tlMasterXbar__monitor___mask_acc_T_22  ; 
  assign   tlMasterXbar__monitor__mask_eq_23  =  tlMasterXbar__monitor__mask_eq_17  &  tlMasterXbar__monitor__mask_bit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_23  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_23  ; 
  assign   tlMasterXbar__monitor__mask_lo_hi_hi_1  =  tlMasterXbar__monitor__mask_acc_9  |  tlMasterXbar__monitor___mask_acc_T_23  ; 
  assign   tlMasterXbar__monitor__mask_eq_24  =  tlMasterXbar__monitor__mask_eq_18  &  tlMasterXbar__monitor__mask_nbit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_24  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_24  ; 
  assign   tlMasterXbar__monitor__mask_hi_lo_lo_1  =  tlMasterXbar__monitor__mask_acc_10  |  tlMasterXbar__monitor___mask_acc_T_24  ; 
  assign   tlMasterXbar__monitor__mask_eq_25  =  tlMasterXbar__monitor__mask_eq_18  &  tlMasterXbar__monitor__mask_bit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_25  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_25  ; 
  assign   tlMasterXbar__monitor__mask_hi_lo_hi_1  =  tlMasterXbar__monitor__mask_acc_10  |  tlMasterXbar__monitor___mask_acc_T_25  ; 
  assign   tlMasterXbar__monitor__mask_eq_26  =  tlMasterXbar__monitor__mask_eq_19  &  tlMasterXbar__monitor__mask_nbit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_26  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_26  ; 
  assign   tlMasterXbar__monitor__mask_hi_hi_lo_1  =  tlMasterXbar__monitor__mask_acc_11  |  tlMasterXbar__monitor___mask_acc_T_26  ; 
  assign   tlMasterXbar__monitor__mask_eq_27  =  tlMasterXbar__monitor__mask_eq_19  &  tlMasterXbar__monitor__mask_bit_5  ; 
  assign   tlMasterXbar__monitor___mask_acc_T_27  =  tlMasterXbar__monitor__mask_size_5  &  tlMasterXbar__monitor__mask_eq_27  ; 
  assign   tlMasterXbar__monitor__mask_hi_hi_hi_1  =  tlMasterXbar__monitor__mask_acc_11  |  tlMasterXbar__monitor___mask_acc_T_27  ; 
  assign   tlMasterXbar__monitor__mask_1  ={  tlMasterXbar__monitor__mask_hi_hi_hi_1  ,  tlMasterXbar__monitor__mask_hi_hi_lo_1  ,  tlMasterXbar__monitor__mask_hi_lo_hi_1  ,  tlMasterXbar__monitor__mask_hi_lo_lo_1  ,  tlMasterXbar__monitor__mask_lo_hi_hi_1  ,  tlMasterXbar__monitor__mask_lo_hi_lo_1  ,  tlMasterXbar__monitor__mask_lo_lo_hi_1  ,  tlMasterXbar__monitor__mask_lo_lo_lo_1  }; 
  assign   tlMasterXbar__monitor__legal_source  =  tlMasterXbar__monitor__io_in_b_bits_source  ==  tlMasterXbar__monitor__io_in_b_bits_source  ; 
  assign   tlMasterXbar__monitor___T_960  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h6; 
  assign   tlMasterXbar__monitor___T_963  =4'h6==  tlMasterXbar__monitor__io_in_b_bits_size  ; 
  assign   tlMasterXbar__monitor___T_964  =~  tlMasterXbar__monitor__io_in_b_bits_source  &  tlMasterXbar__monitor___T_963  ; 
  assign   tlMasterXbar__monitor___T_968  =  tlMasterXbar__monitor__io_in_b_bits_size  <=4'hc; 
  assign   tlMasterXbar__monitor___T_1006  =  tlMasterXbar__monitor___address_ok_T_19  |  tlMasterXbar__monitor___address_ok_T_4  ; 
  assign   tlMasterXbar__monitor___T_1007  =  tlMasterXbar__monitor___T_1006  |  tlMasterXbar__monitor___address_ok_T_24  ; 
  assign   tlMasterXbar__monitor___T_1008  =  tlMasterXbar__monitor___T_1007  |  tlMasterXbar__monitor___address_ok_T_14  ; 
  assign   tlMasterXbar__monitor___T_1009  =  tlMasterXbar__monitor___T_1008  |  tlMasterXbar__monitor___address_ok_T_9  ; 
  assign   tlMasterXbar__monitor___T_1010  =  tlMasterXbar__monitor___T_1009  |  tlMasterXbar__monitor___address_ok_T_34  ; 
  assign   tlMasterXbar__monitor___T_1011  =  tlMasterXbar__monitor___T_1010  |  tlMasterXbar__monitor___address_ok_T_29  ; 
  assign   tlMasterXbar__monitor___T_1012  =  tlMasterXbar__monitor___T_968  &  tlMasterXbar__monitor___T_1011  ; 
  assign   tlMasterXbar__monitor___T_1014  =  tlMasterXbar__monitor___T_964  &  tlMasterXbar__monitor___T_1012  ; 
  assign   tlMasterXbar__monitor___T_1016  =  tlMasterXbar__monitor___T_1014  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1019  =  tlMasterXbar__monitor__address_ok  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1022  =  tlMasterXbar__monitor__legal_source  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1025  =  tlMasterXbar__monitor__is_aligned_1  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1027  =  tlMasterXbar__monitor__io_in_b_bits_param  <=2'h2; 
  assign   tlMasterXbar__monitor___T_1029  =  tlMasterXbar__monitor___T_1027  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1031  =  tlMasterXbar__monitor__io_in_b_bits_mask  ==  tlMasterXbar__monitor__mask_1  ; 
  assign   tlMasterXbar__monitor___T_1033  =  tlMasterXbar__monitor___T_1031  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1037  =~  tlMasterXbar__monitor__io_in_b_bits_corrupt  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1039  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h4; 
  assign   tlMasterXbar__monitor___T_1100  =  tlMasterXbar__monitor__io_in_b_bits_param  ==2'h0; 
  assign   tlMasterXbar__monitor___T_1102  =  tlMasterXbar__monitor___T_1100  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1112  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h0; 
  assign   tlMasterXbar__monitor___T_1181  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h1; 
  assign   tlMasterXbar__monitor___T_1247  =  tlMasterXbar__monitor__io_in_b_bits_mask  &~  tlMasterXbar__monitor__mask_1  ; 
  assign   tlMasterXbar__monitor___T_1248  =  tlMasterXbar__monitor___T_1247  ==8'h0; 
  assign   tlMasterXbar__monitor___T_1250  =  tlMasterXbar__monitor___T_1248  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1252  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h2; 
  assign   tlMasterXbar__monitor___T_1321  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h3; 
  assign   tlMasterXbar__monitor___T_1390  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h5; 
  assign   tlMasterXbar__monitor__source_ok_2  =~  tlMasterXbar__monitor__io_in_c_bits_source  |  tlMasterXbar__monitor__io_in_c_bits_source  ; 
  assign   tlMasterXbar__monitor___is_aligned_mask_T_7  =27'hfff<<  tlMasterXbar__monitor__io_in_c_bits_size  ; 
  assign   tlMasterXbar__monitor__is_aligned_mask_2  =~  tlMasterXbar__monitor___is_aligned_mask_T_7  [11:0]; 
  assign   tlMasterXbar__monitor___GEN_88  ={20'b0,  tlMasterXbar__monitor__is_aligned_mask_2  }; 
  assign   tlMasterXbar__monitor___is_aligned_T_2  =  tlMasterXbar__monitor__io_in_c_bits_address  &  tlMasterXbar__monitor___GEN_88  ; 
  assign   tlMasterXbar__monitor__is_aligned_2  =  tlMasterXbar__monitor___is_aligned_T_2  ==32'h0; 
  assign   tlMasterXbar__monitor___address_ok_T_40  =  tlMasterXbar__monitor__io_in_c_bits_address  ^32'h3000; 
  assign   tlMasterXbar__monitor___address_ok_T_41  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_40  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_43  =$signed(  tlMasterXbar__monitor___address_ok_T_41  )&-33'sh1000; 
  assign   tlMasterXbar__monitor___address_ok_T_44  =$signed(  tlMasterXbar__monitor___address_ok_T_43  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_45  =  tlMasterXbar__monitor__io_in_c_bits_address  ^32'hc000000; 
  assign   tlMasterXbar__monitor___address_ok_T_46  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_45  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_48  =$signed(  tlMasterXbar__monitor___address_ok_T_46  )&-33'sh4000000; 
  assign   tlMasterXbar__monitor___address_ok_T_49  =$signed(  tlMasterXbar__monitor___address_ok_T_48  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_50  =  tlMasterXbar__monitor__io_in_c_bits_address  ^32'h2000000; 
  assign   tlMasterXbar__monitor___address_ok_T_51  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_50  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_53  =$signed(  tlMasterXbar__monitor___address_ok_T_51  )&-33'sh10000; 
  assign   tlMasterXbar__monitor___address_ok_T_54  =$signed(  tlMasterXbar__monitor___address_ok_T_53  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_56  ={1'b0,$signed(  tlMasterXbar__monitor__io_in_c_bits_address  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_58  =$signed(  tlMasterXbar__monitor___address_ok_T_56  )&-33'sh1000; 
  assign   tlMasterXbar__monitor___address_ok_T_59  =$signed(  tlMasterXbar__monitor___address_ok_T_58  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_60  =  tlMasterXbar__monitor__io_in_c_bits_address  ^32'h10000; 
  assign   tlMasterXbar__monitor___address_ok_T_61  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_60  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_63  =$signed(  tlMasterXbar__monitor___address_ok_T_61  )&-33'sh10000; 
  assign   tlMasterXbar__monitor___address_ok_T_64  =$signed(  tlMasterXbar__monitor___address_ok_T_63  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_65  =  tlMasterXbar__monitor__io_in_c_bits_address  ^32'h80000000; 
  assign   tlMasterXbar__monitor___address_ok_T_66  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_65  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_68  =$signed(  tlMasterXbar__monitor___address_ok_T_66  )&-33'sh10000000; 
  assign   tlMasterXbar__monitor___address_ok_T_69  =$signed(  tlMasterXbar__monitor___address_ok_T_68  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_70  =  tlMasterXbar__monitor__io_in_c_bits_address  ^32'h60000000; 
  assign   tlMasterXbar__monitor___address_ok_T_71  ={1'b0,$signed(  tlMasterXbar__monitor___address_ok_T_70  )}; 
  assign   tlMasterXbar__monitor___address_ok_T_73  =$signed(  tlMasterXbar__monitor___address_ok_T_71  )&-33'sh20000000; 
  assign   tlMasterXbar__monitor___address_ok_T_74  =$signed(  tlMasterXbar__monitor___address_ok_T_73  )==33'sh0; 
  assign   tlMasterXbar__monitor___address_ok_T_75  =  tlMasterXbar__monitor___address_ok_T_44  |  tlMasterXbar__monitor___address_ok_T_49  ; 
  assign   tlMasterXbar__monitor___address_ok_T_76  =  tlMasterXbar__monitor___address_ok_T_75  |  tlMasterXbar__monitor___address_ok_T_54  ; 
  assign   tlMasterXbar__monitor___address_ok_T_77  =  tlMasterXbar__monitor___address_ok_T_76  |  tlMasterXbar__monitor___address_ok_T_59  ; 
  assign   tlMasterXbar__monitor___address_ok_T_78  =  tlMasterXbar__monitor___address_ok_T_77  |  tlMasterXbar__monitor___address_ok_T_64  ; 
  assign   tlMasterXbar__monitor___address_ok_T_79  =  tlMasterXbar__monitor___address_ok_T_78  |  tlMasterXbar__monitor___address_ok_T_69  ; 
  assign   tlMasterXbar__monitor__address_ok_1  =  tlMasterXbar__monitor___address_ok_T_79  |  tlMasterXbar__monitor___address_ok_T_74  ; 
  assign   tlMasterXbar__monitor___T_1483  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h4; 
  assign   tlMasterXbar__monitor___T_1485  =  tlMasterXbar__monitor__address_ok_1  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1488  =  tlMasterXbar__monitor__source_ok_2  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1490  =  tlMasterXbar__monitor__io_in_c_bits_size  >=4'h3; 
  assign   tlMasterXbar__monitor___T_1492  =  tlMasterXbar__monitor___T_1490  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1495  =  tlMasterXbar__monitor__is_aligned_2  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1497  =  tlMasterXbar__monitor__io_in_c_bits_param  <=3'h5; 
  assign   tlMasterXbar__monitor___T_1499  =  tlMasterXbar__monitor___T_1497  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1505  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h5; 
  assign   tlMasterXbar__monitor___T_1523  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h6; 
  assign   tlMasterXbar__monitor___T_1525  =  tlMasterXbar__monitor__io_in_c_bits_size  <=4'hc; 
  assign   tlMasterXbar__monitor___T_1530  =  tlMasterXbar__monitor___T_1525  &  tlMasterXbar__monitor__source_ok_2  ; 
  assign   tlMasterXbar__monitor___T_1563  =  tlMasterXbar__monitor___address_ok_T_59  |  tlMasterXbar__monitor___address_ok_T_44  ; 
  assign   tlMasterXbar__monitor___T_1564  =  tlMasterXbar__monitor___T_1563  |  tlMasterXbar__monitor___address_ok_T_64  ; 
  assign   tlMasterXbar__monitor___T_1565  =  tlMasterXbar__monitor___T_1564  |  tlMasterXbar__monitor___address_ok_T_54  ; 
  assign   tlMasterXbar__monitor___T_1566  =  tlMasterXbar__monitor___T_1565  |  tlMasterXbar__monitor___address_ok_T_49  ; 
  assign   tlMasterXbar__monitor___T_1567  =  tlMasterXbar__monitor___T_1566  |  tlMasterXbar__monitor___address_ok_T_74  ; 
  assign   tlMasterXbar__monitor___T_1570  =  tlMasterXbar__monitor__io_in_c_bits_size  <=4'h6; 
  assign   tlMasterXbar__monitor___T_1578  =  tlMasterXbar__monitor___T_1570  &  tlMasterXbar__monitor___address_ok_T_69  ; 
  assign   tlMasterXbar__monitor___T_1581  =  tlMasterXbar__monitor___T_1530  &  tlMasterXbar__monitor___T_1578  ; 
  assign   tlMasterXbar__monitor___T_1583  =  tlMasterXbar__monitor___T_1581  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1587  =4'h6==  tlMasterXbar__monitor__io_in_c_bits_size  ; 
  assign   tlMasterXbar__monitor___T_1588  =~  tlMasterXbar__monitor__io_in_c_bits_source  &  tlMasterXbar__monitor___T_1587  ; 
  assign   tlMasterXbar__monitor___T_1635  =  tlMasterXbar__monitor___T_1567  |  tlMasterXbar__monitor___address_ok_T_69  ; 
  assign   tlMasterXbar__monitor___T_1636  =  tlMasterXbar__monitor___T_1525  &  tlMasterXbar__monitor___T_1635  ; 
  assign   tlMasterXbar__monitor___T_1638  =  tlMasterXbar__monitor___T_1588  &  tlMasterXbar__monitor___T_1636  ; 
  assign   tlMasterXbar__monitor___T_1640  =  tlMasterXbar__monitor___T_1638  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1660  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h7; 
  assign   tlMasterXbar__monitor___T_1793  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h0; 
  assign   tlMasterXbar__monitor___T_1803  =  tlMasterXbar__monitor__io_in_c_bits_param  ==3'h0; 
  assign   tlMasterXbar__monitor___T_1805  =  tlMasterXbar__monitor___T_1803  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1811  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h1; 
  assign   tlMasterXbar__monitor___T_1825  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h2; 
  assign   tlMasterXbar__monitor___a_first_T  =  tlMasterXbar__monitor__io_in_a_ready  &  tlMasterXbar__monitor__io_in_a_valid  ; 
  assign   tlMasterXbar__monitor__a_first_beats1_decode  =  tlMasterXbar__monitor__is_aligned_mask  [11:3]; 
  assign   tlMasterXbar__monitor__a_first_beats1_opdata  =~  tlMasterXbar__monitor__io_in_a_bits_opcode  [2]; 
  assign   tlMasterXbar__monitor__a_first_counter1  =  tlMasterXbar__monitor__a_first_counter  -9'h1; 
  assign   tlMasterXbar__monitor__a_first  =  tlMasterXbar__monitor__a_first_counter  ==9'h0; 
  assign   tlMasterXbar__monitor___T_1847  =  tlMasterXbar__monitor__io_in_a_valid  &~  tlMasterXbar__monitor__a_first  ; 
  assign   tlMasterXbar__monitor___T_1848  =  tlMasterXbar__monitor__io_in_a_bits_opcode  ==  tlMasterXbar__monitor__opcode  ; 
  assign   tlMasterXbar__monitor___T_1850  =  tlMasterXbar__monitor___T_1848  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1852  =  tlMasterXbar__monitor__io_in_a_bits_param  ==  tlMasterXbar__monitor__param  ; 
  assign   tlMasterXbar__monitor___T_1854  =  tlMasterXbar__monitor___T_1852  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1856  =  tlMasterXbar__monitor__io_in_a_bits_size  ==  tlMasterXbar__monitor__size  ; 
  assign   tlMasterXbar__monitor___T_1858  =  tlMasterXbar__monitor___T_1856  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1860  =  tlMasterXbar__monitor__io_in_a_bits_source  ==  tlMasterXbar__monitor__source  ; 
  assign   tlMasterXbar__monitor___T_1862  =  tlMasterXbar__monitor___T_1860  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1864  =  tlMasterXbar__monitor__io_in_a_bits_address  ==  tlMasterXbar__monitor__address  ; 
  assign   tlMasterXbar__monitor___T_1866  =  tlMasterXbar__monitor___T_1864  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1869  =  tlMasterXbar__monitor___a_first_T  &  tlMasterXbar__monitor__a_first  ; 
  assign   tlMasterXbar__monitor___d_first_T  =  tlMasterXbar__monitor__io_in_d_ready  &  tlMasterXbar__monitor__io_in_d_valid  ; 
  assign   tlMasterXbar__monitor___d_first_beats1_decode_T_1  =27'hfff<<  tlMasterXbar__monitor__io_in_d_bits_size  ; 
  assign   tlMasterXbar__monitor__d_first_beats1_decode  =~  tlMasterXbar__monitor___d_first_beats1_decode_T_1  [11:3]; 
  assign   tlMasterXbar__monitor__d_first_beats1_opdata  =  tlMasterXbar__monitor__io_in_d_bits_opcode  [0]; 
  assign   tlMasterXbar__monitor__d_first_counter1  =  tlMasterXbar__monitor__d_first_counter  -9'h1; 
  assign   tlMasterXbar__monitor__d_first  =  tlMasterXbar__monitor__d_first_counter  ==9'h0; 
  assign   tlMasterXbar__monitor___T_1871  =  tlMasterXbar__monitor__io_in_d_valid  &~  tlMasterXbar__monitor__d_first  ; 
  assign   tlMasterXbar__monitor___T_1872  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor__opcode_1  ; 
  assign   tlMasterXbar__monitor___T_1874  =  tlMasterXbar__monitor___T_1872  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1876  =  tlMasterXbar__monitor__io_in_d_bits_param  ==  tlMasterXbar__monitor__param_1  ; 
  assign   tlMasterXbar__monitor___T_1878  =  tlMasterXbar__monitor___T_1876  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1880  =  tlMasterXbar__monitor__io_in_d_bits_size  ==  tlMasterXbar__monitor__size_1  ; 
  assign   tlMasterXbar__monitor___T_1882  =  tlMasterXbar__monitor___T_1880  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1884  =  tlMasterXbar__monitor__io_in_d_bits_source  ==  tlMasterXbar__monitor__source_1  ; 
  assign   tlMasterXbar__monitor___T_1886  =  tlMasterXbar__monitor___T_1884  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1888  =  tlMasterXbar__monitor__io_in_d_bits_sink  ==  tlMasterXbar__monitor__sink  ; 
  assign   tlMasterXbar__monitor___T_1890  =  tlMasterXbar__monitor___T_1888  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1892  =  tlMasterXbar__monitor__io_in_d_bits_denied  ==  tlMasterXbar__monitor__denied  ; 
  assign   tlMasterXbar__monitor___T_1894  =  tlMasterXbar__monitor___T_1892  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1897  =  tlMasterXbar__monitor___d_first_T  &  tlMasterXbar__monitor__d_first  ; 
  assign   tlMasterXbar__monitor__b_first_done  =  tlMasterXbar__monitor__io_in_b_ready  &  tlMasterXbar__monitor__io_in_b_valid  ; 
  assign   tlMasterXbar__monitor__b_first_counter1  =  tlMasterXbar__monitor__b_first_counter  -9'h1; 
  assign   tlMasterXbar__monitor__b_first  =  tlMasterXbar__monitor__b_first_counter  ==9'h0; 
  assign   tlMasterXbar__monitor___T_1899  =  tlMasterXbar__monitor__io_in_b_valid  &~  tlMasterXbar__monitor__b_first  ; 
  assign   tlMasterXbar__monitor___T_1900  =  tlMasterXbar__monitor__io_in_b_bits_opcode  ==  tlMasterXbar__monitor__opcode_2  ; 
  assign   tlMasterXbar__monitor___T_1902  =  tlMasterXbar__monitor___T_1900  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1904  =  tlMasterXbar__monitor__io_in_b_bits_param  ==  tlMasterXbar__monitor__param_2  ; 
  assign   tlMasterXbar__monitor___T_1906  =  tlMasterXbar__monitor___T_1904  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1908  =  tlMasterXbar__monitor__io_in_b_bits_size  ==  tlMasterXbar__monitor__size_2  ; 
  assign   tlMasterXbar__monitor___T_1910  =  tlMasterXbar__monitor___T_1908  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1912  =  tlMasterXbar__monitor__io_in_b_bits_source  ==  tlMasterXbar__monitor__source_2  ; 
  assign   tlMasterXbar__monitor___T_1914  =  tlMasterXbar__monitor___T_1912  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1916  =  tlMasterXbar__monitor__io_in_b_bits_address  ==  tlMasterXbar__monitor__address_1  ; 
  assign   tlMasterXbar__monitor___T_1918  =  tlMasterXbar__monitor___T_1916  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1921  =  tlMasterXbar__monitor__b_first_done  &  tlMasterXbar__monitor__b_first  ; 
  assign   tlMasterXbar__monitor___c_first_T  =  tlMasterXbar__monitor__io_in_c_ready  &  tlMasterXbar__monitor__io_in_c_valid  ; 
  assign   tlMasterXbar__monitor__c_first_beats1_decode  =  tlMasterXbar__monitor__is_aligned_mask_2  [11:3]; 
  assign   tlMasterXbar__monitor__c_first_beats1_opdata  =  tlMasterXbar__monitor__io_in_c_bits_opcode  [0]; 
  assign   tlMasterXbar__monitor__c_first_counter1  =  tlMasterXbar__monitor__c_first_counter  -9'h1; 
  assign   tlMasterXbar__monitor__c_first  =  tlMasterXbar__monitor__c_first_counter  ==9'h0; 
  assign   tlMasterXbar__monitor___T_1923  =  tlMasterXbar__monitor__io_in_c_valid  &~  tlMasterXbar__monitor__c_first  ; 
  assign   tlMasterXbar__monitor___T_1924  =  tlMasterXbar__monitor__io_in_c_bits_opcode  ==  tlMasterXbar__monitor__opcode_3  ; 
  assign   tlMasterXbar__monitor___T_1926  =  tlMasterXbar__monitor___T_1924  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1928  =  tlMasterXbar__monitor__io_in_c_bits_param  ==  tlMasterXbar__monitor__param_3  ; 
  assign   tlMasterXbar__monitor___T_1930  =  tlMasterXbar__monitor___T_1928  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1932  =  tlMasterXbar__monitor__io_in_c_bits_size  ==  tlMasterXbar__monitor__size_3  ; 
  assign   tlMasterXbar__monitor___T_1934  =  tlMasterXbar__monitor___T_1932  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1936  =  tlMasterXbar__monitor__io_in_c_bits_source  ==  tlMasterXbar__monitor__source_3  ; 
  assign   tlMasterXbar__monitor___T_1938  =  tlMasterXbar__monitor___T_1936  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1940  =  tlMasterXbar__monitor__io_in_c_bits_address  ==  tlMasterXbar__monitor__address_2  ; 
  assign   tlMasterXbar__monitor___T_1942  =  tlMasterXbar__monitor___T_1940  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1945  =  tlMasterXbar__monitor___c_first_T  &  tlMasterXbar__monitor__c_first  ; 
  assign   tlMasterXbar__monitor__a_first_counter1_1  =  tlMasterXbar__monitor__a_first_counter_1  -9'h1; 
  assign   tlMasterXbar__monitor__a_first_1  =  tlMasterXbar__monitor__a_first_counter_1  ==9'h0; 
  assign   tlMasterXbar__monitor__d_first_counter1_1  =  tlMasterXbar__monitor__d_first_counter_1  -9'h1; 
  assign   tlMasterXbar__monitor__d_first_1  =  tlMasterXbar__monitor__d_first_counter_1  ==9'h0; 
  assign   tlMasterXbar__monitor___GEN_89  ={  tlMasterXbar__monitor__io_in_d_bits_source  ,2'h0}; 
  assign   tlMasterXbar__monitor___a_opcode_lookup_T  ={1'b0,  tlMasterXbar__monitor___GEN_89  }; 
  assign   tlMasterXbar__monitor___a_opcode_lookup_T_1  =  tlMasterXbar__monitor__inflight_opcodes  >>  tlMasterXbar__monitor___a_opcode_lookup_T  ; 
  assign   tlMasterXbar__monitor___a_opcode_lookup_T_5  =16'h10-16'h1; 
  assign   tlMasterXbar__monitor___GEN_90  ={8'b0,  tlMasterXbar__monitor___a_opcode_lookup_T_1  }; 
  assign   tlMasterXbar__monitor___a_opcode_lookup_T_6  =  tlMasterXbar__monitor___GEN_90  &  tlMasterXbar__monitor___a_opcode_lookup_T_5  ; 
  assign   tlMasterXbar__monitor___a_opcode_lookup_T_7  ={1'b0,  tlMasterXbar__monitor___a_opcode_lookup_T_6  [15:1]}; 
  assign   tlMasterXbar__monitor___a_size_lookup_T  ={  tlMasterXbar__monitor__io_in_d_bits_source  ,3'h0}; 
  assign   tlMasterXbar__monitor___a_size_lookup_T_1  =  tlMasterXbar__monitor__inflight_sizes  >>  tlMasterXbar__monitor___a_size_lookup_T  ; 
  assign   tlMasterXbar__monitor___a_size_lookup_T_5  =16'h100-16'h1; 
  assign   tlMasterXbar__monitor___a_size_lookup_T_6  =  tlMasterXbar__monitor___a_size_lookup_T_1  &  tlMasterXbar__monitor___a_size_lookup_T_5  ; 
  assign   tlMasterXbar__monitor___a_size_lookup_T_7  ={1'b0,  tlMasterXbar__monitor___a_size_lookup_T_6  [15:1]}; 
  assign   tlMasterXbar__monitor___T_1946  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__a_first_1  ; 
  assign   tlMasterXbar__monitor___a_set_wo_ready_T  =2'h1<<  tlMasterXbar__monitor__io_in_a_bits_source  ; 
  assign   tlMasterXbar__monitor__a_set_wo_ready  =  tlMasterXbar__monitor___T_1946   ?   tlMasterXbar__monitor___a_set_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___T_1949  =  tlMasterXbar__monitor___a_first_T  &  tlMasterXbar__monitor__a_first_1  ; 
  assign   tlMasterXbar__monitor___a_opcodes_set_interm_T  ={  tlMasterXbar__monitor__io_in_a_bits_opcode  ,1'h0}; 
  assign   tlMasterXbar__monitor___a_opcodes_set_interm_T_1  =  tlMasterXbar__monitor___a_opcodes_set_interm_T  |4'h1; 
  assign   tlMasterXbar__monitor___a_sizes_set_interm_T  ={  tlMasterXbar__monitor__io_in_a_bits_size  ,1'h0}; 
  assign   tlMasterXbar__monitor___a_sizes_set_interm_T_1  =  tlMasterXbar__monitor___a_sizes_set_interm_T  |5'h1; 
  assign   tlMasterXbar__monitor___GEN_93  ={  tlMasterXbar__monitor__io_in_a_bits_source  ,2'h0}; 
  assign   tlMasterXbar__monitor___a_opcodes_set_T  ={1'b0,  tlMasterXbar__monitor___GEN_93  }; 
  assign   tlMasterXbar__monitor__a_opcodes_set_interm  =  tlMasterXbar__monitor___T_1949   ?   tlMasterXbar__monitor___a_opcodes_set_interm_T_1  :4'h0; 
  assign   tlMasterXbar__monitor___GEN_94  ={15'b0,  tlMasterXbar__monitor__a_opcodes_set_interm  }; 
  assign   tlMasterXbar__monitor___a_opcodes_set_T_1  =  tlMasterXbar__monitor___GEN_94  <<  tlMasterXbar__monitor___a_opcodes_set_T  ; 
  assign   tlMasterXbar__monitor___a_sizes_set_T  ={  tlMasterXbar__monitor__io_in_a_bits_source  ,3'h0}; 
  assign   tlMasterXbar__monitor__a_sizes_set_interm  =  tlMasterXbar__monitor___T_1949   ?   tlMasterXbar__monitor___a_sizes_set_interm_T_1  :5'h0; 
  assign   tlMasterXbar__monitor___GEN_95  ={15'b0,  tlMasterXbar__monitor__a_sizes_set_interm  }; 
  assign   tlMasterXbar__monitor___a_sizes_set_T_1  =  tlMasterXbar__monitor___GEN_95  <<  tlMasterXbar__monitor___a_sizes_set_T  ; 
  assign   tlMasterXbar__monitor___T_1951  =  tlMasterXbar__monitor__inflight  >>  tlMasterXbar__monitor__io_in_a_bits_source  ; 
  assign   tlMasterXbar__monitor___T_1955  =~  tlMasterXbar__monitor___T_1951  [0]|  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__a_set  =  tlMasterXbar__monitor___T_1949   ?   tlMasterXbar__monitor___a_set_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___GEN_31  =  tlMasterXbar__monitor___T_1949   ?   tlMasterXbar__monitor___a_opcodes_set_T_1  :19'h0; 
  assign   tlMasterXbar__monitor___GEN_32  =  tlMasterXbar__monitor___T_1949   ?   tlMasterXbar__monitor___a_sizes_set_T_1  :20'h0; 
  assign   tlMasterXbar__monitor___T_1957  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__d_first_1  ; 
  assign   tlMasterXbar__monitor___T_1960  =  tlMasterXbar__monitor___T_1957  &~  tlMasterXbar__monitor___T_807  ; 
  assign   tlMasterXbar__monitor___d_clr_wo_ready_T  =2'h1<<  tlMasterXbar__monitor__io_in_d_bits_source  ; 
  assign   tlMasterXbar__monitor__d_clr_wo_ready  =  tlMasterXbar__monitor___T_1960   ?   tlMasterXbar__monitor___d_clr_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___T_1962  =  tlMasterXbar__monitor___d_first_T  &  tlMasterXbar__monitor__d_first_1  ; 
  assign   tlMasterXbar__monitor___T_1965  =  tlMasterXbar__monitor___T_1962  &~  tlMasterXbar__monitor___T_807  ; 
  assign   tlMasterXbar__monitor___GEN_97  ={15'b0,  tlMasterXbar__monitor___a_opcode_lookup_T_5  }; 
  assign   tlMasterXbar__monitor___d_opcodes_clr_T_5  =  tlMasterXbar__monitor___GEN_97  <<  tlMasterXbar__monitor___a_opcode_lookup_T  ; 
  assign   tlMasterXbar__monitor___GEN_98  ={15'b0,  tlMasterXbar__monitor___a_size_lookup_T_5  }; 
  assign   tlMasterXbar__monitor___d_sizes_clr_T_5  =  tlMasterXbar__monitor___GEN_98  <<  tlMasterXbar__monitor___a_size_lookup_T  ; 
  assign   tlMasterXbar__monitor__d_clr  =  tlMasterXbar__monitor___T_1965   ?   tlMasterXbar__monitor___d_clr_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___GEN_35  =  tlMasterXbar__monitor___T_1965   ?   tlMasterXbar__monitor___d_opcodes_clr_T_5  :31'h0; 
  assign   tlMasterXbar__monitor___GEN_36  =  tlMasterXbar__monitor___T_1965   ?   tlMasterXbar__monitor___d_sizes_clr_T_5  :31'h0; 
  assign   tlMasterXbar__monitor___same_cycle_resp_T_2  =  tlMasterXbar__monitor__io_in_a_bits_source  ==  tlMasterXbar__monitor__io_in_d_bits_source  ; 
  assign   tlMasterXbar__monitor__same_cycle_resp  =  tlMasterXbar__monitor___T_1946  &  tlMasterXbar__monitor___same_cycle_resp_T_2  ; 
  assign   tlMasterXbar__monitor___T_1970  =  tlMasterXbar__monitor__inflight  >>  tlMasterXbar__monitor__io_in_d_bits_source  ; 
  assign   tlMasterXbar__monitor___T_1972  =  tlMasterXbar__monitor___T_1970  [0]|  tlMasterXbar__monitor__same_cycle_resp  ; 
  assign   tlMasterXbar__monitor___T_1974  =  tlMasterXbar__monitor___T_1972  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___GEN_39  =3'h2==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h1:3'h0; 
  assign   tlMasterXbar__monitor___GEN_40  =3'h3==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h1:  tlMasterXbar__monitor___GEN_39  ; 
  assign   tlMasterXbar__monitor___GEN_41  =3'h4==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h1:  tlMasterXbar__monitor___GEN_40  ; 
  assign   tlMasterXbar__monitor___GEN_42  =3'h5==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h2:  tlMasterXbar__monitor___GEN_41  ; 
  assign   tlMasterXbar__monitor___GEN_43  =3'h6==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h4:  tlMasterXbar__monitor___GEN_42  ; 
  assign   tlMasterXbar__monitor___GEN_44  =3'h7==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h4:  tlMasterXbar__monitor___GEN_43  ; 
  assign   tlMasterXbar__monitor___T_1976  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor___GEN_44  ; 
  assign   tlMasterXbar__monitor___GEN_51  =3'h6==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h5:  tlMasterXbar__monitor___GEN_42  ; 
  assign   tlMasterXbar__monitor___GEN_52  =3'h7==  tlMasterXbar__monitor__io_in_a_bits_opcode   ? 3'h4:  tlMasterXbar__monitor___GEN_51  ; 
  assign   tlMasterXbar__monitor___T_1977  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor___GEN_52  ; 
  assign   tlMasterXbar__monitor___T_1978  =  tlMasterXbar__monitor___T_1976  |  tlMasterXbar__monitor___T_1977  ; 
  assign   tlMasterXbar__monitor___T_1980  =  tlMasterXbar__monitor___T_1978  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1982  =  tlMasterXbar__monitor__io_in_a_bits_size  ==  tlMasterXbar__monitor__io_in_d_bits_size  ; 
  assign   tlMasterXbar__monitor___T_1984  =  tlMasterXbar__monitor___T_1982  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__a_opcode_lookup  =  tlMasterXbar__monitor___a_opcode_lookup_T_7  [3:0]; 
  assign   tlMasterXbar__monitor___GEN_55  =3'h2==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h1:3'h0; 
  assign   tlMasterXbar__monitor___GEN_56  =3'h3==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h1:  tlMasterXbar__monitor___GEN_55  ; 
  assign   tlMasterXbar__monitor___GEN_57  =3'h4==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h1:  tlMasterXbar__monitor___GEN_56  ; 
  assign   tlMasterXbar__monitor___GEN_58  =3'h5==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h2:  tlMasterXbar__monitor___GEN_57  ; 
  assign   tlMasterXbar__monitor___GEN_59  =3'h6==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h4:  tlMasterXbar__monitor___GEN_58  ; 
  assign   tlMasterXbar__monitor___GEN_60  =3'h7==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h4:  tlMasterXbar__monitor___GEN_59  ; 
  assign   tlMasterXbar__monitor___T_1987  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor___GEN_60  ; 
  assign   tlMasterXbar__monitor___GEN_67  =3'h6==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h5:  tlMasterXbar__monitor___GEN_58  ; 
  assign   tlMasterXbar__monitor___GEN_68  =3'h7==  tlMasterXbar__monitor__a_opcode_lookup  [2:0] ? 3'h4:  tlMasterXbar__monitor___GEN_67  ; 
  assign   tlMasterXbar__monitor___T_1989  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor___GEN_68  ; 
  assign   tlMasterXbar__monitor___T_1990  =  tlMasterXbar__monitor___T_1987  |  tlMasterXbar__monitor___T_1989  ; 
  assign   tlMasterXbar__monitor___T_1992  =  tlMasterXbar__monitor___T_1990  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__a_size_lookup  =  tlMasterXbar__monitor___a_size_lookup_T_7  [7:0]; 
  assign   tlMasterXbar__monitor___GEN_99  ={4'b0,  tlMasterXbar__monitor__io_in_d_bits_size  }; 
  assign   tlMasterXbar__monitor___T_1994  =  tlMasterXbar__monitor___GEN_99  ==  tlMasterXbar__monitor__a_size_lookup  ; 
  assign   tlMasterXbar__monitor___T_1996  =  tlMasterXbar__monitor___T_1994  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_1999  =  tlMasterXbar__monitor___T_1957  &  tlMasterXbar__monitor__a_first_1  ; 
  assign   tlMasterXbar__monitor___T_2000  =  tlMasterXbar__monitor___T_1999  &  tlMasterXbar__monitor__io_in_a_valid  ; 
  assign   tlMasterXbar__monitor___T_2002  =  tlMasterXbar__monitor___T_2000  &  tlMasterXbar__monitor___same_cycle_resp_T_2  ; 
  assign   tlMasterXbar__monitor___T_2004  =  tlMasterXbar__monitor___T_2002  &~  tlMasterXbar__monitor___T_807  ; 
  assign   tlMasterXbar__monitor___T_2006  =~  tlMasterXbar__monitor__io_in_d_ready  |  tlMasterXbar__monitor__io_in_a_ready  ; 
  assign   tlMasterXbar__monitor___T_2008  =  tlMasterXbar__monitor___T_2006  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_2010  =  tlMasterXbar__monitor__a_set_wo_ready  !=  tlMasterXbar__monitor__d_clr_wo_ready  ; 
  assign   tlMasterXbar__monitor___T_2011  =|  tlMasterXbar__monitor__a_set_wo_ready  ; 
  assign   tlMasterXbar__monitor___T_2013  =  tlMasterXbar__monitor___T_2010  |~  tlMasterXbar__monitor___T_2011  ; 
  assign   tlMasterXbar__monitor___T_2015  =  tlMasterXbar__monitor___T_2013  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___inflight_T  =  tlMasterXbar__monitor__inflight  |  tlMasterXbar__monitor__a_set  ; 
  assign   tlMasterXbar__monitor___inflight_T_2  =  tlMasterXbar__monitor___inflight_T  &~  tlMasterXbar__monitor__d_clr  ; 
  assign   tlMasterXbar__monitor__a_opcodes_set  =  tlMasterXbar__monitor___GEN_31  [7:0]; 
  assign   tlMasterXbar__monitor___inflight_opcodes_T  =  tlMasterXbar__monitor__inflight_opcodes  |  tlMasterXbar__monitor__a_opcodes_set  ; 
  assign   tlMasterXbar__monitor__d_opcodes_clr  =  tlMasterXbar__monitor___GEN_35  [7:0]; 
  assign   tlMasterXbar__monitor___inflight_opcodes_T_2  =  tlMasterXbar__monitor___inflight_opcodes_T  &~  tlMasterXbar__monitor__d_opcodes_clr  ; 
  assign   tlMasterXbar__monitor__a_sizes_set  =  tlMasterXbar__monitor___GEN_32  [15:0]; 
  assign   tlMasterXbar__monitor___inflight_sizes_T  =  tlMasterXbar__monitor__inflight_sizes  |  tlMasterXbar__monitor__a_sizes_set  ; 
  assign   tlMasterXbar__monitor__d_sizes_clr  =  tlMasterXbar__monitor___GEN_36  [15:0]; 
  assign   tlMasterXbar__monitor___inflight_sizes_T_2  =  tlMasterXbar__monitor___inflight_sizes_T  &~  tlMasterXbar__monitor__d_sizes_clr  ; 
  assign   tlMasterXbar__monitor___T_2017  =|  tlMasterXbar__monitor__inflight  ; 
  assign   tlMasterXbar__monitor___T_2019  =  tlMasterXbar__monitor__plusarg_reader_out  ==32'h0; 
  assign   tlMasterXbar__monitor___T_2020  =~  tlMasterXbar__monitor___T_2017  |  tlMasterXbar__monitor___T_2019  ; 
  assign   tlMasterXbar__monitor___T_2021  =  tlMasterXbar__monitor__watchdog  <  tlMasterXbar__monitor__plusarg_reader_out  ; 
  assign   tlMasterXbar__monitor___T_2022  =  tlMasterXbar__monitor___T_2020  |  tlMasterXbar__monitor___T_2021  ; 
  assign   tlMasterXbar__monitor___T_2024  =  tlMasterXbar__monitor___T_2022  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___watchdog_T_1  =  tlMasterXbar__monitor__watchdog  +32'h1; 
  assign   tlMasterXbar__monitor___T_2028  =  tlMasterXbar__monitor___a_first_T  |  tlMasterXbar__monitor___d_first_T  ; 
  assign   tlMasterXbar__monitor__c_first_counter1_1  =  tlMasterXbar__monitor__c_first_counter_1  -9'h1; 
  assign   tlMasterXbar__monitor__c_first_1  =  tlMasterXbar__monitor__c_first_counter_1  ==9'h0; 
  assign   tlMasterXbar__monitor__d_first_counter1_2  =  tlMasterXbar__monitor__d_first_counter_2  -9'h1; 
  assign   tlMasterXbar__monitor__d_first_2  =  tlMasterXbar__monitor__d_first_counter_2  ==9'h0; 
  assign   tlMasterXbar__monitor___c_size_lookup_T_1  =  tlMasterXbar__monitor__inflight_sizes_1  >>  tlMasterXbar__monitor___a_size_lookup_T  ; 
  assign   tlMasterXbar__monitor___c_size_lookup_T_6  =  tlMasterXbar__monitor___c_size_lookup_T_1  &  tlMasterXbar__monitor___a_size_lookup_T_5  ; 
  assign   tlMasterXbar__monitor___c_size_lookup_T_7  ={1'b0,  tlMasterXbar__monitor___c_size_lookup_T_6  [15:1]}; 
  assign   tlMasterXbar__monitor___T_2029  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__c_first_1  ; 
  assign   tlMasterXbar__monitor___T_2032  =  tlMasterXbar__monitor__io_in_c_bits_opcode  [2]&  tlMasterXbar__monitor__io_in_c_bits_opcode  [1]; 
  assign   tlMasterXbar__monitor___T_2033  =  tlMasterXbar__monitor___T_2029  &  tlMasterXbar__monitor___T_2032  ; 
  assign   tlMasterXbar__monitor___c_set_wo_ready_T  =2'h1<<  tlMasterXbar__monitor__io_in_c_bits_source  ; 
  assign   tlMasterXbar__monitor__c_set_wo_ready  =  tlMasterXbar__monitor___T_2033   ?   tlMasterXbar__monitor___c_set_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___T_2035  =  tlMasterXbar__monitor___c_first_T  &  tlMasterXbar__monitor__c_first_1  ; 
  assign   tlMasterXbar__monitor___T_2039  =  tlMasterXbar__monitor___T_2035  &  tlMasterXbar__monitor___T_2032  ; 
  assign   tlMasterXbar__monitor___c_sizes_set_interm_T  ={  tlMasterXbar__monitor__io_in_c_bits_size  ,1'h0}; 
  assign   tlMasterXbar__monitor___c_sizes_set_interm_T_1  =  tlMasterXbar__monitor___c_sizes_set_interm_T  |5'h1; 
  assign   tlMasterXbar__monitor___c_sizes_set_T  ={  tlMasterXbar__monitor__io_in_c_bits_source  ,3'h0}; 
  assign   tlMasterXbar__monitor__c_sizes_set_interm  =  tlMasterXbar__monitor___T_2039   ?   tlMasterXbar__monitor___c_sizes_set_interm_T_1  :5'h0; 
  assign   tlMasterXbar__monitor___GEN_106  ={15'b0,  tlMasterXbar__monitor__c_sizes_set_interm  }; 
  assign   tlMasterXbar__monitor___c_sizes_set_T_1  =  tlMasterXbar__monitor___GEN_106  <<  tlMasterXbar__monitor___c_sizes_set_T  ; 
  assign   tlMasterXbar__monitor___T_2040  =  tlMasterXbar__monitor__inflight_1  >>  tlMasterXbar__monitor__io_in_c_bits_source  ; 
  assign   tlMasterXbar__monitor___T_2044  =~  tlMasterXbar__monitor___T_2040  [0]|  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__c_set  =  tlMasterXbar__monitor___T_2039   ?   tlMasterXbar__monitor___c_set_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___GEN_77  =  tlMasterXbar__monitor___T_2039   ?   tlMasterXbar__monitor___c_sizes_set_T_1  :20'h0; 
  assign   tlMasterXbar__monitor___T_2046  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__d_first_2  ; 
  assign   tlMasterXbar__monitor___T_2048  =  tlMasterXbar__monitor___T_2046  &  tlMasterXbar__monitor___T_807  ; 
  assign   tlMasterXbar__monitor__d_clr_wo_ready_1  =  tlMasterXbar__monitor___T_2048   ?   tlMasterXbar__monitor___d_clr_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___T_2050  =  tlMasterXbar__monitor___d_first_T  &  tlMasterXbar__monitor__d_first_2  ; 
  assign   tlMasterXbar__monitor___T_2052  =  tlMasterXbar__monitor___T_2050  &  tlMasterXbar__monitor___T_807  ; 
  assign   tlMasterXbar__monitor__d_clr_1  =  tlMasterXbar__monitor___T_2052   ?   tlMasterXbar__monitor___d_clr_wo_ready_T  :2'h0; 
  assign   tlMasterXbar__monitor___GEN_81  =  tlMasterXbar__monitor___T_2052   ?   tlMasterXbar__monitor___d_sizes_clr_T_5  :31'h0; 
  assign   tlMasterXbar__monitor___same_cycle_resp_T_8  =  tlMasterXbar__monitor__io_in_c_bits_source  ==  tlMasterXbar__monitor__io_in_d_bits_source  ; 
  assign   tlMasterXbar__monitor__same_cycle_resp_1  =  tlMasterXbar__monitor___T_2033  &  tlMasterXbar__monitor___same_cycle_resp_T_8  ; 
  assign   tlMasterXbar__monitor___T_2056  =  tlMasterXbar__monitor__inflight_1  >>  tlMasterXbar__monitor__io_in_d_bits_source  ; 
  assign   tlMasterXbar__monitor___T_2058  =  tlMasterXbar__monitor___T_2056  [0]|  tlMasterXbar__monitor__same_cycle_resp_1  ; 
  assign   tlMasterXbar__monitor___T_2060  =  tlMasterXbar__monitor___T_2058  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_2062  =  tlMasterXbar__monitor__io_in_d_bits_size  ==  tlMasterXbar__monitor__io_in_c_bits_size  ; 
  assign   tlMasterXbar__monitor___T_2064  =  tlMasterXbar__monitor___T_2062  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__c_size_lookup  =  tlMasterXbar__monitor___c_size_lookup_T_7  [7:0]; 
  assign   tlMasterXbar__monitor___T_2066  =  tlMasterXbar__monitor___GEN_99  ==  tlMasterXbar__monitor__c_size_lookup  ; 
  assign   tlMasterXbar__monitor___T_2068  =  tlMasterXbar__monitor___T_2066  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_2071  =  tlMasterXbar__monitor___T_2046  &  tlMasterXbar__monitor__c_first_1  ; 
  assign   tlMasterXbar__monitor___T_2072  =  tlMasterXbar__monitor___T_2071  &  tlMasterXbar__monitor__io_in_c_valid  ; 
  assign   tlMasterXbar__monitor___T_2074  =  tlMasterXbar__monitor___T_2072  &  tlMasterXbar__monitor___same_cycle_resp_T_8  ; 
  assign   tlMasterXbar__monitor___T_2075  =  tlMasterXbar__monitor___T_2074  &  tlMasterXbar__monitor___T_807  ; 
  assign   tlMasterXbar__monitor___T_2077  =~  tlMasterXbar__monitor__io_in_d_ready  |  tlMasterXbar__monitor__io_in_c_ready  ; 
  assign   tlMasterXbar__monitor___T_2079  =  tlMasterXbar__monitor___T_2077  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___T_2081  =|  tlMasterXbar__monitor__c_set_wo_ready  ; 
  assign   tlMasterXbar__monitor___T_2082  =  tlMasterXbar__monitor__c_set_wo_ready  !=  tlMasterXbar__monitor__d_clr_wo_ready_1  ; 
  assign   tlMasterXbar__monitor___T_2084  =  tlMasterXbar__monitor___T_2082  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___inflight_T_3  =  tlMasterXbar__monitor__inflight_1  |  tlMasterXbar__monitor__c_set  ; 
  assign   tlMasterXbar__monitor___inflight_T_5  =  tlMasterXbar__monitor___inflight_T_3  &~  tlMasterXbar__monitor__d_clr_1  ; 
  assign   tlMasterXbar__monitor__c_sizes_set  =  tlMasterXbar__monitor___GEN_77  [15:0]; 
  assign   tlMasterXbar__monitor___inflight_sizes_T_3  =  tlMasterXbar__monitor__inflight_sizes_1  |  tlMasterXbar__monitor__c_sizes_set  ; 
  assign   tlMasterXbar__monitor__d_sizes_clr_1  =  tlMasterXbar__monitor___GEN_81  [15:0]; 
  assign   tlMasterXbar__monitor___inflight_sizes_T_5  =  tlMasterXbar__monitor___inflight_sizes_T_3  &~  tlMasterXbar__monitor__d_sizes_clr_1  ; 
  assign   tlMasterXbar__monitor___T_2086  =|  tlMasterXbar__monitor__inflight_1  ; 
  assign   tlMasterXbar__monitor___T_2088  =  tlMasterXbar__monitor__plusarg_reader_1_out  ==32'h0; 
  assign   tlMasterXbar__monitor___T_2089  =~  tlMasterXbar__monitor___T_2086  |  tlMasterXbar__monitor___T_2088  ; 
  assign   tlMasterXbar__monitor___T_2090  =  tlMasterXbar__monitor__watchdog_1  <  tlMasterXbar__monitor__plusarg_reader_1_out  ; 
  assign   tlMasterXbar__monitor___T_2091  =  tlMasterXbar__monitor___T_2089  |  tlMasterXbar__monitor___T_2090  ; 
  assign   tlMasterXbar__monitor___T_2093  =  tlMasterXbar__monitor___T_2091  |  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor___watchdog_T_3  =  tlMasterXbar__monitor__watchdog_1  +32'h1; 
  assign   tlMasterXbar__monitor___T_2097  =  tlMasterXbar__monitor___c_first_T  |  tlMasterXbar__monitor___d_first_T  ; 
  assign   tlMasterXbar__monitor__d_first_counter1_3  =  tlMasterXbar__monitor__d_first_counter_3  -9'h1; 
  assign   tlMasterXbar__monitor__d_first_3  =  tlMasterXbar__monitor__d_first_counter_3  ==9'h0; 
  assign   tlMasterXbar__monitor___T_2099  =  tlMasterXbar__monitor___d_first_T  &  tlMasterXbar__monitor__d_first_3  ; 
  assign   tlMasterXbar__monitor___T_2103  =  tlMasterXbar__monitor__io_in_d_bits_opcode  [2]&~  tlMasterXbar__monitor__io_in_d_bits_opcode  [1]; 
  assign   tlMasterXbar__monitor___T_2104  =  tlMasterXbar__monitor___T_2099  &  tlMasterXbar__monitor___T_2103  ; 
  assign   tlMasterXbar__monitor___d_set_T  =4'h1<<  tlMasterXbar__monitor__io_in_d_bits_sink  ; 
  assign   tlMasterXbar__monitor___T_2105  =  tlMasterXbar__monitor__inflight_2  >>  tlMasterXbar__monitor__io_in_d_bits_sink  ; 
  assign   tlMasterXbar__monitor___T_2109  =~  tlMasterXbar__monitor___T_2105  [0]|  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__d_set  =  tlMasterXbar__monitor___T_2104   ?   tlMasterXbar__monitor___d_set_T  :4'h0; 
  assign   tlMasterXbar__monitor___T_2111  =  tlMasterXbar__monitor__io_in_e_ready  &  tlMasterXbar__monitor__io_in_e_valid  ; 
  assign   tlMasterXbar__monitor___e_clr_T  =4'h1<<  tlMasterXbar__monitor__io_in_e_bits_sink  ; 
  assign   tlMasterXbar__monitor___T_2114  =  tlMasterXbar__monitor__d_set  |  tlMasterXbar__monitor__inflight_2  ; 
  assign   tlMasterXbar__monitor___T_2115  =  tlMasterXbar__monitor___T_2114  >>  tlMasterXbar__monitor__io_in_e_bits_sink  ; 
  assign   tlMasterXbar__monitor___T_2118  =  tlMasterXbar__monitor___T_2115  [0]|  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__e_clr  =  tlMasterXbar__monitor___T_2111   ?   tlMasterXbar__monitor___e_clr_T  :4'h0; 
  assign   tlMasterXbar__monitor___inflight_T_6  =  tlMasterXbar__monitor__inflight_2  |  tlMasterXbar__monitor__d_set  ; 
  assign   tlMasterXbar__monitor___inflight_T_8  =  tlMasterXbar__monitor___inflight_T_6  &~  tlMasterXbar__monitor__e_clr  ; 
  assign   tlMasterXbar__monitor___GEN_111  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_24  ; 
  assign   tlMasterXbar__monitor___GEN_125  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_166  ; 
  assign   tlMasterXbar__monitor___GEN_141  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_312  ; 
  assign   tlMasterXbar__monitor___GEN_153  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_397  ; 
  assign   tlMasterXbar__monitor___GEN_163  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_483  ; 
  assign   tlMasterXbar__monitor___GEN_173  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_571  ; 
  assign   tlMasterXbar__monitor___GEN_183  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_647  ; 
  assign   tlMasterXbar__monitor___GEN_193  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor___T_723  ; 
  assign   tlMasterXbar__monitor___GEN_203  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor___T_807  ; 
  assign   tlMasterXbar__monitor___GEN_213  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor___T_827  ; 
  assign   tlMasterXbar__monitor___GEN_223  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor___T_855  ; 
  assign   tlMasterXbar__monitor___GEN_233  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor___T_884  ; 
  assign   tlMasterXbar__monitor___GEN_239  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor___T_901  ; 
  assign   tlMasterXbar__monitor___GEN_245  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor___T_919  ; 
  assign   tlMasterXbar__monitor___GEN_251  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor___T_960  ; 
  assign   tlMasterXbar__monitor___GEN_265  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor___T_1039  ; 
  assign   tlMasterXbar__monitor___GEN_279  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor___T_1112  ; 
  assign   tlMasterXbar__monitor___GEN_291  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor___T_1181  ; 
  assign   tlMasterXbar__monitor___GEN_303  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor___T_1252  ; 
  assign   tlMasterXbar__monitor___GEN_313  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor___T_1321  ; 
  assign   tlMasterXbar__monitor___GEN_323  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor___T_1390  ; 
  assign   tlMasterXbar__monitor___GEN_335  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor___T_1483  ; 
  assign   tlMasterXbar__monitor___GEN_345  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor___T_1505  ; 
  assign   tlMasterXbar__monitor___GEN_355  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor___T_1523  ; 
  assign   tlMasterXbar__monitor___GEN_367  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor___T_1660  ; 
  assign   tlMasterXbar__monitor___GEN_379  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor___T_1793  ; 
  assign   tlMasterXbar__monitor___GEN_387  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor___T_1811  ; 
  assign   tlMasterXbar__monitor___GEN_395  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor___T_1825  ; 
  assign   tlMasterXbar__monitor___GEN_403  =  tlMasterXbar__monitor___T_1960  &  tlMasterXbar__monitor__same_cycle_resp  ; 
  assign   tlMasterXbar__monitor___GEN_408  =  tlMasterXbar__monitor___T_1960  &~  tlMasterXbar__monitor__same_cycle_resp  ; 
  assign   tlMasterXbar__monitor___GEN_415  =  tlMasterXbar__monitor___T_2048  &  tlMasterXbar__monitor__same_cycle_resp_1  ; 
  assign   tlMasterXbar__monitor___GEN_418  =  tlMasterXbar__monitor___T_2048  &~  tlMasterXbar__monitor__same_cycle_resp_1  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_covSum  =30'h0; 
  assign   tlMasterXbar__monitor__io_covSum  =  tlMasterXbar__monitor__TLMonitor_23_covSum  ; 
  assign   tlMasterXbar__monitor__stopEn0  =  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_84  ; 
  assign   tlMasterXbar__monitor__stopEn1  =  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_141  ; 
  assign   tlMasterXbar__monitor__stopEn2  =  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn3  =  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_148  ; 
  assign   tlMasterXbar__monitor__stopEn4  =  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn5  =  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_155  ; 
  assign   tlMasterXbar__monitor__stopEn6  =  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_160  ; 
  assign   tlMasterXbar__monitor__stopEn7  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_84  ; 
  assign   tlMasterXbar__monitor__stopEn8  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_141  ; 
  assign   tlMasterXbar__monitor__stopEn9  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn10  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_148  ; 
  assign   tlMasterXbar__monitor__stopEn11  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn12  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_155  ; 
  assign   tlMasterXbar__monitor__stopEn13  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_301  ; 
  assign   tlMasterXbar__monitor__stopEn14  =  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_160  ; 
  assign   tlMasterXbar__monitor__stopEn15  =  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_322  ; 
  assign   tlMasterXbar__monitor__stopEn16  =  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_377  ; 
  assign   tlMasterXbar__monitor__stopEn17  =  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn18  =  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn19  =  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_387  ; 
  assign   tlMasterXbar__monitor__stopEn20  =  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_391  ; 
  assign   tlMasterXbar__monitor__stopEn21  =  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_467  ; 
  assign   tlMasterXbar__monitor__stopEn22  =  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn23  =  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn24  =  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_387  ; 
  assign   tlMasterXbar__monitor__stopEn25  =  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_391  ; 
  assign   tlMasterXbar__monitor__stopEn26  =  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_467  ; 
  assign   tlMasterXbar__monitor__stopEn27  =  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn28  =  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn29  =  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_387  ; 
  assign   tlMasterXbar__monitor__stopEn30  =  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_569  ; 
  assign   tlMasterXbar__monitor__stopEn31  =  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_631  ; 
  assign   tlMasterXbar__monitor__stopEn32  =  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn33  =  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn34  =  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_641  ; 
  assign   tlMasterXbar__monitor__stopEn35  =  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_391  ; 
  assign   tlMasterXbar__monitor__stopEn36  =  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_631  ; 
  assign   tlMasterXbar__monitor__stopEn37  =  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn38  =  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn39  =  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_717  ; 
  assign   tlMasterXbar__monitor__stopEn40  =  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_391  ; 
  assign   tlMasterXbar__monitor__stopEn41  =  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_783  ; 
  assign   tlMasterXbar__monitor__stopEn42  =  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_144  ; 
  assign   tlMasterXbar__monitor__stopEn43  =  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_151  ; 
  assign   tlMasterXbar__monitor__stopEn44  =  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_793  ; 
  assign   tlMasterXbar__monitor__stopEn45  =  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_391  ; 
  assign   tlMasterXbar__monitor__stopEn46  =  tlMasterXbar__monitor__io_in_d_valid  &~  tlMasterXbar__monitor___T_805  ; 
  assign   tlMasterXbar__monitor__stopEn47  =  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_809  ; 
  assign   tlMasterXbar__monitor__stopEn48  =  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_813  ; 
  assign   tlMasterXbar__monitor__stopEn49  =  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_817  ; 
  assign   tlMasterXbar__monitor__stopEn50  =  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_821  ; 
  assign   tlMasterXbar__monitor__stopEn51  =  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_825  ; 
  assign   tlMasterXbar__monitor__stopEn52  =  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_809  ; 
  assign   tlMasterXbar__monitor__stopEn53  =  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_813  ; 
  assign   tlMasterXbar__monitor__stopEn54  =  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_840  ; 
  assign   tlMasterXbar__monitor__stopEn55  =  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_844  ; 
  assign   tlMasterXbar__monitor__stopEn56  =  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_821  ; 
  assign   tlMasterXbar__monitor__stopEn57  =  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_809  ; 
  assign   tlMasterXbar__monitor__stopEn58  =  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_813  ; 
  assign   tlMasterXbar__monitor__stopEn59  =  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_840  ; 
  assign   tlMasterXbar__monitor__stopEn60  =  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_844  ; 
  assign   tlMasterXbar__monitor__stopEn61  =  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_877  ; 
  assign   tlMasterXbar__monitor__stopEn62  =  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_809  ; 
  assign   tlMasterXbar__monitor__stopEn63  =  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_817  ; 
  assign   tlMasterXbar__monitor__stopEn64  =  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_821  ; 
  assign   tlMasterXbar__monitor__stopEn65  =  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_809  ; 
  assign   tlMasterXbar__monitor__stopEn66  =  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_817  ; 
  assign   tlMasterXbar__monitor__stopEn67  =  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_877  ; 
  assign   tlMasterXbar__monitor__stopEn68  =  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_809  ; 
  assign   tlMasterXbar__monitor__stopEn69  =  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_817  ; 
  assign   tlMasterXbar__monitor__stopEn70  =  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_821  ; 
  assign   tlMasterXbar__monitor__stopEn71  =  tlMasterXbar__monitor__io_in_b_valid  &~  tlMasterXbar__monitor___T_938  ; 
  assign   tlMasterXbar__monitor__stopEn72  =  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1016  ; 
  assign   tlMasterXbar__monitor__stopEn73  =  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1019  ; 
  assign   tlMasterXbar__monitor__stopEn74  =  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1022  ; 
  assign   tlMasterXbar__monitor__stopEn75  =  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1025  ; 
  assign   tlMasterXbar__monitor__stopEn76  =  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1029  ; 
  assign   tlMasterXbar__monitor__stopEn77  =  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1033  ; 
  assign   tlMasterXbar__monitor__stopEn78  =  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1037  ; 
  assign   tlMasterXbar__monitor__stopEn79  =  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__stopEn80  =  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1019  ; 
  assign   tlMasterXbar__monitor__stopEn81  =  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1022  ; 
  assign   tlMasterXbar__monitor__stopEn82  =  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1025  ; 
  assign   tlMasterXbar__monitor__stopEn83  =  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1102  ; 
  assign   tlMasterXbar__monitor__stopEn84  =  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1033  ; 
  assign   tlMasterXbar__monitor__stopEn85  =  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1037  ; 
  assign   tlMasterXbar__monitor__stopEn86  =  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__stopEn87  =  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1019  ; 
  assign   tlMasterXbar__monitor__stopEn88  =  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1022  ; 
  assign   tlMasterXbar__monitor__stopEn89  =  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1025  ; 
  assign   tlMasterXbar__monitor__stopEn90  =  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1102  ; 
  assign   tlMasterXbar__monitor__stopEn91  =  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1033  ; 
  assign   tlMasterXbar__monitor__stopEn92  =  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__stopEn93  =  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1019  ; 
  assign   tlMasterXbar__monitor__stopEn94  =  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1022  ; 
  assign   tlMasterXbar__monitor__stopEn95  =  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1025  ; 
  assign   tlMasterXbar__monitor__stopEn96  =  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1102  ; 
  assign   tlMasterXbar__monitor__stopEn97  =  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1250  ; 
  assign   tlMasterXbar__monitor__stopEn98  =  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__stopEn99  =  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1019  ; 
  assign   tlMasterXbar__monitor__stopEn100  =  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1022  ; 
  assign   tlMasterXbar__monitor__stopEn101  =  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1025  ; 
  assign   tlMasterXbar__monitor__stopEn102  =  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1033  ; 
  assign   tlMasterXbar__monitor__stopEn103  =  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__stopEn104  =  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1019  ; 
  assign   tlMasterXbar__monitor__stopEn105  =  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1022  ; 
  assign   tlMasterXbar__monitor__stopEn106  =  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1025  ; 
  assign   tlMasterXbar__monitor__stopEn107  =  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1033  ; 
  assign   tlMasterXbar__monitor__stopEn108  =  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor__reset  ; 
  assign   tlMasterXbar__monitor__stopEn109  =  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1019  ; 
  assign   tlMasterXbar__monitor__stopEn110  =  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1022  ; 
  assign   tlMasterXbar__monitor__stopEn111  =  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1025  ; 
  assign   tlMasterXbar__monitor__stopEn112  =  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1033  ; 
  assign   tlMasterXbar__monitor__stopEn113  =  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1037  ; 
  assign   tlMasterXbar__monitor__stopEn114  =  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1485  ; 
  assign   tlMasterXbar__monitor__stopEn115  =  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1488  ; 
  assign   tlMasterXbar__monitor__stopEn116  =  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1492  ; 
  assign   tlMasterXbar__monitor__stopEn117  =  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1495  ; 
  assign   tlMasterXbar__monitor__stopEn118  =  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1499  ; 
  assign   tlMasterXbar__monitor__stopEn119  =  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1485  ; 
  assign   tlMasterXbar__monitor__stopEn120  =  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1488  ; 
  assign   tlMasterXbar__monitor__stopEn121  =  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1492  ; 
  assign   tlMasterXbar__monitor__stopEn122  =  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1495  ; 
  assign   tlMasterXbar__monitor__stopEn123  =  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1499  ; 
  assign   tlMasterXbar__monitor__stopEn124  =  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1583  ; 
  assign   tlMasterXbar__monitor__stopEn125  =  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1640  ; 
  assign   tlMasterXbar__monitor__stopEn126  =  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1488  ; 
  assign   tlMasterXbar__monitor__stopEn127  =  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1492  ; 
  assign   tlMasterXbar__monitor__stopEn128  =  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1495  ; 
  assign   tlMasterXbar__monitor__stopEn129  =  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1499  ; 
  assign   tlMasterXbar__monitor__stopEn130  =  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1583  ; 
  assign   tlMasterXbar__monitor__stopEn131  =  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1640  ; 
  assign   tlMasterXbar__monitor__stopEn132  =  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1488  ; 
  assign   tlMasterXbar__monitor__stopEn133  =  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1492  ; 
  assign   tlMasterXbar__monitor__stopEn134  =  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1495  ; 
  assign   tlMasterXbar__monitor__stopEn135  =  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1499  ; 
  assign   tlMasterXbar__monitor__stopEn136  =  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1485  ; 
  assign   tlMasterXbar__monitor__stopEn137  =  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1488  ; 
  assign   tlMasterXbar__monitor__stopEn138  =  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1495  ; 
  assign   tlMasterXbar__monitor__stopEn139  =  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1805  ; 
  assign   tlMasterXbar__monitor__stopEn140  =  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1485  ; 
  assign   tlMasterXbar__monitor__stopEn141  =  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1488  ; 
  assign   tlMasterXbar__monitor__stopEn142  =  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1495  ; 
  assign   tlMasterXbar__monitor__stopEn143  =  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1805  ; 
  assign   tlMasterXbar__monitor__stopEn144  =  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1485  ; 
  assign   tlMasterXbar__monitor__stopEn145  =  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1488  ; 
  assign   tlMasterXbar__monitor__stopEn146  =  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1495  ; 
  assign   tlMasterXbar__monitor__stopEn147  =  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1805  ; 
  assign   tlMasterXbar__monitor__stopEn148  =  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1850  ; 
  assign   tlMasterXbar__monitor__stopEn149  =  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1854  ; 
  assign   tlMasterXbar__monitor__stopEn150  =  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1858  ; 
  assign   tlMasterXbar__monitor__stopEn151  =  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1862  ; 
  assign   tlMasterXbar__monitor__stopEn152  =  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1866  ; 
  assign   tlMasterXbar__monitor__stopEn153  =  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1874  ; 
  assign   tlMasterXbar__monitor__stopEn154  =  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1878  ; 
  assign   tlMasterXbar__monitor__stopEn155  =  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1882  ; 
  assign   tlMasterXbar__monitor__stopEn156  =  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1886  ; 
  assign   tlMasterXbar__monitor__stopEn157  =  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1890  ; 
  assign   tlMasterXbar__monitor__stopEn158  =  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1894  ; 
  assign   tlMasterXbar__monitor__stopEn159  =  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1902  ; 
  assign   tlMasterXbar__monitor__stopEn160  =  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1906  ; 
  assign   tlMasterXbar__monitor__stopEn161  =  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1910  ; 
  assign   tlMasterXbar__monitor__stopEn162  =  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1914  ; 
  assign   tlMasterXbar__monitor__stopEn163  =  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1918  ; 
  assign   tlMasterXbar__monitor__stopEn164  =  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1926  ; 
  assign   tlMasterXbar__monitor__stopEn165  =  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1930  ; 
  assign   tlMasterXbar__monitor__stopEn166  =  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1934  ; 
  assign   tlMasterXbar__monitor__stopEn167  =  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1938  ; 
  assign   tlMasterXbar__monitor__stopEn168  =  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1942  ; 
  assign   tlMasterXbar__monitor__stopEn169  =  tlMasterXbar__monitor___T_1949  &~  tlMasterXbar__monitor___T_1955  ; 
  assign   tlMasterXbar__monitor__stopEn170  =  tlMasterXbar__monitor___T_1960  &~  tlMasterXbar__monitor___T_1974  ; 
  assign   tlMasterXbar__monitor__stopEn171  =  tlMasterXbar__monitor___GEN_403  &~  tlMasterXbar__monitor___T_1980  ; 
  assign   tlMasterXbar__monitor__stopEn172  =  tlMasterXbar__monitor___GEN_403  &~  tlMasterXbar__monitor___T_1984  ; 
  assign   tlMasterXbar__monitor__stopEn173  =  tlMasterXbar__monitor___GEN_408  &~  tlMasterXbar__monitor___T_1992  ; 
  assign   tlMasterXbar__monitor__stopEn174  =  tlMasterXbar__monitor___GEN_408  &~  tlMasterXbar__monitor___T_1996  ; 
  assign   tlMasterXbar__monitor__stopEn175  =  tlMasterXbar__monitor___T_2004  &~  tlMasterXbar__monitor___T_2008  ; 
  assign   tlMasterXbar__monitor__stopEn176  =~  tlMasterXbar__monitor___T_2015  ; 
  assign   tlMasterXbar__monitor__stopEn177  =~  tlMasterXbar__monitor___T_2024  ; 
  assign   tlMasterXbar__monitor__stopEn178  =  tlMasterXbar__monitor___T_2039  &~  tlMasterXbar__monitor___T_2044  ; 
  assign   tlMasterXbar__monitor__stopEn179  =  tlMasterXbar__monitor___T_2048  &~  tlMasterXbar__monitor___T_2060  ; 
  assign   tlMasterXbar__monitor__stopEn180  =  tlMasterXbar__monitor___GEN_415  &~  tlMasterXbar__monitor___T_2064  ; 
  assign   tlMasterXbar__monitor__stopEn181  =  tlMasterXbar__monitor___GEN_418  &~  tlMasterXbar__monitor___T_2068  ; 
  assign   tlMasterXbar__monitor__stopEn182  =  tlMasterXbar__monitor___T_2075  &~  tlMasterXbar__monitor___T_2079  ; 
  assign   tlMasterXbar__monitor__stopEn183  =  tlMasterXbar__monitor___T_2081  &~  tlMasterXbar__monitor___T_2084  ; 
  assign   tlMasterXbar__monitor__stopEn184  =~  tlMasterXbar__monitor___T_2093  ; 
  assign   tlMasterXbar__monitor__stopEn185  =  tlMasterXbar__monitor___T_2104  &~  tlMasterXbar__monitor___T_2109  ; 
  assign   tlMasterXbar__monitor__stopEn186  =  tlMasterXbar__monitor___T_2111  &~  tlMasterXbar__monitor___T_2118  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or63  =  tlMasterXbar__monitor__stopEn0  |  tlMasterXbar__monitor__stopEn1  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or130  =  tlMasterXbar__monitor__stopEn3  |  tlMasterXbar__monitor__stopEn4  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or64  =  tlMasterXbar__monitor__stopEn2  |  tlMasterXbar__monitor__TLMonitor_23_or130  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or31  =  tlMasterXbar__monitor__TLMonitor_23_or63  |  tlMasterXbar__monitor__TLMonitor_23_or64  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or132  =  tlMasterXbar__monitor__stopEn6  |  tlMasterXbar__monitor__stopEn7  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or65  =  tlMasterXbar__monitor__stopEn5  |  tlMasterXbar__monitor__TLMonitor_23_or132  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or134  =  tlMasterXbar__monitor__stopEn9  |  tlMasterXbar__monitor__stopEn10  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or66  =  tlMasterXbar__monitor__stopEn8  |  tlMasterXbar__monitor__TLMonitor_23_or134  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or32  =  tlMasterXbar__monitor__TLMonitor_23_or65  |  tlMasterXbar__monitor__TLMonitor_23_or66  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or15  =  tlMasterXbar__monitor__TLMonitor_23_or31  |  tlMasterXbar__monitor__TLMonitor_23_or32  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or136  =  tlMasterXbar__monitor__stopEn12  |  tlMasterXbar__monitor__stopEn13  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or67  =  tlMasterXbar__monitor__stopEn11  |  tlMasterXbar__monitor__TLMonitor_23_or136  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or138  =  tlMasterXbar__monitor__stopEn15  |  tlMasterXbar__monitor__stopEn16  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or68  =  tlMasterXbar__monitor__stopEn14  |  tlMasterXbar__monitor__TLMonitor_23_or138  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or33  =  tlMasterXbar__monitor__TLMonitor_23_or67  |  tlMasterXbar__monitor__TLMonitor_23_or68  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or140  =  tlMasterXbar__monitor__stopEn18  |  tlMasterXbar__monitor__stopEn19  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or69  =  tlMasterXbar__monitor__stopEn17  |  tlMasterXbar__monitor__TLMonitor_23_or140  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or142  =  tlMasterXbar__monitor__stopEn21  |  tlMasterXbar__monitor__stopEn22  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or70  =  tlMasterXbar__monitor__stopEn20  |  tlMasterXbar__monitor__TLMonitor_23_or142  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or34  =  tlMasterXbar__monitor__TLMonitor_23_or69  |  tlMasterXbar__monitor__TLMonitor_23_or70  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or16  =  tlMasterXbar__monitor__TLMonitor_23_or33  |  tlMasterXbar__monitor__TLMonitor_23_or34  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or7  =  tlMasterXbar__monitor__TLMonitor_23_or15  |  tlMasterXbar__monitor__TLMonitor_23_or16  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or144  =  tlMasterXbar__monitor__stopEn24  |  tlMasterXbar__monitor__stopEn25  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or71  =  tlMasterXbar__monitor__stopEn23  |  tlMasterXbar__monitor__TLMonitor_23_or144  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or146  =  tlMasterXbar__monitor__stopEn27  |  tlMasterXbar__monitor__stopEn28  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or72  =  tlMasterXbar__monitor__stopEn26  |  tlMasterXbar__monitor__TLMonitor_23_or146  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or35  =  tlMasterXbar__monitor__TLMonitor_23_or71  |  tlMasterXbar__monitor__TLMonitor_23_or72  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or148  =  tlMasterXbar__monitor__stopEn30  |  tlMasterXbar__monitor__stopEn31  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or73  =  tlMasterXbar__monitor__stopEn29  |  tlMasterXbar__monitor__TLMonitor_23_or148  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or150  =  tlMasterXbar__monitor__stopEn33  |  tlMasterXbar__monitor__stopEn34  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or74  =  tlMasterXbar__monitor__stopEn32  |  tlMasterXbar__monitor__TLMonitor_23_or150  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or36  =  tlMasterXbar__monitor__TLMonitor_23_or73  |  tlMasterXbar__monitor__TLMonitor_23_or74  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or17  =  tlMasterXbar__monitor__TLMonitor_23_or35  |  tlMasterXbar__monitor__TLMonitor_23_or36  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or152  =  tlMasterXbar__monitor__stopEn36  |  tlMasterXbar__monitor__stopEn37  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or75  =  tlMasterXbar__monitor__stopEn35  |  tlMasterXbar__monitor__TLMonitor_23_or152  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or154  =  tlMasterXbar__monitor__stopEn39  |  tlMasterXbar__monitor__stopEn40  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or76  =  tlMasterXbar__monitor__stopEn38  |  tlMasterXbar__monitor__TLMonitor_23_or154  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or37  =  tlMasterXbar__monitor__TLMonitor_23_or75  |  tlMasterXbar__monitor__TLMonitor_23_or76  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or156  =  tlMasterXbar__monitor__stopEn42  |  tlMasterXbar__monitor__stopEn43  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or77  =  tlMasterXbar__monitor__stopEn41  |  tlMasterXbar__monitor__TLMonitor_23_or156  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or158  =  tlMasterXbar__monitor__stopEn45  |  tlMasterXbar__monitor__stopEn46  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or78  =  tlMasterXbar__monitor__stopEn44  |  tlMasterXbar__monitor__TLMonitor_23_or158  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or38  =  tlMasterXbar__monitor__TLMonitor_23_or77  |  tlMasterXbar__monitor__TLMonitor_23_or78  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or18  =  tlMasterXbar__monitor__TLMonitor_23_or37  |  tlMasterXbar__monitor__TLMonitor_23_or38  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or8  =  tlMasterXbar__monitor__TLMonitor_23_or17  |  tlMasterXbar__monitor__TLMonitor_23_or18  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or3  =  tlMasterXbar__monitor__TLMonitor_23_or7  |  tlMasterXbar__monitor__TLMonitor_23_or8  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or79  =  tlMasterXbar__monitor__stopEn47  |  tlMasterXbar__monitor__stopEn48  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or162  =  tlMasterXbar__monitor__stopEn50  |  tlMasterXbar__monitor__stopEn51  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or80  =  tlMasterXbar__monitor__stopEn49  |  tlMasterXbar__monitor__TLMonitor_23_or162  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or39  =  tlMasterXbar__monitor__TLMonitor_23_or79  |  tlMasterXbar__monitor__TLMonitor_23_or80  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or164  =  tlMasterXbar__monitor__stopEn53  |  tlMasterXbar__monitor__stopEn54  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or81  =  tlMasterXbar__monitor__stopEn52  |  tlMasterXbar__monitor__TLMonitor_23_or164  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or166  =  tlMasterXbar__monitor__stopEn56  |  tlMasterXbar__monitor__stopEn57  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or82  =  tlMasterXbar__monitor__stopEn55  |  tlMasterXbar__monitor__TLMonitor_23_or166  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or40  =  tlMasterXbar__monitor__TLMonitor_23_or81  |  tlMasterXbar__monitor__TLMonitor_23_or82  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or19  =  tlMasterXbar__monitor__TLMonitor_23_or39  |  tlMasterXbar__monitor__TLMonitor_23_or40  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or168  =  tlMasterXbar__monitor__stopEn59  |  tlMasterXbar__monitor__stopEn60  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or83  =  tlMasterXbar__monitor__stopEn58  |  tlMasterXbar__monitor__TLMonitor_23_or168  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or170  =  tlMasterXbar__monitor__stopEn62  |  tlMasterXbar__monitor__stopEn63  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or84  =  tlMasterXbar__monitor__stopEn61  |  tlMasterXbar__monitor__TLMonitor_23_or170  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or41  =  tlMasterXbar__monitor__TLMonitor_23_or83  |  tlMasterXbar__monitor__TLMonitor_23_or84  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or172  =  tlMasterXbar__monitor__stopEn65  |  tlMasterXbar__monitor__stopEn66  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or85  =  tlMasterXbar__monitor__stopEn64  |  tlMasterXbar__monitor__TLMonitor_23_or172  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or174  =  tlMasterXbar__monitor__stopEn68  |  tlMasterXbar__monitor__stopEn69  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or86  =  tlMasterXbar__monitor__stopEn67  |  tlMasterXbar__monitor__TLMonitor_23_or174  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or42  =  tlMasterXbar__monitor__TLMonitor_23_or85  |  tlMasterXbar__monitor__TLMonitor_23_or86  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or20  =  tlMasterXbar__monitor__TLMonitor_23_or41  |  tlMasterXbar__monitor__TLMonitor_23_or42  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or9  =  tlMasterXbar__monitor__TLMonitor_23_or19  |  tlMasterXbar__monitor__TLMonitor_23_or20  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or176  =  tlMasterXbar__monitor__stopEn71  |  tlMasterXbar__monitor__stopEn72  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or87  =  tlMasterXbar__monitor__stopEn70  |  tlMasterXbar__monitor__TLMonitor_23_or176  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or178  =  tlMasterXbar__monitor__stopEn74  |  tlMasterXbar__monitor__stopEn75  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or88  =  tlMasterXbar__monitor__stopEn73  |  tlMasterXbar__monitor__TLMonitor_23_or178  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or43  =  tlMasterXbar__monitor__TLMonitor_23_or87  |  tlMasterXbar__monitor__TLMonitor_23_or88  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or180  =  tlMasterXbar__monitor__stopEn77  |  tlMasterXbar__monitor__stopEn78  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or89  =  tlMasterXbar__monitor__stopEn76  |  tlMasterXbar__monitor__TLMonitor_23_or180  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or182  =  tlMasterXbar__monitor__stopEn80  |  tlMasterXbar__monitor__stopEn81  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or90  =  tlMasterXbar__monitor__stopEn79  |  tlMasterXbar__monitor__TLMonitor_23_or182  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or44  =  tlMasterXbar__monitor__TLMonitor_23_or89  |  tlMasterXbar__monitor__TLMonitor_23_or90  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or21  =  tlMasterXbar__monitor__TLMonitor_23_or43  |  tlMasterXbar__monitor__TLMonitor_23_or44  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or184  =  tlMasterXbar__monitor__stopEn83  |  tlMasterXbar__monitor__stopEn84  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or91  =  tlMasterXbar__monitor__stopEn82  |  tlMasterXbar__monitor__TLMonitor_23_or184  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or186  =  tlMasterXbar__monitor__stopEn86  |  tlMasterXbar__monitor__stopEn87  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or92  =  tlMasterXbar__monitor__stopEn85  |  tlMasterXbar__monitor__TLMonitor_23_or186  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or45  =  tlMasterXbar__monitor__TLMonitor_23_or91  |  tlMasterXbar__monitor__TLMonitor_23_or92  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or188  =  tlMasterXbar__monitor__stopEn89  |  tlMasterXbar__monitor__stopEn90  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or93  =  tlMasterXbar__monitor__stopEn88  |  tlMasterXbar__monitor__TLMonitor_23_or188  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or190  =  tlMasterXbar__monitor__stopEn92  |  tlMasterXbar__monitor__stopEn93  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or94  =  tlMasterXbar__monitor__stopEn91  |  tlMasterXbar__monitor__TLMonitor_23_or190  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or46  =  tlMasterXbar__monitor__TLMonitor_23_or93  |  tlMasterXbar__monitor__TLMonitor_23_or94  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or22  =  tlMasterXbar__monitor__TLMonitor_23_or45  |  tlMasterXbar__monitor__TLMonitor_23_or46  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or10  =  tlMasterXbar__monitor__TLMonitor_23_or21  |  tlMasterXbar__monitor__TLMonitor_23_or22  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or4  =  tlMasterXbar__monitor__TLMonitor_23_or9  |  tlMasterXbar__monitor__TLMonitor_23_or10  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or1  =  tlMasterXbar__monitor__TLMonitor_23_or3  |  tlMasterXbar__monitor__TLMonitor_23_or4  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or95  =  tlMasterXbar__monitor__stopEn94  |  tlMasterXbar__monitor__stopEn95  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or194  =  tlMasterXbar__monitor__stopEn97  |  tlMasterXbar__monitor__stopEn98  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or96  =  tlMasterXbar__monitor__stopEn96  |  tlMasterXbar__monitor__TLMonitor_23_or194  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or47  =  tlMasterXbar__monitor__TLMonitor_23_or95  |  tlMasterXbar__monitor__TLMonitor_23_or96  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or196  =  tlMasterXbar__monitor__stopEn100  |  tlMasterXbar__monitor__stopEn101  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or97  =  tlMasterXbar__monitor__stopEn99  |  tlMasterXbar__monitor__TLMonitor_23_or196  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or198  =  tlMasterXbar__monitor__stopEn103  |  tlMasterXbar__monitor__stopEn104  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or98  =  tlMasterXbar__monitor__stopEn102  |  tlMasterXbar__monitor__TLMonitor_23_or198  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or48  =  tlMasterXbar__monitor__TLMonitor_23_or97  |  tlMasterXbar__monitor__TLMonitor_23_or98  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or23  =  tlMasterXbar__monitor__TLMonitor_23_or47  |  tlMasterXbar__monitor__TLMonitor_23_or48  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or200  =  tlMasterXbar__monitor__stopEn106  |  tlMasterXbar__monitor__stopEn107  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or99  =  tlMasterXbar__monitor__stopEn105  |  tlMasterXbar__monitor__TLMonitor_23_or200  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or202  =  tlMasterXbar__monitor__stopEn109  |  tlMasterXbar__monitor__stopEn110  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or100  =  tlMasterXbar__monitor__stopEn108  |  tlMasterXbar__monitor__TLMonitor_23_or202  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or49  =  tlMasterXbar__monitor__TLMonitor_23_or99  |  tlMasterXbar__monitor__TLMonitor_23_or100  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or204  =  tlMasterXbar__monitor__stopEn112  |  tlMasterXbar__monitor__stopEn113  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or101  =  tlMasterXbar__monitor__stopEn111  |  tlMasterXbar__monitor__TLMonitor_23_or204  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or206  =  tlMasterXbar__monitor__stopEn115  |  tlMasterXbar__monitor__stopEn116  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or102  =  tlMasterXbar__monitor__stopEn114  |  tlMasterXbar__monitor__TLMonitor_23_or206  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or50  =  tlMasterXbar__monitor__TLMonitor_23_or101  |  tlMasterXbar__monitor__TLMonitor_23_or102  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or24  =  tlMasterXbar__monitor__TLMonitor_23_or49  |  tlMasterXbar__monitor__TLMonitor_23_or50  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or11  =  tlMasterXbar__monitor__TLMonitor_23_or23  |  tlMasterXbar__monitor__TLMonitor_23_or24  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or208  =  tlMasterXbar__monitor__stopEn118  |  tlMasterXbar__monitor__stopEn119  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or103  =  tlMasterXbar__monitor__stopEn117  |  tlMasterXbar__monitor__TLMonitor_23_or208  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or210  =  tlMasterXbar__monitor__stopEn121  |  tlMasterXbar__monitor__stopEn122  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or104  =  tlMasterXbar__monitor__stopEn120  |  tlMasterXbar__monitor__TLMonitor_23_or210  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or51  =  tlMasterXbar__monitor__TLMonitor_23_or103  |  tlMasterXbar__monitor__TLMonitor_23_or104  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or212  =  tlMasterXbar__monitor__stopEn124  |  tlMasterXbar__monitor__stopEn125  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or105  =  tlMasterXbar__monitor__stopEn123  |  tlMasterXbar__monitor__TLMonitor_23_or212  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or214  =  tlMasterXbar__monitor__stopEn127  |  tlMasterXbar__monitor__stopEn128  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or106  =  tlMasterXbar__monitor__stopEn126  |  tlMasterXbar__monitor__TLMonitor_23_or214  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or52  =  tlMasterXbar__monitor__TLMonitor_23_or105  |  tlMasterXbar__monitor__TLMonitor_23_or106  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or25  =  tlMasterXbar__monitor__TLMonitor_23_or51  |  tlMasterXbar__monitor__TLMonitor_23_or52  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or216  =  tlMasterXbar__monitor__stopEn130  |  tlMasterXbar__monitor__stopEn131  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or107  =  tlMasterXbar__monitor__stopEn129  |  tlMasterXbar__monitor__TLMonitor_23_or216  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or218  =  tlMasterXbar__monitor__stopEn133  |  tlMasterXbar__monitor__stopEn134  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or108  =  tlMasterXbar__monitor__stopEn132  |  tlMasterXbar__monitor__TLMonitor_23_or218  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or53  =  tlMasterXbar__monitor__TLMonitor_23_or107  |  tlMasterXbar__monitor__TLMonitor_23_or108  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or220  =  tlMasterXbar__monitor__stopEn136  |  tlMasterXbar__monitor__stopEn137  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or109  =  tlMasterXbar__monitor__stopEn135  |  tlMasterXbar__monitor__TLMonitor_23_or220  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or222  =  tlMasterXbar__monitor__stopEn139  |  tlMasterXbar__monitor__stopEn140  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or110  =  tlMasterXbar__monitor__stopEn138  |  tlMasterXbar__monitor__TLMonitor_23_or222  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or54  =  tlMasterXbar__monitor__TLMonitor_23_or109  |  tlMasterXbar__monitor__TLMonitor_23_or110  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or26  =  tlMasterXbar__monitor__TLMonitor_23_or53  |  tlMasterXbar__monitor__TLMonitor_23_or54  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or12  =  tlMasterXbar__monitor__TLMonitor_23_or25  |  tlMasterXbar__monitor__TLMonitor_23_or26  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or5  =  tlMasterXbar__monitor__TLMonitor_23_or11  |  tlMasterXbar__monitor__TLMonitor_23_or12  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or224  =  tlMasterXbar__monitor__stopEn142  |  tlMasterXbar__monitor__stopEn143  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or111  =  tlMasterXbar__monitor__stopEn141  |  tlMasterXbar__monitor__TLMonitor_23_or224  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or226  =  tlMasterXbar__monitor__stopEn145  |  tlMasterXbar__monitor__stopEn146  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or112  =  tlMasterXbar__monitor__stopEn144  |  tlMasterXbar__monitor__TLMonitor_23_or226  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or55  =  tlMasterXbar__monitor__TLMonitor_23_or111  |  tlMasterXbar__monitor__TLMonitor_23_or112  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or228  =  tlMasterXbar__monitor__stopEn148  |  tlMasterXbar__monitor__stopEn149  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or113  =  tlMasterXbar__monitor__stopEn147  |  tlMasterXbar__monitor__TLMonitor_23_or228  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or230  =  tlMasterXbar__monitor__stopEn151  |  tlMasterXbar__monitor__stopEn152  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or114  =  tlMasterXbar__monitor__stopEn150  |  tlMasterXbar__monitor__TLMonitor_23_or230  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or56  =  tlMasterXbar__monitor__TLMonitor_23_or113  |  tlMasterXbar__monitor__TLMonitor_23_or114  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or27  =  tlMasterXbar__monitor__TLMonitor_23_or55  |  tlMasterXbar__monitor__TLMonitor_23_or56  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or232  =  tlMasterXbar__monitor__stopEn154  |  tlMasterXbar__monitor__stopEn155  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or115  =  tlMasterXbar__monitor__stopEn153  |  tlMasterXbar__monitor__TLMonitor_23_or232  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or234  =  tlMasterXbar__monitor__stopEn157  |  tlMasterXbar__monitor__stopEn158  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or116  =  tlMasterXbar__monitor__stopEn156  |  tlMasterXbar__monitor__TLMonitor_23_or234  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or57  =  tlMasterXbar__monitor__TLMonitor_23_or115  |  tlMasterXbar__monitor__TLMonitor_23_or116  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or236  =  tlMasterXbar__monitor__stopEn160  |  tlMasterXbar__monitor__stopEn161  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or117  =  tlMasterXbar__monitor__stopEn159  |  tlMasterXbar__monitor__TLMonitor_23_or236  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or238  =  tlMasterXbar__monitor__stopEn163  |  tlMasterXbar__monitor__stopEn164  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or118  =  tlMasterXbar__monitor__stopEn162  |  tlMasterXbar__monitor__TLMonitor_23_or238  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or58  =  tlMasterXbar__monitor__TLMonitor_23_or117  |  tlMasterXbar__monitor__TLMonitor_23_or118  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or28  =  tlMasterXbar__monitor__TLMonitor_23_or57  |  tlMasterXbar__monitor__TLMonitor_23_or58  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or13  =  tlMasterXbar__monitor__TLMonitor_23_or27  |  tlMasterXbar__monitor__TLMonitor_23_or28  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or240  =  tlMasterXbar__monitor__stopEn166  |  tlMasterXbar__monitor__stopEn167  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or119  =  tlMasterXbar__monitor__stopEn165  |  tlMasterXbar__monitor__TLMonitor_23_or240  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or242  =  tlMasterXbar__monitor__stopEn169  |  tlMasterXbar__monitor__stopEn170  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or120  =  tlMasterXbar__monitor__stopEn168  |  tlMasterXbar__monitor__TLMonitor_23_or242  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or59  =  tlMasterXbar__monitor__TLMonitor_23_or119  |  tlMasterXbar__monitor__TLMonitor_23_or120  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or244  =  tlMasterXbar__monitor__stopEn172  |  tlMasterXbar__monitor__stopEn173  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or121  =  tlMasterXbar__monitor__stopEn171  |  tlMasterXbar__monitor__TLMonitor_23_or244  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or246  =  tlMasterXbar__monitor__stopEn175  |  tlMasterXbar__monitor__stopEn176  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or122  =  tlMasterXbar__monitor__stopEn174  |  tlMasterXbar__monitor__TLMonitor_23_or246  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or60  =  tlMasterXbar__monitor__TLMonitor_23_or121  |  tlMasterXbar__monitor__TLMonitor_23_or122  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or29  =  tlMasterXbar__monitor__TLMonitor_23_or59  |  tlMasterXbar__monitor__TLMonitor_23_or60  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or248  =  tlMasterXbar__monitor__stopEn178  |  tlMasterXbar__monitor__stopEn179  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or123  =  tlMasterXbar__monitor__stopEn177  |  tlMasterXbar__monitor__TLMonitor_23_or248  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or250  =  tlMasterXbar__monitor__stopEn181  |  tlMasterXbar__monitor__stopEn182  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or124  =  tlMasterXbar__monitor__stopEn180  |  tlMasterXbar__monitor__TLMonitor_23_or250  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or61  =  tlMasterXbar__monitor__TLMonitor_23_or123  |  tlMasterXbar__monitor__TLMonitor_23_or124  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or252  =  tlMasterXbar__monitor__stopEn184  |  tlMasterXbar__monitor__stopEn185  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or125  =  tlMasterXbar__monitor__stopEn183  |  tlMasterXbar__monitor__TLMonitor_23_or252  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or254  =  tlMasterXbar__monitor__plusarg_reader_metaAssert_wire  |  tlMasterXbar__monitor__plusarg_reader_1_metaAssert_wire  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or126  =  tlMasterXbar__monitor__stopEn186  |  tlMasterXbar__monitor__TLMonitor_23_or254  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or62  =  tlMasterXbar__monitor__TLMonitor_23_or125  |  tlMasterXbar__monitor__TLMonitor_23_or126  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or30  =  tlMasterXbar__monitor__TLMonitor_23_or61  |  tlMasterXbar__monitor__TLMonitor_23_or62  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or14  =  tlMasterXbar__monitor__TLMonitor_23_or29  |  tlMasterXbar__monitor__TLMonitor_23_or30  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or6  =  tlMasterXbar__monitor__TLMonitor_23_or13  |  tlMasterXbar__monitor__TLMonitor_23_or14  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or2  =  tlMasterXbar__monitor__TLMonitor_23_or5  |  tlMasterXbar__monitor__TLMonitor_23_or6  ; 
  assign   tlMasterXbar__monitor__TLMonitor_23_or0  =  tlMasterXbar__monitor__TLMonitor_23_or1  |  tlMasterXbar__monitor__TLMonitor_23_or2  ; 
  assign   tlMasterXbar__monitor__metaAssert  =  tlMasterXbar__monitor__TLMonitor_23_metaAssert  ; initial
    begin 
    end  
  always @( posedge   tlMasterXbar__monitor__clock  )
       begin 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__a_first_counter   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__a_first_counter   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___a_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__a_first  )
                       begin 
                         if (  tlMasterXbar__monitor__a_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__a_first_counter   <=  tlMasterXbar__monitor__a_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__a_first_counter   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__a_first_counter   <=  tlMasterXbar__monitor__a_first_counter1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__opcode   <=3'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1869  )
               begin  
                  tlMasterXbar__monitor__opcode   <=  tlMasterXbar__monitor__io_in_a_bits_opcode  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__param   <=3'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1869  )
               begin  
                  tlMasterXbar__monitor__param   <=  tlMasterXbar__monitor__io_in_a_bits_param  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__size   <=4'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1869  )
               begin  
                  tlMasterXbar__monitor__size   <=  tlMasterXbar__monitor__io_in_a_bits_size  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__source   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1869  )
               begin  
                  tlMasterXbar__monitor__source   <=  tlMasterXbar__monitor__io_in_a_bits_source  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__address   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1869  )
               begin  
                  tlMasterXbar__monitor__address   <=  tlMasterXbar__monitor__io_in_a_bits_address  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__d_first_counter   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__d_first_counter   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___d_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__d_first  )
                       begin 
                         if (  tlMasterXbar__monitor__d_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__d_first_counter   <=  tlMasterXbar__monitor__d_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__d_first_counter   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__d_first_counter   <=  tlMasterXbar__monitor__d_first_counter1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__opcode_1   <=3'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1897  )
               begin  
                  tlMasterXbar__monitor__opcode_1   <=  tlMasterXbar__monitor__io_in_d_bits_opcode  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__param_1   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1897  )
               begin  
                  tlMasterXbar__monitor__param_1   <=  tlMasterXbar__monitor__io_in_d_bits_param  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__size_1   <=4'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1897  )
               begin  
                  tlMasterXbar__monitor__size_1   <=  tlMasterXbar__monitor__io_in_d_bits_size  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__source_1   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1897  )
               begin  
                  tlMasterXbar__monitor__source_1   <=  tlMasterXbar__monitor__io_in_d_bits_source  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__sink   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1897  )
               begin  
                  tlMasterXbar__monitor__sink   <=  tlMasterXbar__monitor__io_in_d_bits_sink  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__denied   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1897  )
               begin  
                  tlMasterXbar__monitor__denied   <=  tlMasterXbar__monitor__io_in_d_bits_denied  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__b_first_counter   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__b_first_counter   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor__b_first_done  )
                  begin 
                    if (  tlMasterXbar__monitor__b_first  )
                       begin  
                          tlMasterXbar__monitor__b_first_counter   <=9'h0;
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__b_first_counter   <=  tlMasterXbar__monitor__b_first_counter1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__opcode_2   <=3'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1921  )
               begin  
                  tlMasterXbar__monitor__opcode_2   <=  tlMasterXbar__monitor__io_in_b_bits_opcode  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__param_2   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1921  )
               begin  
                  tlMasterXbar__monitor__param_2   <=  tlMasterXbar__monitor__io_in_b_bits_param  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__size_2   <=4'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1921  )
               begin  
                  tlMasterXbar__monitor__size_2   <=  tlMasterXbar__monitor__io_in_b_bits_size  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__source_2   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1921  )
               begin  
                  tlMasterXbar__monitor__source_2   <=  tlMasterXbar__monitor__io_in_b_bits_source  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__address_1   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1921  )
               begin  
                  tlMasterXbar__monitor__address_1   <=  tlMasterXbar__monitor__io_in_b_bits_address  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__c_first_counter   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__c_first_counter   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___c_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__c_first  )
                       begin 
                         if (  tlMasterXbar__monitor__c_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__c_first_counter   <=  tlMasterXbar__monitor__c_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__c_first_counter   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__c_first_counter   <=  tlMasterXbar__monitor__c_first_counter1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__opcode_3   <=3'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1945  )
               begin  
                  tlMasterXbar__monitor__opcode_3   <=  tlMasterXbar__monitor__io_in_c_bits_opcode  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__param_3   <=3'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1945  )
               begin  
                  tlMasterXbar__monitor__param_3   <=  tlMasterXbar__monitor__io_in_c_bits_param  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__size_3   <=4'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1945  )
               begin  
                  tlMasterXbar__monitor__size_3   <=  tlMasterXbar__monitor__io_in_c_bits_size  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__source_3   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1945  )
               begin  
                  tlMasterXbar__monitor__source_3   <=  tlMasterXbar__monitor__io_in_c_bits_source  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__address_2   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor___T_1945  )
               begin  
                  tlMasterXbar__monitor__address_2   <=  tlMasterXbar__monitor__io_in_c_bits_address  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__inflight   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__inflight   <=2'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor__inflight   <=  tlMasterXbar__monitor___inflight_T_2  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__inflight_opcodes   <=8'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__inflight_opcodes   <=8'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor__inflight_opcodes   <=  tlMasterXbar__monitor___inflight_opcodes_T_2  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__inflight_sizes   <=16'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__inflight_sizes   <=16'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor__inflight_sizes   <=  tlMasterXbar__monitor___inflight_sizes_T_2  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__a_first_counter_1   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__a_first_counter_1   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___a_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__a_first_1  )
                       begin 
                         if (  tlMasterXbar__monitor__a_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__a_first_counter_1   <=  tlMasterXbar__monitor__a_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__a_first_counter_1   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__a_first_counter_1   <=  tlMasterXbar__monitor__a_first_counter1_1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__d_first_counter_1   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__d_first_counter_1   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___d_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__d_first_1  )
                       begin 
                         if (  tlMasterXbar__monitor__d_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__d_first_counter_1   <=  tlMasterXbar__monitor__d_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__d_first_counter_1   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__d_first_counter_1   <=  tlMasterXbar__monitor__d_first_counter1_1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__watchdog   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__watchdog   <=32'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___T_2028  )
                  begin  
                     tlMasterXbar__monitor__watchdog   <=32'h0;
                  end 
                else 
                  begin  
                     tlMasterXbar__monitor__watchdog   <=  tlMasterXbar__monitor___watchdog_T_1  ;
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__inflight_1   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__inflight_1   <=2'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor__inflight_1   <=  tlMasterXbar__monitor___inflight_T_5  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__inflight_sizes_1   <=16'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__inflight_sizes_1   <=16'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor__inflight_sizes_1   <=  tlMasterXbar__monitor___inflight_sizes_T_5  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__c_first_counter_1   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__c_first_counter_1   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___c_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__c_first_1  )
                       begin 
                         if (  tlMasterXbar__monitor__c_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__c_first_counter_1   <=  tlMasterXbar__monitor__c_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__c_first_counter_1   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__c_first_counter_1   <=  tlMasterXbar__monitor__c_first_counter1_1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__d_first_counter_2   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__d_first_counter_2   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___d_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__d_first_2  )
                       begin 
                         if (  tlMasterXbar__monitor__d_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__d_first_counter_2   <=  tlMasterXbar__monitor__d_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__d_first_counter_2   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__d_first_counter_2   <=  tlMasterXbar__monitor__d_first_counter1_2  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__watchdog_1   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__watchdog_1   <=32'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___T_2097  )
                  begin  
                     tlMasterXbar__monitor__watchdog_1   <=32'h0;
                  end 
                else 
                  begin  
                     tlMasterXbar__monitor__watchdog_1   <=  tlMasterXbar__monitor___watchdog_T_3  ;
                  end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__inflight_2   <=4'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__inflight_2   <=4'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor__inflight_2   <=  tlMasterXbar__monitor___inflight_T_8  ;
               end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__d_first_counter_3   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor__reset  )
               begin  
                  tlMasterXbar__monitor__d_first_counter_3   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor___d_first_T  )
                  begin 
                    if (  tlMasterXbar__monitor__d_first_3  )
                       begin 
                         if (  tlMasterXbar__monitor__d_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor__d_first_counter_3   <=  tlMasterXbar__monitor__d_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor__d_first_counter_3   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor__d_first_counter_3   <=  tlMasterXbar__monitor__d_first_counter1_3  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_84  )
            begin $display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_84  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_141  )
            begin $display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_141  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_148  )
            begin $display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_148  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_155  )
            begin $display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_155  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_160  )
            begin $display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_111  &~  tlMasterXbar__monitor___T_160  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_84  )
            begin $display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_84  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_141  )
            begin $display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_141  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_148  )
            begin $display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_148  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_155  )
            begin $display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_155  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_301  )
            begin $display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_301  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_160  )
            begin $display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_125  &~  tlMasterXbar__monitor___T_160  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_322  )
            begin $display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_322  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_377  )
            begin $display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_377  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel Get carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel Get address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_387  )
            begin $display("Assertion failed: 'A' channel Get carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_387  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_391  )
            begin $display("Assertion failed: 'A' channel Get contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_141  &~  tlMasterXbar__monitor___T_391  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_467  )
            begin $display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_467  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_387  )
            begin $display("Assertion failed: 'A' channel PutFull carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_387  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_391  )
            begin $display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_153  &~  tlMasterXbar__monitor___T_391  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_467  )
            begin $display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_467  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_387  )
            begin $display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_387  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_569  )
            begin $display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_163  &~  tlMasterXbar__monitor___T_569  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_631  )
            begin $display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_631  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_641  )
            begin $display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_641  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_391  )
            begin $display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_173  &~  tlMasterXbar__monitor___T_391  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_631  )
            begin $display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_631  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel Logical address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_717  )
            begin $display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_717  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_391  )
            begin $display("Assertion failed: 'A' channel Logical contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_183  &~  tlMasterXbar__monitor___T_391  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_783  )
            begin $display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_783  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_144  )
            begin $display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_144  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_151  )
            begin $display("Assertion failed: 'A' channel Hint address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_151  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_793  )
            begin $display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_793  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_391  )
            begin $display("Assertion failed: 'A' channel Hint contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_193  &~  tlMasterXbar__monitor___T_391  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor__io_in_d_valid  &~  tlMasterXbar__monitor___T_805  )
            begin $display("Assertion failed: 'D' channel has invalid opcode (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor__io_in_d_valid  &~  tlMasterXbar__monitor___T_805  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_809  )
            begin $display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_809  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_813  )
            begin $display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_813  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_817  )
            begin $display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_817  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_821  )
            begin $display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_821  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_825  )
            begin $display("Assertion failed: 'D' channel ReleaseAck is denied (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_203  &~  tlMasterXbar__monitor___T_825  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_809  )
            begin $display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_809  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_813  )
            begin $display("Assertion failed: 'D' channel Grant smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_813  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_840  )
            begin $display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_840  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_844  )
            begin $display("Assertion failed: 'D' channel Grant carries toN param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_844  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_821  )
            begin $display("Assertion failed: 'D' channel Grant is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_213  &~  tlMasterXbar__monitor___T_821  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_809  )
            begin $display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_809  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_813  )
            begin $display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_813  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_840  )
            begin $display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_840  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_844  )
            begin $display("Assertion failed: 'D' channel GrantData carries toN param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_844  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_877  )
            begin $display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_223  &~  tlMasterXbar__monitor___T_877  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_809  )
            begin $display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_809  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_817  )
            begin $display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_817  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_821  )
            begin $display("Assertion failed: 'D' channel AccessAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_233  &~  tlMasterXbar__monitor___T_821  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_809  )
            begin $display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_809  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_817  )
            begin $display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_817  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_877  )
            begin $display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_239  &~  tlMasterXbar__monitor___T_877  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_809  )
            begin $display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_809  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_817  )
            begin $display("Assertion failed: 'D' channel HintAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_817  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_821  )
            begin $display("Assertion failed: 'D' channel HintAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_245  &~  tlMasterXbar__monitor___T_821  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor__io_in_b_valid  &~  tlMasterXbar__monitor___T_938  )
            begin $display("Assertion failed: 'B' channel has invalid opcode (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor__io_in_b_valid  &~  tlMasterXbar__monitor___T_938  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1016  )
            begin $display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1016  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("Assertion failed: 'B' channel Probe carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("Assertion failed: 'B' channel Probe address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1029  )
            begin $display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1029  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("Assertion failed: 'B' channel Probe contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1037  )
            begin $display("Assertion failed: 'B' channel Probe is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_251  &~  tlMasterXbar__monitor___T_1037  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor__reset  )
            begin $display("Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor__reset  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("Assertion failed: 'B' channel Get carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("Assertion failed: 'B' channel Get carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("Assertion failed: 'B' channel Get address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1102  )
            begin $display("Assertion failed: 'B' channel Get carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1102  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("Assertion failed: 'B' channel Get contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1037  )
            begin $display("Assertion failed: 'B' channel Get is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_265  &~  tlMasterXbar__monitor___T_1037  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor__reset  )
            begin $display("Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor__reset  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("Assertion failed: 'B' channel PutFull carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("Assertion failed: 'B' channel PutFull carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("Assertion failed: 'B' channel PutFull address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1102  )
            begin $display("Assertion failed: 'B' channel PutFull carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1102  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("Assertion failed: 'B' channel PutFull contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_279  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor__reset  )
            begin $display("Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor__reset  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("Assertion failed: 'B' channel PutPartial address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1102  )
            begin $display("Assertion failed: 'B' channel PutPartial carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1102  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1250  )
            begin $display("Assertion failed: 'B' channel PutPartial contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_291  &~  tlMasterXbar__monitor___T_1250  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor__reset  )
            begin $display("Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor__reset  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_303  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor__reset  )
            begin $display("Assertion failed: 'B' channel carries Logical type unsupported by client (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor__reset  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("Assertion failed: 'B' channel Logical carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("Assertion failed: 'B' channel Logical carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("Assertion failed: 'B' channel Logical address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("Assertion failed: 'B' channel Logical contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_313  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor__reset  )
            begin $display("Assertion failed: 'B' channel carries Hint type unsupported by client (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor__reset  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("Assertion failed: 'B' channel Hint carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1019  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("Assertion failed: 'B' channel Hint carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1022  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("Assertion failed: 'B' channel Hint address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1025  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("Assertion failed: 'B' channel Hint contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1033  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1037  )
            begin $display("Assertion failed: 'B' channel Hint is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_323  &~  tlMasterXbar__monitor___T_1037  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_335  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_345  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1583  )
            begin $display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1583  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1640  )
            begin $display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1640  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("Assertion failed: 'C' channel Release carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("Assertion failed: 'C' channel Release smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("Assertion failed: 'C' channel Release address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("Assertion failed: 'C' channel Release carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_355  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1583  )
            begin $display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1583  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1640  )
            begin $display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1640  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1492  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_367  &~  tlMasterXbar__monitor___T_1499  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1805  )
            begin $display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_379  &~  tlMasterXbar__monitor___T_1805  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1805  )
            begin $display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_387  &~  tlMasterXbar__monitor___T_1805  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1485  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("Assertion failed: 'C' channel HintAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1488  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1495  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1805  )
            begin $display("Assertion failed: 'C' channel HintAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_395  &~  tlMasterXbar__monitor___T_1805  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1850  )
            begin $display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1850  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1854  )
            begin $display("Assertion failed: 'A' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1854  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1858  )
            begin $display("Assertion failed: 'A' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1858  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1862  )
            begin $display("Assertion failed: 'A' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1862  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1866  )
            begin $display("Assertion failed: 'A' channel address changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1847  &~  tlMasterXbar__monitor___T_1866  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1874  )
            begin $display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1874  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1878  )
            begin $display("Assertion failed: 'D' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1878  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1882  )
            begin $display("Assertion failed: 'D' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1882  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1886  )
            begin $display("Assertion failed: 'D' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1886  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1890  )
            begin $display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1890  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1894  )
            begin $display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1871  &~  tlMasterXbar__monitor___T_1894  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1902  )
            begin $display("Assertion failed: 'B' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1902  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1906  )
            begin $display("Assertion failed: 'B' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1906  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1910  )
            begin $display("Assertion failed: 'B' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1910  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1914  )
            begin $display("Assertion failed: 'B' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1914  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1918  )
            begin $display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1899  &~  tlMasterXbar__monitor___T_1918  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1926  )
            begin $display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1926  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1930  )
            begin $display("Assertion failed: 'C' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1930  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1934  )
            begin $display("Assertion failed: 'C' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1934  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1938  )
            begin $display("Assertion failed: 'C' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1938  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1942  )
            begin $display("Assertion failed: 'C' channel address changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1923  &~  tlMasterXbar__monitor___T_1942  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1949  &~  tlMasterXbar__monitor___T_1955  )
            begin $display("Assertion failed: 'A' channel re-used a source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1949  &~  tlMasterXbar__monitor___T_1955  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_1960  &~  tlMasterXbar__monitor___T_1974  )
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_1960  &~  tlMasterXbar__monitor___T_1974  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_403  &~  tlMasterXbar__monitor___T_1980  )
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_403  &~  tlMasterXbar__monitor___T_1980  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_403  &~  tlMasterXbar__monitor___T_1984  )
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_403  &~  tlMasterXbar__monitor___T_1984  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_408  &~  tlMasterXbar__monitor___T_1992  )
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_408  &~  tlMasterXbar__monitor___T_1992  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_408  &~  tlMasterXbar__monitor___T_1996  )
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_408  &~  tlMasterXbar__monitor___T_1996  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_2004  &~  tlMasterXbar__monitor___T_2008  )
            begin $display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_2004  &~  tlMasterXbar__monitor___T_2008  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar__monitor___T_2015  )
            begin $display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (~  tlMasterXbar__monitor___T_2015  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar__monitor___T_2024  )
            begin $display("Assertion failed: TileLink timeout expired (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~  tlMasterXbar__monitor___T_2024  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_2039  &~  tlMasterXbar__monitor___T_2044  )
            begin $display("Assertion failed: 'C' channel re-used a source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_2039  &~  tlMasterXbar__monitor___T_2044  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_2048  &~  tlMasterXbar__monitor___T_2060  )
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_2048  &~  tlMasterXbar__monitor___T_2060  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_415  &~  tlMasterXbar__monitor___T_2064  )
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_415  &~  tlMasterXbar__monitor___T_2064  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___GEN_418  &~  tlMasterXbar__monitor___T_2068  )
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___GEN_418  &~  tlMasterXbar__monitor___T_2068  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_2075  &~  tlMasterXbar__monitor___T_2079  )
            begin $display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_2075  &~  tlMasterXbar__monitor___T_2079  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_2081  &~  tlMasterXbar__monitor___T_2084  )
            begin $display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_2081  &~  tlMasterXbar__monitor___T_2084  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar__monitor___T_2093  )
            begin $display("Assertion failed: TileLink timeout expired (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~  tlMasterXbar__monitor___T_2093  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_2104  &~  tlMasterXbar__monitor___T_2109  )
            begin $display("Assertion failed: 'D' channel re-used a sink ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_2104  &~  tlMasterXbar__monitor___T_2109  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor___T_2111  &~  tlMasterXbar__monitor___T_2118  )
            begin $display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor___T_2111  &~  tlMasterXbar__monitor___T_2118  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor__metaReset  )
            begin  
               tlMasterXbar__monitor__TLMonitor_23_metaAssert   <=1'h0;
            end 
          else 
            begin  
               tlMasterXbar__monitor__TLMonitor_23_metaAssert   <=  tlMasterXbar__monitor__TLMonitor_23_metaAssert  |  tlMasterXbar__monitor__TLMonitor_23_or0  ;
            end 
       end
 
assign tlMasterXbar__monitor__clock = tlMasterXbar__monitor_clock;
assign tlMasterXbar__monitor__reset = tlMasterXbar__monitor_reset;
assign tlMasterXbar__monitor__io_in_a_ready = tlMasterXbar__monitor_io_in_a_ready;
assign tlMasterXbar__monitor__io_in_a_valid = tlMasterXbar__monitor_io_in_a_valid;
assign tlMasterXbar__monitor__io_in_a_bits_opcode = tlMasterXbar__monitor_io_in_a_bits_opcode;
assign tlMasterXbar__monitor__io_in_a_bits_param = tlMasterXbar__monitor_io_in_a_bits_param;
assign tlMasterXbar__monitor__io_in_a_bits_size = tlMasterXbar__monitor_io_in_a_bits_size;
assign tlMasterXbar__monitor__io_in_a_bits_source = tlMasterXbar__monitor_io_in_a_bits_source;
assign tlMasterXbar__monitor__io_in_a_bits_address = tlMasterXbar__monitor_io_in_a_bits_address;
assign tlMasterXbar__monitor__io_in_a_bits_mask = tlMasterXbar__monitor_io_in_a_bits_mask;
assign tlMasterXbar__monitor__io_in_b_ready = tlMasterXbar__monitor_io_in_b_ready;
assign tlMasterXbar__monitor__io_in_b_valid = tlMasterXbar__monitor_io_in_b_valid;
assign tlMasterXbar__monitor__io_in_b_bits_opcode = tlMasterXbar__monitor_io_in_b_bits_opcode;
assign tlMasterXbar__monitor__io_in_b_bits_param = tlMasterXbar__monitor_io_in_b_bits_param;
assign tlMasterXbar__monitor__io_in_b_bits_size = tlMasterXbar__monitor_io_in_b_bits_size;
assign tlMasterXbar__monitor__io_in_b_bits_source = tlMasterXbar__monitor_io_in_b_bits_source;
assign tlMasterXbar__monitor__io_in_b_bits_address = tlMasterXbar__monitor_io_in_b_bits_address;
assign tlMasterXbar__monitor__io_in_b_bits_mask = tlMasterXbar__monitor_io_in_b_bits_mask;
assign tlMasterXbar__monitor__io_in_b_bits_corrupt = tlMasterXbar__monitor_io_in_b_bits_corrupt;
assign tlMasterXbar__monitor__io_in_c_ready = tlMasterXbar__monitor_io_in_c_ready;
assign tlMasterXbar__monitor__io_in_c_valid = tlMasterXbar__monitor_io_in_c_valid;
assign tlMasterXbar__monitor__io_in_c_bits_opcode = tlMasterXbar__monitor_io_in_c_bits_opcode;
assign tlMasterXbar__monitor__io_in_c_bits_param = tlMasterXbar__monitor_io_in_c_bits_param;
assign tlMasterXbar__monitor__io_in_c_bits_size = tlMasterXbar__monitor_io_in_c_bits_size;
assign tlMasterXbar__monitor__io_in_c_bits_source = tlMasterXbar__monitor_io_in_c_bits_source;
assign tlMasterXbar__monitor__io_in_c_bits_address = tlMasterXbar__monitor_io_in_c_bits_address;
assign tlMasterXbar__monitor__io_in_d_ready = tlMasterXbar__monitor_io_in_d_ready;
assign tlMasterXbar__monitor__io_in_d_valid = tlMasterXbar__monitor_io_in_d_valid;
assign tlMasterXbar__monitor__io_in_d_bits_opcode = tlMasterXbar__monitor_io_in_d_bits_opcode;
assign tlMasterXbar__monitor__io_in_d_bits_param = tlMasterXbar__monitor_io_in_d_bits_param;
assign tlMasterXbar__monitor__io_in_d_bits_size = tlMasterXbar__monitor_io_in_d_bits_size;
assign tlMasterXbar__monitor__io_in_d_bits_source = tlMasterXbar__monitor_io_in_d_bits_source;
assign tlMasterXbar__monitor__io_in_d_bits_sink = tlMasterXbar__monitor_io_in_d_bits_sink;
assign tlMasterXbar__monitor__io_in_d_bits_denied = tlMasterXbar__monitor_io_in_d_bits_denied;
assign tlMasterXbar__monitor__io_in_d_bits_corrupt = tlMasterXbar__monitor_io_in_d_bits_corrupt;
assign tlMasterXbar__monitor__io_in_e_ready = tlMasterXbar__monitor_io_in_e_ready;
assign tlMasterXbar__monitor__io_in_e_valid = tlMasterXbar__monitor_io_in_e_valid;
assign tlMasterXbar__monitor__io_in_e_bits_sink = tlMasterXbar__monitor_io_in_e_bits_sink;
assign tlMasterXbar__monitor_io_covSum = tlMasterXbar__monitor__io_covSum;
assign tlMasterXbar__monitor_metaAssert = tlMasterXbar__monitor__metaAssert;
assign tlMasterXbar__monitor__metaReset = tlMasterXbar__monitor_metaReset;
  
  
wire  tlMasterXbar__monitor_1__clock;
wire  tlMasterXbar__monitor_1__reset;
wire  tlMasterXbar__monitor_1__io_in_a_ready;
wire  tlMasterXbar__monitor_1__io_in_a_valid;
wire [31:0] tlMasterXbar__monitor_1__io_in_a_bits_address;
wire  tlMasterXbar__monitor_1__io_in_d_valid;
wire [2:0] tlMasterXbar__monitor_1__io_in_d_bits_opcode;
wire [1:0] tlMasterXbar__monitor_1__io_in_d_bits_param;
wire [3:0] tlMasterXbar__monitor_1__io_in_d_bits_size;
wire [1:0] tlMasterXbar__monitor_1__io_in_d_bits_sink;
wire  tlMasterXbar__monitor_1__io_in_d_bits_denied;
wire  tlMasterXbar__monitor_1__io_in_d_bits_corrupt;
wire [29:0] tlMasterXbar__monitor_1__io_covSum;
wire  tlMasterXbar__monitor_1__metaAssert;
wire  tlMasterXbar__monitor_1__metaReset;
 
   wire[31:0]  tlMasterXbar__monitor_1__plusarg_reader_out  ; 
   wire[31:0]  tlMasterXbar__monitor_1__plusarg_reader_1_out  ; 
   wire[31:0]  tlMasterXbar__monitor_1___is_aligned_T  ; 
   wire  tlMasterXbar__monitor_1__is_aligned  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_7  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_26  ; 
   wire  tlMasterXbar__monitor_1___T_27  ; 
   wire[31:0]  tlMasterXbar__monitor_1___T_28  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_29  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_31  ; 
   wire  tlMasterXbar__monitor_1___T_32  ; 
   wire[31:0]  tlMasterXbar__monitor_1___T_33  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_34  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_36  ; 
   wire  tlMasterXbar__monitor_1___T_37  ; 
   wire[31:0]  tlMasterXbar__monitor_1___T_38  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_39  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_41  ; 
   wire  tlMasterXbar__monitor_1___T_42  ; 
   wire[31:0]  tlMasterXbar__monitor_1___T_43  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_44  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_46  ; 
   wire  tlMasterXbar__monitor_1___T_47  ; 
   wire[31:0]  tlMasterXbar__monitor_1___T_48  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_49  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_51  ; 
   wire  tlMasterXbar__monitor_1___T_52  ; 
   wire[31:0]  tlMasterXbar__monitor_1___T_63  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_64  ; 
   wire[32:0]  tlMasterXbar__monitor_1___T_66  ; 
   wire  tlMasterXbar__monitor_1___T_67  ; 
   wire  tlMasterXbar__monitor_1___T_134  ; 
   wire  tlMasterXbar__monitor_1___T_341  ; 
   wire  tlMasterXbar__monitor_1___T_342  ; 
   wire  tlMasterXbar__monitor_1___T_343  ; 
   wire  tlMasterXbar__monitor_1___T_344  ; 
   wire  tlMasterXbar__monitor_1___T_345  ; 
   wire  tlMasterXbar__monitor_1___T_348  ; 
   wire  tlMasterXbar__monitor_1___T_350  ; 
   wire  tlMasterXbar__monitor_1___T_766  ; 
   wire  tlMasterXbar__monitor_1___T_768  ; 
   wire  tlMasterXbar__monitor_1___T_770  ; 
   wire  tlMasterXbar__monitor_1___T_774  ; 
   wire  tlMasterXbar__monitor_1___T_776  ; 
   wire  tlMasterXbar__monitor_1___T_778  ; 
   wire  tlMasterXbar__monitor_1___T_780  ; 
   wire  tlMasterXbar__monitor_1___T_784  ; 
   wire  tlMasterXbar__monitor_1___T_788  ; 
   wire  tlMasterXbar__monitor_1___T_790  ; 
   wire  tlMasterXbar__monitor_1___T_801  ; 
   wire  tlMasterXbar__monitor_1___T_803  ; 
   wire  tlMasterXbar__monitor_1___T_805  ; 
   wire  tlMasterXbar__monitor_1___T_807  ; 
   wire  tlMasterXbar__monitor_1___T_818  ; 
   wire  tlMasterXbar__monitor_1___T_838  ; 
   wire  tlMasterXbar__monitor_1___T_840  ; 
   wire  tlMasterXbar__monitor_1___T_847  ; 
   wire  tlMasterXbar__monitor_1___T_864  ; 
   wire  tlMasterXbar__monitor_1___T_882  ; 
   wire  tlMasterXbar__monitor_1__a_first_done  ; 
   reg[8:0]  tlMasterXbar__monitor_1__a_first_counter  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_0  ; 
   wire[8:0]  tlMasterXbar__monitor_1__a_first_counter1  ; 
   wire  tlMasterXbar__monitor_1__a_first  ; 
   reg[31:0]  tlMasterXbar__monitor_1__address  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_1  ; 
   wire  tlMasterXbar__monitor_1___T_912  ; 
   wire  tlMasterXbar__monitor_1___T_929  ; 
   wire  tlMasterXbar__monitor_1___T_931  ; 
   wire  tlMasterXbar__monitor_1___T_934  ; 
   wire[26:0]  tlMasterXbar__monitor_1___d_first_beats1_decode_T_1  ; 
   wire[8:0]  tlMasterXbar__monitor_1__d_first_beats1_decode  ; 
   wire  tlMasterXbar__monitor_1__d_first_beats1_opdata  ; 
   reg[8:0]  tlMasterXbar__monitor_1__d_first_counter  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_2  ; 
   wire[8:0]  tlMasterXbar__monitor_1__d_first_counter1  ; 
   wire  tlMasterXbar__monitor_1__d_first  ; 
   reg[2:0]  tlMasterXbar__monitor_1__opcode_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_3  ; 
   reg[1:0]  tlMasterXbar__monitor_1__param_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_4  ; 
   reg[3:0]  tlMasterXbar__monitor_1__size_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_5  ; 
   reg[1:0]  tlMasterXbar__monitor_1__sink  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_6  ; 
   reg  tlMasterXbar__monitor_1__denied  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_7  ; 
   wire  tlMasterXbar__monitor_1___T_936  ; 
   wire  tlMasterXbar__monitor_1___T_937  ; 
   wire  tlMasterXbar__monitor_1___T_939  ; 
   wire  tlMasterXbar__monitor_1___T_941  ; 
   wire  tlMasterXbar__monitor_1___T_943  ; 
   wire  tlMasterXbar__monitor_1___T_945  ; 
   wire  tlMasterXbar__monitor_1___T_947  ; 
   wire  tlMasterXbar__monitor_1___T_953  ; 
   wire  tlMasterXbar__monitor_1___T_955  ; 
   wire  tlMasterXbar__monitor_1___T_957  ; 
   wire  tlMasterXbar__monitor_1___T_959  ; 
   wire  tlMasterXbar__monitor_1___T_962  ; 
   reg  tlMasterXbar__monitor_1__inflight  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_8  ; 
   reg[3:0]  tlMasterXbar__monitor_1__inflight_opcodes  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_9  ; 
   reg[7:0]  tlMasterXbar__monitor_1__inflight_sizes  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_10  ; 
   reg[8:0]  tlMasterXbar__monitor_1__a_first_counter_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_11  ; 
   wire[8:0]  tlMasterXbar__monitor_1__a_first_counter1_1  ; 
   wire  tlMasterXbar__monitor_1__a_first_1  ; 
   reg[8:0]  tlMasterXbar__monitor_1__d_first_counter_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_12  ; 
   wire[8:0]  tlMasterXbar__monitor_1__d_first_counter1_1  ; 
   wire  tlMasterXbar__monitor_1__d_first_1  ; 
   wire[15:0]  tlMasterXbar__monitor_1___a_opcode_lookup_T_5  ; 
   wire[15:0]  tlMasterXbar__monitor_1___GEN_71  ; 
   wire[15:0]  tlMasterXbar__monitor_1___a_opcode_lookup_T_6  ; 
   wire[15:0]  tlMasterXbar__monitor_1___a_opcode_lookup_T_7  ; 
   wire[15:0]  tlMasterXbar__monitor_1___a_size_lookup_T_5  ; 
   wire[15:0]  tlMasterXbar__monitor_1___GEN_73  ; 
   wire[15:0]  tlMasterXbar__monitor_1___a_size_lookup_T_6  ; 
   wire[15:0]  tlMasterXbar__monitor_1___a_size_lookup_T_7  ; 
   wire  tlMasterXbar__monitor_1___T_963  ; 
   wire[1:0]  tlMasterXbar__monitor_1___GEN_15  ; 
   wire  tlMasterXbar__monitor_1___T_966  ; 
   wire[3:0]  tlMasterXbar__monitor_1__a_opcodes_set_interm  ; 
   wire[18:0]  tlMasterXbar__monitor_1___a_opcodes_set_T_1  ; 
   wire[4:0]  tlMasterXbar__monitor_1__a_sizes_set_interm  ; 
   wire[19:0]  tlMasterXbar__monitor_1___a_sizes_set_T_1  ; 
   wire  tlMasterXbar__monitor_1___T_972  ; 
   wire[1:0]  tlMasterXbar__monitor_1___GEN_16  ; 
   wire[18:0]  tlMasterXbar__monitor_1___GEN_19  ; 
   wire[19:0]  tlMasterXbar__monitor_1___GEN_20  ; 
   wire  tlMasterXbar__monitor_1___T_974  ; 
   wire  tlMasterXbar__monitor_1___T_977  ; 
   wire[1:0]  tlMasterXbar__monitor_1___GEN_21  ; 
   wire[30:0]  tlMasterXbar__monitor_1___d_opcodes_clr_T_5  ; 
   wire[30:0]  tlMasterXbar__monitor_1___d_sizes_clr_T_5  ; 
   wire[30:0]  tlMasterXbar__monitor_1___GEN_23  ; 
   wire[30:0]  tlMasterXbar__monitor_1___GEN_24  ; 
   wire  tlMasterXbar__monitor_1___T_989  ; 
   wire  tlMasterXbar__monitor_1___T_991  ; 
   wire  tlMasterXbar__monitor_1___T_995  ; 
   wire  tlMasterXbar__monitor_1___T_997  ; 
   wire  tlMasterXbar__monitor_1___T_999  ; 
   wire  tlMasterXbar__monitor_1___T_1001  ; 
   wire[3:0]  tlMasterXbar__monitor_1__a_opcode_lookup  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_43  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_44  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_45  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_46  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_47  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_48  ; 
   wire  tlMasterXbar__monitor_1___T_1004  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_55  ; 
   wire[2:0]  tlMasterXbar__monitor_1___GEN_56  ; 
   wire  tlMasterXbar__monitor_1___T_1006  ; 
   wire  tlMasterXbar__monitor_1___T_1007  ; 
   wire  tlMasterXbar__monitor_1___T_1009  ; 
   wire[7:0]  tlMasterXbar__monitor_1__a_size_lookup  ; 
   wire[7:0]  tlMasterXbar__monitor_1___GEN_75  ; 
   wire  tlMasterXbar__monitor_1___T_1011  ; 
   wire  tlMasterXbar__monitor_1___T_1013  ; 
   wire  tlMasterXbar__monitor_1___T_1016  ; 
   wire  tlMasterXbar__monitor_1___T_1017  ; 
   wire  tlMasterXbar__monitor_1___T_1021  ; 
   wire  tlMasterXbar__monitor_1___T_1025  ; 
   wire  tlMasterXbar__monitor_1__a_set_wo_ready  ; 
   wire  tlMasterXbar__monitor_1__d_clr_wo_ready  ; 
   wire  tlMasterXbar__monitor_1___T_1027  ; 
   wire  tlMasterXbar__monitor_1___T_1028  ; 
   wire  tlMasterXbar__monitor_1___T_1030  ; 
   wire  tlMasterXbar__monitor_1___T_1032  ; 
   wire  tlMasterXbar__monitor_1__a_set  ; 
   wire  tlMasterXbar__monitor_1___inflight_T  ; 
   wire  tlMasterXbar__monitor_1___inflight_T_2  ; 
   wire[3:0]  tlMasterXbar__monitor_1__a_opcodes_set  ; 
   wire[3:0]  tlMasterXbar__monitor_1___inflight_opcodes_T  ; 
   wire[3:0]  tlMasterXbar__monitor_1__d_opcodes_clr  ; 
   wire[3:0]  tlMasterXbar__monitor_1___inflight_opcodes_T_2  ; 
   wire[7:0]  tlMasterXbar__monitor_1__a_sizes_set  ; 
   wire[7:0]  tlMasterXbar__monitor_1___inflight_sizes_T  ; 
   wire[7:0]  tlMasterXbar__monitor_1__d_sizes_clr  ; 
   wire[7:0]  tlMasterXbar__monitor_1___inflight_sizes_T_2  ; 
   reg[31:0]  tlMasterXbar__monitor_1__watchdog  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_13  ; 
   wire  tlMasterXbar__monitor_1___T_1034  ; 
   wire  tlMasterXbar__monitor_1___T_1036  ; 
   wire  tlMasterXbar__monitor_1___T_1037  ; 
   wire  tlMasterXbar__monitor_1___T_1038  ; 
   wire  tlMasterXbar__monitor_1___T_1039  ; 
   wire  tlMasterXbar__monitor_1___T_1041  ; 
   wire[31:0]  tlMasterXbar__monitor_1___watchdog_T_1  ; 
   wire  tlMasterXbar__monitor_1___T_1045  ; 
   reg  tlMasterXbar__monitor_1__inflight_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_14  ; 
   reg[7:0]  tlMasterXbar__monitor_1__inflight_sizes_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_15  ; 
   reg[8:0]  tlMasterXbar__monitor_1__d_first_counter_2  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_16  ; 
   wire[8:0]  tlMasterXbar__monitor_1__d_first_counter1_2  ; 
   wire  tlMasterXbar__monitor_1__d_first_2  ; 
   wire[15:0]  tlMasterXbar__monitor_1___GEN_78  ; 
   wire[15:0]  tlMasterXbar__monitor_1___c_size_lookup_T_6  ; 
   wire[15:0]  tlMasterXbar__monitor_1___c_size_lookup_T_7  ; 
   wire  tlMasterXbar__monitor_1___T_1063  ; 
   wire  tlMasterXbar__monitor_1___T_1065  ; 
   wire[1:0]  tlMasterXbar__monitor_1___GEN_66  ; 
   wire[30:0]  tlMasterXbar__monitor_1___GEN_69  ; 
   wire  tlMasterXbar__monitor_1___T_1077  ; 
   wire[7:0]  tlMasterXbar__monitor_1__c_size_lookup  ; 
   wire  tlMasterXbar__monitor_1___T_1083  ; 
   wire  tlMasterXbar__monitor_1___T_1085  ; 
   wire  tlMasterXbar__monitor_1___T_1098  ; 
   wire  tlMasterXbar__monitor_1__d_clr_wo_ready_1  ; 
   wire  tlMasterXbar__monitor_1___T_1101  ; 
   wire  tlMasterXbar__monitor_1___inflight_T_5  ; 
   wire[7:0]  tlMasterXbar__monitor_1__d_sizes_clr_1  ; 
   wire[7:0]  tlMasterXbar__monitor_1___inflight_sizes_T_5  ; 
   reg[31:0]  tlMasterXbar__monitor_1__watchdog_1  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_17  ; 
   wire  tlMasterXbar__monitor_1___T_1103  ; 
   wire  tlMasterXbar__monitor_1___T_1105  ; 
   wire  tlMasterXbar__monitor_1___T_1106  ; 
   wire  tlMasterXbar__monitor_1___T_1107  ; 
   wire  tlMasterXbar__monitor_1___T_1108  ; 
   wire  tlMasterXbar__monitor_1___T_1110  ; 
   wire[31:0]  tlMasterXbar__monitor_1___watchdog_T_3  ; 
   wire  tlMasterXbar__monitor_1___GEN_81  ; 
   wire  tlMasterXbar__monitor_1___GEN_89  ; 
   wire  tlMasterXbar__monitor_1___GEN_97  ; 
   wire  tlMasterXbar__monitor_1___GEN_105  ; 
   wire  tlMasterXbar__monitor_1___GEN_109  ; 
   wire  tlMasterXbar__monitor_1___GEN_113  ; 
   wire  tlMasterXbar__monitor_1___GEN_117  ; 
   wire  tlMasterXbar__monitor_1___GEN_122  ; 
   wire[29:0]  tlMasterXbar__monitor_1__TLMonitor_24_covSum  ; 
   wire  tlMasterXbar__monitor_1__stopEn0  ; 
   wire  tlMasterXbar__monitor_1__stopEn1  ; 
   wire  tlMasterXbar__monitor_1__stopEn2  ; 
   wire  tlMasterXbar__monitor_1__stopEn3  ; 
   wire  tlMasterXbar__monitor_1__stopEn4  ; 
   wire  tlMasterXbar__monitor_1__stopEn5  ; 
   wire  tlMasterXbar__monitor_1__stopEn6  ; 
   wire  tlMasterXbar__monitor_1__stopEn7  ; 
   wire  tlMasterXbar__monitor_1__stopEn8  ; 
   wire  tlMasterXbar__monitor_1__stopEn9  ; 
   wire  tlMasterXbar__monitor_1__stopEn10  ; 
   wire  tlMasterXbar__monitor_1__stopEn11  ; 
   wire  tlMasterXbar__monitor_1__stopEn12  ; 
   wire  tlMasterXbar__monitor_1__stopEn13  ; 
   wire  tlMasterXbar__monitor_1__stopEn14  ; 
   wire  tlMasterXbar__monitor_1__stopEn15  ; 
   wire  tlMasterXbar__monitor_1__stopEn16  ; 
   wire  tlMasterXbar__monitor_1__stopEn17  ; 
   wire  tlMasterXbar__monitor_1__stopEn18  ; 
   wire  tlMasterXbar__monitor_1__stopEn19  ; 
   wire  tlMasterXbar__monitor_1__stopEn20  ; 
   wire  tlMasterXbar__monitor_1__stopEn21  ; 
   wire  tlMasterXbar__monitor_1__stopEn22  ; 
   wire  tlMasterXbar__monitor_1__stopEn23  ; 
   wire  tlMasterXbar__monitor_1__stopEn24  ; 
   wire  tlMasterXbar__monitor_1__stopEn25  ; 
   wire  tlMasterXbar__monitor_1__stopEn26  ; 
   wire  tlMasterXbar__monitor_1__stopEn27  ; 
   wire  tlMasterXbar__monitor_1__stopEn28  ; 
   wire  tlMasterXbar__monitor_1__stopEn29  ; 
   wire  tlMasterXbar__monitor_1__stopEn30  ; 
   wire  tlMasterXbar__monitor_1__stopEn31  ; 
   wire  tlMasterXbar__monitor_1__stopEn32  ; 
   wire  tlMasterXbar__monitor_1__stopEn33  ; 
   wire  tlMasterXbar__monitor_1__stopEn34  ; 
   wire  tlMasterXbar__monitor_1__stopEn35  ; 
   wire  tlMasterXbar__monitor_1__stopEn36  ; 
   wire  tlMasterXbar__monitor_1__stopEn37  ; 
   wire  tlMasterXbar__monitor_1__stopEn38  ; 
   wire  tlMasterXbar__monitor_1__stopEn39  ; 
   wire  tlMasterXbar__monitor_1__plusarg_reader_metaAssert_wire  ; 
   wire  tlMasterXbar__monitor_1__plusarg_reader_1_metaAssert_wire  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or15  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or34  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or16  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or7  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or17  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or38  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or18  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or8  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or3  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or19  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or42  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or20  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or9  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or44  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or21  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or46  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or22  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or10  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or4  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or1  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or23  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or50  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or24  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or11  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or25  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or54  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or26  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or12  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or5  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or27  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or58  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or28  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or13  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or60  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or29  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or62  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or30  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or14  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or6  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or2  ; 
   wire  tlMasterXbar__monitor_1__TLMonitor_24_or0  ; 
   reg  tlMasterXbar__monitor_1__TLMonitor_24_metaAssert  ; 
   reg[31:0]  tlMasterXbar__monitor_1___RAND_18  ; 
  assign   tlMasterXbar__monitor_1___is_aligned_T  =  tlMasterXbar__monitor_1__io_in_a_bits_address  &32'h3f; 
  assign   tlMasterXbar__monitor_1__is_aligned  =  tlMasterXbar__monitor_1___is_aligned_T  ==32'h0; 
  assign   tlMasterXbar__monitor_1___T_7  ={1'b0,$signed(  tlMasterXbar__monitor_1__io_in_a_bits_address  )}; 
  assign   tlMasterXbar__monitor_1___T_26  =$signed(  tlMasterXbar__monitor_1___T_7  )&-33'sh1000; 
  assign   tlMasterXbar__monitor_1___T_27  =$signed(  tlMasterXbar__monitor_1___T_26  )==33'sh0; 
  assign   tlMasterXbar__monitor_1___T_28  =  tlMasterXbar__monitor_1__io_in_a_bits_address  ^32'h3000; 
  assign   tlMasterXbar__monitor_1___T_29  ={1'b0,$signed(  tlMasterXbar__monitor_1___T_28  )}; 
  assign   tlMasterXbar__monitor_1___T_31  =$signed(  tlMasterXbar__monitor_1___T_29  )&-33'sh1000; 
  assign   tlMasterXbar__monitor_1___T_32  =$signed(  tlMasterXbar__monitor_1___T_31  )==33'sh0; 
  assign   tlMasterXbar__monitor_1___T_33  =  tlMasterXbar__monitor_1__io_in_a_bits_address  ^32'h10000; 
  assign   tlMasterXbar__monitor_1___T_34  ={1'b0,$signed(  tlMasterXbar__monitor_1___T_33  )}; 
  assign   tlMasterXbar__monitor_1___T_36  =$signed(  tlMasterXbar__monitor_1___T_34  )&-33'sh10000; 
  assign   tlMasterXbar__monitor_1___T_37  =$signed(  tlMasterXbar__monitor_1___T_36  )==33'sh0; 
  assign   tlMasterXbar__monitor_1___T_38  =  tlMasterXbar__monitor_1__io_in_a_bits_address  ^32'h2000000; 
  assign   tlMasterXbar__monitor_1___T_39  ={1'b0,$signed(  tlMasterXbar__monitor_1___T_38  )}; 
  assign   tlMasterXbar__monitor_1___T_41  =$signed(  tlMasterXbar__monitor_1___T_39  )&-33'sh10000; 
  assign   tlMasterXbar__monitor_1___T_42  =$signed(  tlMasterXbar__monitor_1___T_41  )==33'sh0; 
  assign   tlMasterXbar__monitor_1___T_43  =  tlMasterXbar__monitor_1__io_in_a_bits_address  ^32'hc000000; 
  assign   tlMasterXbar__monitor_1___T_44  ={1'b0,$signed(  tlMasterXbar__monitor_1___T_43  )}; 
  assign   tlMasterXbar__monitor_1___T_46  =$signed(  tlMasterXbar__monitor_1___T_44  )&-33'sh4000000; 
  assign   tlMasterXbar__monitor_1___T_47  =$signed(  tlMasterXbar__monitor_1___T_46  )==33'sh0; 
  assign   tlMasterXbar__monitor_1___T_48  =  tlMasterXbar__monitor_1__io_in_a_bits_address  ^32'h60000000; 
  assign   tlMasterXbar__monitor_1___T_49  ={1'b0,$signed(  tlMasterXbar__monitor_1___T_48  )}; 
  assign   tlMasterXbar__monitor_1___T_51  =$signed(  tlMasterXbar__monitor_1___T_49  )&-33'sh20000000; 
  assign   tlMasterXbar__monitor_1___T_52  =$signed(  tlMasterXbar__monitor_1___T_51  )==33'sh0; 
  assign   tlMasterXbar__monitor_1___T_63  =  tlMasterXbar__monitor_1__io_in_a_bits_address  ^32'h80000000; 
  assign   tlMasterXbar__monitor_1___T_64  ={1'b0,$signed(  tlMasterXbar__monitor_1___T_63  )}; 
  assign   tlMasterXbar__monitor_1___T_66  =$signed(  tlMasterXbar__monitor_1___T_64  )&-33'sh10000000; 
  assign   tlMasterXbar__monitor_1___T_67  =$signed(  tlMasterXbar__monitor_1___T_66  )==33'sh0; 
  assign   tlMasterXbar__monitor_1___T_134  =  tlMasterXbar__monitor_1__is_aligned  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_341  =  tlMasterXbar__monitor_1___T_27  |  tlMasterXbar__monitor_1___T_37  ; 
  assign   tlMasterXbar__monitor_1___T_342  =  tlMasterXbar__monitor_1___T_341  |  tlMasterXbar__monitor_1___T_42  ; 
  assign   tlMasterXbar__monitor_1___T_343  =  tlMasterXbar__monitor_1___T_342  |  tlMasterXbar__monitor_1___T_47  ; 
  assign   tlMasterXbar__monitor_1___T_344  =  tlMasterXbar__monitor_1___T_343  |  tlMasterXbar__monitor_1___T_52  ; 
  assign   tlMasterXbar__monitor_1___T_345  =  tlMasterXbar__monitor_1___T_344  |  tlMasterXbar__monitor_1___T_67  ; 
  assign   tlMasterXbar__monitor_1___T_348  =  tlMasterXbar__monitor_1___T_32  |  tlMasterXbar__monitor_1___T_345  ; 
  assign   tlMasterXbar__monitor_1___T_350  =  tlMasterXbar__monitor_1___T_348  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_766  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  <=3'h6; 
  assign   tlMasterXbar__monitor_1___T_768  =  tlMasterXbar__monitor_1___T_766  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_770  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h6; 
  assign   tlMasterXbar__monitor_1___T_774  =  tlMasterXbar__monitor_1__io_in_d_bits_size  >=4'h3; 
  assign   tlMasterXbar__monitor_1___T_776  =  tlMasterXbar__monitor_1___T_774  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_778  =  tlMasterXbar__monitor_1__io_in_d_bits_param  ==2'h0; 
  assign   tlMasterXbar__monitor_1___T_780  =  tlMasterXbar__monitor_1___T_778  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_784  =~  tlMasterXbar__monitor_1__io_in_d_bits_corrupt  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_788  =~  tlMasterXbar__monitor_1__io_in_d_bits_denied  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_790  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h4; 
  assign   tlMasterXbar__monitor_1___T_801  =  tlMasterXbar__monitor_1__io_in_d_bits_param  <=2'h2; 
  assign   tlMasterXbar__monitor_1___T_803  =  tlMasterXbar__monitor_1___T_801  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_805  =  tlMasterXbar__monitor_1__io_in_d_bits_param  !=2'h2; 
  assign   tlMasterXbar__monitor_1___T_807  =  tlMasterXbar__monitor_1___T_805  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_818  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h5; 
  assign   tlMasterXbar__monitor_1___T_838  =~  tlMasterXbar__monitor_1__io_in_d_bits_denied  |  tlMasterXbar__monitor_1__io_in_d_bits_corrupt  ; 
  assign   tlMasterXbar__monitor_1___T_840  =  tlMasterXbar__monitor_1___T_838  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_847  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h0; 
  assign   tlMasterXbar__monitor_1___T_864  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h1; 
  assign   tlMasterXbar__monitor_1___T_882  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h2; 
  assign   tlMasterXbar__monitor_1__a_first_done  =  tlMasterXbar__monitor_1__io_in_a_ready  &  tlMasterXbar__monitor_1__io_in_a_valid  ; 
  assign   tlMasterXbar__monitor_1__a_first_counter1  =  tlMasterXbar__monitor_1__a_first_counter  -9'h1; 
  assign   tlMasterXbar__monitor_1__a_first  =  tlMasterXbar__monitor_1__a_first_counter  ==9'h0; 
  assign   tlMasterXbar__monitor_1___T_912  =  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1__a_first  ; 
  assign   tlMasterXbar__monitor_1___T_929  =  tlMasterXbar__monitor_1__io_in_a_bits_address  ==  tlMasterXbar__monitor_1__address  ; 
  assign   tlMasterXbar__monitor_1___T_931  =  tlMasterXbar__monitor_1___T_929  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_934  =  tlMasterXbar__monitor_1__a_first_done  &  tlMasterXbar__monitor_1__a_first  ; 
  assign   tlMasterXbar__monitor_1___d_first_beats1_decode_T_1  =27'hfff<<  tlMasterXbar__monitor_1__io_in_d_bits_size  ; 
  assign   tlMasterXbar__monitor_1__d_first_beats1_decode  =~  tlMasterXbar__monitor_1___d_first_beats1_decode_T_1  [11:3]; 
  assign   tlMasterXbar__monitor_1__d_first_beats1_opdata  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  [0]; 
  assign   tlMasterXbar__monitor_1__d_first_counter1  =  tlMasterXbar__monitor_1__d_first_counter  -9'h1; 
  assign   tlMasterXbar__monitor_1__d_first  =  tlMasterXbar__monitor_1__d_first_counter  ==9'h0; 
  assign   tlMasterXbar__monitor_1___T_936  =  tlMasterXbar__monitor_1__io_in_d_valid  &~  tlMasterXbar__monitor_1__d_first  ; 
  assign   tlMasterXbar__monitor_1___T_937  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==  tlMasterXbar__monitor_1__opcode_1  ; 
  assign   tlMasterXbar__monitor_1___T_939  =  tlMasterXbar__monitor_1___T_937  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_941  =  tlMasterXbar__monitor_1__io_in_d_bits_param  ==  tlMasterXbar__monitor_1__param_1  ; 
  assign   tlMasterXbar__monitor_1___T_943  =  tlMasterXbar__monitor_1___T_941  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_945  =  tlMasterXbar__monitor_1__io_in_d_bits_size  ==  tlMasterXbar__monitor_1__size_1  ; 
  assign   tlMasterXbar__monitor_1___T_947  =  tlMasterXbar__monitor_1___T_945  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_953  =  tlMasterXbar__monitor_1__io_in_d_bits_sink  ==  tlMasterXbar__monitor_1__sink  ; 
  assign   tlMasterXbar__monitor_1___T_955  =  tlMasterXbar__monitor_1___T_953  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_957  =  tlMasterXbar__monitor_1__io_in_d_bits_denied  ==  tlMasterXbar__monitor_1__denied  ; 
  assign   tlMasterXbar__monitor_1___T_959  =  tlMasterXbar__monitor_1___T_957  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_962  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__d_first  ; 
  assign   tlMasterXbar__monitor_1__a_first_counter1_1  =  tlMasterXbar__monitor_1__a_first_counter_1  -9'h1; 
  assign   tlMasterXbar__monitor_1__a_first_1  =  tlMasterXbar__monitor_1__a_first_counter_1  ==9'h0; 
  assign   tlMasterXbar__monitor_1__d_first_counter1_1  =  tlMasterXbar__monitor_1__d_first_counter_1  -9'h1; 
  assign   tlMasterXbar__monitor_1__d_first_1  =  tlMasterXbar__monitor_1__d_first_counter_1  ==9'h0; 
  assign   tlMasterXbar__monitor_1___a_opcode_lookup_T_5  =16'h10-16'h1; 
  assign   tlMasterXbar__monitor_1___GEN_71  ={12'b0,  tlMasterXbar__monitor_1__inflight_opcodes  }; 
  assign   tlMasterXbar__monitor_1___a_opcode_lookup_T_6  =  tlMasterXbar__monitor_1___GEN_71  &  tlMasterXbar__monitor_1___a_opcode_lookup_T_5  ; 
  assign   tlMasterXbar__monitor_1___a_opcode_lookup_T_7  ={1'b0,  tlMasterXbar__monitor_1___a_opcode_lookup_T_6  [15:1]}; 
  assign   tlMasterXbar__monitor_1___a_size_lookup_T_5  =16'h100-16'h1; 
  assign   tlMasterXbar__monitor_1___GEN_73  ={8'b0,  tlMasterXbar__monitor_1__inflight_sizes  }; 
  assign   tlMasterXbar__monitor_1___a_size_lookup_T_6  =  tlMasterXbar__monitor_1___GEN_73  &  tlMasterXbar__monitor_1___a_size_lookup_T_5  ; 
  assign   tlMasterXbar__monitor_1___a_size_lookup_T_7  ={1'b0,  tlMasterXbar__monitor_1___a_size_lookup_T_6  [15:1]}; 
  assign   tlMasterXbar__monitor_1___T_963  =  tlMasterXbar__monitor_1__io_in_a_valid  &  tlMasterXbar__monitor_1__a_first_1  ; 
  assign   tlMasterXbar__monitor_1___GEN_15  =  tlMasterXbar__monitor_1___T_963   ? 2'h1:2'h0; 
  assign   tlMasterXbar__monitor_1___T_966  =  tlMasterXbar__monitor_1__a_first_done  &  tlMasterXbar__monitor_1__a_first_1  ; 
  assign   tlMasterXbar__monitor_1__a_opcodes_set_interm  =  tlMasterXbar__monitor_1___T_966   ? 4'h9:4'h0; 
  assign   tlMasterXbar__monitor_1___a_opcodes_set_T_1  ={15'b0,  tlMasterXbar__monitor_1__a_opcodes_set_interm  }; 
  assign   tlMasterXbar__monitor_1__a_sizes_set_interm  =  tlMasterXbar__monitor_1___T_966   ? 5'hd:5'h0; 
  assign   tlMasterXbar__monitor_1___a_sizes_set_T_1  ={15'b0,  tlMasterXbar__monitor_1__a_sizes_set_interm  }; 
  assign   tlMasterXbar__monitor_1___T_972  =~  tlMasterXbar__monitor_1__inflight  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___GEN_16  =  tlMasterXbar__monitor_1___T_966   ? 2'h1:2'h0; 
  assign   tlMasterXbar__monitor_1___GEN_19  =  tlMasterXbar__monitor_1___T_966   ?   tlMasterXbar__monitor_1___a_opcodes_set_T_1  :19'h0; 
  assign   tlMasterXbar__monitor_1___GEN_20  =  tlMasterXbar__monitor_1___T_966   ?   tlMasterXbar__monitor_1___a_sizes_set_T_1  :20'h0; 
  assign   tlMasterXbar__monitor_1___T_974  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__d_first_1  ; 
  assign   tlMasterXbar__monitor_1___T_977  =  tlMasterXbar__monitor_1___T_974  &~  tlMasterXbar__monitor_1___T_770  ; 
  assign   tlMasterXbar__monitor_1___GEN_21  =  tlMasterXbar__monitor_1___T_977   ? 2'h1:2'h0; 
  assign   tlMasterXbar__monitor_1___d_opcodes_clr_T_5  ={15'b0,  tlMasterXbar__monitor_1___a_opcode_lookup_T_5  }; 
  assign   tlMasterXbar__monitor_1___d_sizes_clr_T_5  ={15'b0,  tlMasterXbar__monitor_1___a_size_lookup_T_5  }; 
  assign   tlMasterXbar__monitor_1___GEN_23  =  tlMasterXbar__monitor_1___T_977   ?   tlMasterXbar__monitor_1___d_opcodes_clr_T_5  :31'h0; 
  assign   tlMasterXbar__monitor_1___GEN_24  =  tlMasterXbar__monitor_1___T_977   ?   tlMasterXbar__monitor_1___d_sizes_clr_T_5  :31'h0; 
  assign   tlMasterXbar__monitor_1___T_989  =  tlMasterXbar__monitor_1__inflight  |  tlMasterXbar__monitor_1___T_963  ; 
  assign   tlMasterXbar__monitor_1___T_991  =  tlMasterXbar__monitor_1___T_989  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_995  =  tlMasterXbar__monitor_1___T_864  |  tlMasterXbar__monitor_1___T_864  ; 
  assign   tlMasterXbar__monitor_1___T_997  =  tlMasterXbar__monitor_1___T_995  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_999  =4'h6==  tlMasterXbar__monitor_1__io_in_d_bits_size  ; 
  assign   tlMasterXbar__monitor_1___T_1001  =  tlMasterXbar__monitor_1___T_999  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1__a_opcode_lookup  =  tlMasterXbar__monitor_1___a_opcode_lookup_T_7  [3:0]; 
  assign   tlMasterXbar__monitor_1___GEN_43  =3'h2==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h1:3'h0; 
  assign   tlMasterXbar__monitor_1___GEN_44  =3'h3==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h1:  tlMasterXbar__monitor_1___GEN_43  ; 
  assign   tlMasterXbar__monitor_1___GEN_45  =3'h4==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h1:  tlMasterXbar__monitor_1___GEN_44  ; 
  assign   tlMasterXbar__monitor_1___GEN_46  =3'h5==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h2:  tlMasterXbar__monitor_1___GEN_45  ; 
  assign   tlMasterXbar__monitor_1___GEN_47  =3'h6==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h4:  tlMasterXbar__monitor_1___GEN_46  ; 
  assign   tlMasterXbar__monitor_1___GEN_48  =3'h7==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h4:  tlMasterXbar__monitor_1___GEN_47  ; 
  assign   tlMasterXbar__monitor_1___T_1004  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==  tlMasterXbar__monitor_1___GEN_48  ; 
  assign   tlMasterXbar__monitor_1___GEN_55  =3'h6==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h5:  tlMasterXbar__monitor_1___GEN_46  ; 
  assign   tlMasterXbar__monitor_1___GEN_56  =3'h7==  tlMasterXbar__monitor_1__a_opcode_lookup  [2:0] ? 3'h4:  tlMasterXbar__monitor_1___GEN_55  ; 
  assign   tlMasterXbar__monitor_1___T_1006  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==  tlMasterXbar__monitor_1___GEN_56  ; 
  assign   tlMasterXbar__monitor_1___T_1007  =  tlMasterXbar__monitor_1___T_1004  |  tlMasterXbar__monitor_1___T_1006  ; 
  assign   tlMasterXbar__monitor_1___T_1009  =  tlMasterXbar__monitor_1___T_1007  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1__a_size_lookup  =  tlMasterXbar__monitor_1___a_size_lookup_T_7  [7:0]; 
  assign   tlMasterXbar__monitor_1___GEN_75  ={4'b0,  tlMasterXbar__monitor_1__io_in_d_bits_size  }; 
  assign   tlMasterXbar__monitor_1___T_1011  =  tlMasterXbar__monitor_1___GEN_75  ==  tlMasterXbar__monitor_1__a_size_lookup  ; 
  assign   tlMasterXbar__monitor_1___T_1013  =  tlMasterXbar__monitor_1___T_1011  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_1016  =  tlMasterXbar__monitor_1___T_974  &  tlMasterXbar__monitor_1__a_first_1  ; 
  assign   tlMasterXbar__monitor_1___T_1017  =  tlMasterXbar__monitor_1___T_1016  &  tlMasterXbar__monitor_1__io_in_a_valid  ; 
  assign   tlMasterXbar__monitor_1___T_1021  =  tlMasterXbar__monitor_1___T_1017  &~  tlMasterXbar__monitor_1___T_770  ; 
  assign   tlMasterXbar__monitor_1___T_1025  =  tlMasterXbar__monitor_1__io_in_a_ready  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1__a_set_wo_ready  =  tlMasterXbar__monitor_1___GEN_15  [0]; 
  assign   tlMasterXbar__monitor_1__d_clr_wo_ready  =  tlMasterXbar__monitor_1___GEN_21  [0]; 
  assign   tlMasterXbar__monitor_1___T_1027  =  tlMasterXbar__monitor_1__a_set_wo_ready  !=  tlMasterXbar__monitor_1__d_clr_wo_ready  ; 
  assign   tlMasterXbar__monitor_1___T_1028  =|  tlMasterXbar__monitor_1__a_set_wo_ready  ; 
  assign   tlMasterXbar__monitor_1___T_1030  =  tlMasterXbar__monitor_1___T_1027  |~  tlMasterXbar__monitor_1___T_1028  ; 
  assign   tlMasterXbar__monitor_1___T_1032  =  tlMasterXbar__monitor_1___T_1030  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1__a_set  =  tlMasterXbar__monitor_1___GEN_16  [0]; 
  assign   tlMasterXbar__monitor_1___inflight_T  =  tlMasterXbar__monitor_1__inflight  |  tlMasterXbar__monitor_1__a_set  ; 
  assign   tlMasterXbar__monitor_1___inflight_T_2  =  tlMasterXbar__monitor_1___inflight_T  &~  tlMasterXbar__monitor_1__d_clr_wo_ready  ; 
  assign   tlMasterXbar__monitor_1__a_opcodes_set  =  tlMasterXbar__monitor_1___GEN_19  [3:0]; 
  assign   tlMasterXbar__monitor_1___inflight_opcodes_T  =  tlMasterXbar__monitor_1__inflight_opcodes  |  tlMasterXbar__monitor_1__a_opcodes_set  ; 
  assign   tlMasterXbar__monitor_1__d_opcodes_clr  =  tlMasterXbar__monitor_1___GEN_23  [3:0]; 
  assign   tlMasterXbar__monitor_1___inflight_opcodes_T_2  =  tlMasterXbar__monitor_1___inflight_opcodes_T  &~  tlMasterXbar__monitor_1__d_opcodes_clr  ; 
  assign   tlMasterXbar__monitor_1__a_sizes_set  =  tlMasterXbar__monitor_1___GEN_20  [7:0]; 
  assign   tlMasterXbar__monitor_1___inflight_sizes_T  =  tlMasterXbar__monitor_1__inflight_sizes  |  tlMasterXbar__monitor_1__a_sizes_set  ; 
  assign   tlMasterXbar__monitor_1__d_sizes_clr  =  tlMasterXbar__monitor_1___GEN_24  [7:0]; 
  assign   tlMasterXbar__monitor_1___inflight_sizes_T_2  =  tlMasterXbar__monitor_1___inflight_sizes_T  &~  tlMasterXbar__monitor_1__d_sizes_clr  ; 
  assign   tlMasterXbar__monitor_1___T_1034  =|  tlMasterXbar__monitor_1__inflight  ; 
  assign   tlMasterXbar__monitor_1___T_1036  =  tlMasterXbar__monitor_1__plusarg_reader_out  ==32'h0; 
  assign   tlMasterXbar__monitor_1___T_1037  =~  tlMasterXbar__monitor_1___T_1034  |  tlMasterXbar__monitor_1___T_1036  ; 
  assign   tlMasterXbar__monitor_1___T_1038  =  tlMasterXbar__monitor_1__watchdog  <  tlMasterXbar__monitor_1__plusarg_reader_out  ; 
  assign   tlMasterXbar__monitor_1___T_1039  =  tlMasterXbar__monitor_1___T_1037  |  tlMasterXbar__monitor_1___T_1038  ; 
  assign   tlMasterXbar__monitor_1___T_1041  =  tlMasterXbar__monitor_1___T_1039  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___watchdog_T_1  =  tlMasterXbar__monitor_1__watchdog  +32'h1; 
  assign   tlMasterXbar__monitor_1___T_1045  =  tlMasterXbar__monitor_1__a_first_done  |  tlMasterXbar__monitor_1__io_in_d_valid  ; 
  assign   tlMasterXbar__monitor_1__d_first_counter1_2  =  tlMasterXbar__monitor_1__d_first_counter_2  -9'h1; 
  assign   tlMasterXbar__monitor_1__d_first_2  =  tlMasterXbar__monitor_1__d_first_counter_2  ==9'h0; 
  assign   tlMasterXbar__monitor_1___GEN_78  ={8'b0,  tlMasterXbar__monitor_1__inflight_sizes_1  }; 
  assign   tlMasterXbar__monitor_1___c_size_lookup_T_6  =  tlMasterXbar__monitor_1___GEN_78  &  tlMasterXbar__monitor_1___a_size_lookup_T_5  ; 
  assign   tlMasterXbar__monitor_1___c_size_lookup_T_7  ={1'b0,  tlMasterXbar__monitor_1___c_size_lookup_T_6  [15:1]}; 
  assign   tlMasterXbar__monitor_1___T_1063  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__d_first_2  ; 
  assign   tlMasterXbar__monitor_1___T_1065  =  tlMasterXbar__monitor_1___T_1063  &  tlMasterXbar__monitor_1___T_770  ; 
  assign   tlMasterXbar__monitor_1___GEN_66  =  tlMasterXbar__monitor_1___T_1065   ? 2'h1:2'h0; 
  assign   tlMasterXbar__monitor_1___GEN_69  =  tlMasterXbar__monitor_1___T_1065   ?   tlMasterXbar__monitor_1___d_sizes_clr_T_5  :31'h0; 
  assign   tlMasterXbar__monitor_1___T_1077  =  tlMasterXbar__monitor_1__inflight_1  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1__c_size_lookup  =  tlMasterXbar__monitor_1___c_size_lookup_T_7  [7:0]; 
  assign   tlMasterXbar__monitor_1___T_1083  =  tlMasterXbar__monitor_1___GEN_75  ==  tlMasterXbar__monitor_1__c_size_lookup  ; 
  assign   tlMasterXbar__monitor_1___T_1085  =  tlMasterXbar__monitor_1___T_1083  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___T_1098  =|1'h0; 
  assign   tlMasterXbar__monitor_1__d_clr_wo_ready_1  =  tlMasterXbar__monitor_1___GEN_66  [0]; 
  assign   tlMasterXbar__monitor_1___T_1101  =  tlMasterXbar__monitor_1__d_clr_wo_ready_1  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___inflight_T_5  =  tlMasterXbar__monitor_1__inflight_1  &~  tlMasterXbar__monitor_1__d_clr_wo_ready_1  ; 
  assign   tlMasterXbar__monitor_1__d_sizes_clr_1  =  tlMasterXbar__monitor_1___GEN_69  [7:0]; 
  assign   tlMasterXbar__monitor_1___inflight_sizes_T_5  =  tlMasterXbar__monitor_1__inflight_sizes_1  &~  tlMasterXbar__monitor_1__d_sizes_clr_1  ; 
  assign   tlMasterXbar__monitor_1___T_1103  =|  tlMasterXbar__monitor_1__inflight_1  ; 
  assign   tlMasterXbar__monitor_1___T_1105  =  tlMasterXbar__monitor_1__plusarg_reader_1_out  ==32'h0; 
  assign   tlMasterXbar__monitor_1___T_1106  =~  tlMasterXbar__monitor_1___T_1103  |  tlMasterXbar__monitor_1___T_1105  ; 
  assign   tlMasterXbar__monitor_1___T_1107  =  tlMasterXbar__monitor_1__watchdog_1  <  tlMasterXbar__monitor_1__plusarg_reader_1_out  ; 
  assign   tlMasterXbar__monitor_1___T_1108  =  tlMasterXbar__monitor_1___T_1106  |  tlMasterXbar__monitor_1___T_1107  ; 
  assign   tlMasterXbar__monitor_1___T_1110  =  tlMasterXbar__monitor_1___T_1108  |  tlMasterXbar__monitor_1__reset  ; 
  assign   tlMasterXbar__monitor_1___watchdog_T_3  =  tlMasterXbar__monitor_1__watchdog_1  +32'h1; 
  assign   tlMasterXbar__monitor_1___GEN_81  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1___T_770  ; 
  assign   tlMasterXbar__monitor_1___GEN_89  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1___T_790  ; 
  assign   tlMasterXbar__monitor_1___GEN_97  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1___T_818  ; 
  assign   tlMasterXbar__monitor_1___GEN_105  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1___T_847  ; 
  assign   tlMasterXbar__monitor_1___GEN_109  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1___T_864  ; 
  assign   tlMasterXbar__monitor_1___GEN_113  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1___T_882  ; 
  assign   tlMasterXbar__monitor_1___GEN_117  =  tlMasterXbar__monitor_1___T_977  &  tlMasterXbar__monitor_1___T_963  ; 
  assign   tlMasterXbar__monitor_1___GEN_122  =  tlMasterXbar__monitor_1___T_977  &~  tlMasterXbar__monitor_1___T_963  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_covSum  =30'h0; 
  assign   tlMasterXbar__monitor_1__io_covSum  =  tlMasterXbar__monitor_1__TLMonitor_24_covSum  ; 
  assign   tlMasterXbar__monitor_1__stopEn0  =  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1___T_350  ; 
  assign   tlMasterXbar__monitor_1__stopEn1  =  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1___T_134  ; 
  assign   tlMasterXbar__monitor_1__stopEn2  =  tlMasterXbar__monitor_1__io_in_d_valid  &~  tlMasterXbar__monitor_1___T_768  ; 
  assign   tlMasterXbar__monitor_1__stopEn3  =  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_776  ; 
  assign   tlMasterXbar__monitor_1__stopEn4  =  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_780  ; 
  assign   tlMasterXbar__monitor_1__stopEn5  =  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_784  ; 
  assign   tlMasterXbar__monitor_1__stopEn6  =  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_788  ; 
  assign   tlMasterXbar__monitor_1__stopEn7  =  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_776  ; 
  assign   tlMasterXbar__monitor_1__stopEn8  =  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_803  ; 
  assign   tlMasterXbar__monitor_1__stopEn9  =  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_807  ; 
  assign   tlMasterXbar__monitor_1__stopEn10  =  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_784  ; 
  assign   tlMasterXbar__monitor_1__stopEn11  =  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_776  ; 
  assign   tlMasterXbar__monitor_1__stopEn12  =  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_803  ; 
  assign   tlMasterXbar__monitor_1__stopEn13  =  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_807  ; 
  assign   tlMasterXbar__monitor_1__stopEn14  =  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_840  ; 
  assign   tlMasterXbar__monitor_1__stopEn15  =  tlMasterXbar__monitor_1___GEN_105  &~  tlMasterXbar__monitor_1___T_780  ; 
  assign   tlMasterXbar__monitor_1__stopEn16  =  tlMasterXbar__monitor_1___GEN_105  &~  tlMasterXbar__monitor_1___T_784  ; 
  assign   tlMasterXbar__monitor_1__stopEn17  =  tlMasterXbar__monitor_1___GEN_109  &~  tlMasterXbar__monitor_1___T_780  ; 
  assign   tlMasterXbar__monitor_1__stopEn18  =  tlMasterXbar__monitor_1___GEN_109  &~  tlMasterXbar__monitor_1___T_840  ; 
  assign   tlMasterXbar__monitor_1__stopEn19  =  tlMasterXbar__monitor_1___GEN_113  &~  tlMasterXbar__monitor_1___T_780  ; 
  assign   tlMasterXbar__monitor_1__stopEn20  =  tlMasterXbar__monitor_1___GEN_113  &~  tlMasterXbar__monitor_1___T_784  ; 
  assign   tlMasterXbar__monitor_1__stopEn21  =  tlMasterXbar__monitor_1___T_912  &~  tlMasterXbar__monitor_1___T_931  ; 
  assign   tlMasterXbar__monitor_1__stopEn22  =  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_939  ; 
  assign   tlMasterXbar__monitor_1__stopEn23  =  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_943  ; 
  assign   tlMasterXbar__monitor_1__stopEn24  =  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_947  ; 
  assign   tlMasterXbar__monitor_1__stopEn25  =  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_955  ; 
  assign   tlMasterXbar__monitor_1__stopEn26  =  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_959  ; 
  assign   tlMasterXbar__monitor_1__stopEn27  =  tlMasterXbar__monitor_1___T_966  &~  tlMasterXbar__monitor_1___T_972  ; 
  assign   tlMasterXbar__monitor_1__stopEn28  =  tlMasterXbar__monitor_1___T_977  &~  tlMasterXbar__monitor_1___T_991  ; 
  assign   tlMasterXbar__monitor_1__stopEn29  =  tlMasterXbar__monitor_1___GEN_117  &~  tlMasterXbar__monitor_1___T_997  ; 
  assign   tlMasterXbar__monitor_1__stopEn30  =  tlMasterXbar__monitor_1___GEN_117  &~  tlMasterXbar__monitor_1___T_1001  ; 
  assign   tlMasterXbar__monitor_1__stopEn31  =  tlMasterXbar__monitor_1___GEN_122  &~  tlMasterXbar__monitor_1___T_1009  ; 
  assign   tlMasterXbar__monitor_1__stopEn32  =  tlMasterXbar__monitor_1___GEN_122  &~  tlMasterXbar__monitor_1___T_1013  ; 
  assign   tlMasterXbar__monitor_1__stopEn33  =  tlMasterXbar__monitor_1___T_1021  &~  tlMasterXbar__monitor_1___T_1025  ; 
  assign   tlMasterXbar__monitor_1__stopEn34  =~  tlMasterXbar__monitor_1___T_1032  ; 
  assign   tlMasterXbar__monitor_1__stopEn35  =~  tlMasterXbar__monitor_1___T_1041  ; 
  assign   tlMasterXbar__monitor_1__stopEn36  =  tlMasterXbar__monitor_1___T_1065  &~  tlMasterXbar__monitor_1___T_1077  ; 
  assign   tlMasterXbar__monitor_1__stopEn37  =  tlMasterXbar__monitor_1___T_1065  &~  tlMasterXbar__monitor_1___T_1085  ; 
  assign   tlMasterXbar__monitor_1__stopEn38  =  tlMasterXbar__monitor_1___T_1098  &~  tlMasterXbar__monitor_1___T_1101  ; 
  assign   tlMasterXbar__monitor_1__stopEn39  =~  tlMasterXbar__monitor_1___T_1110  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or15  =  tlMasterXbar__monitor_1__stopEn0  |  tlMasterXbar__monitor_1__stopEn1  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or34  =  tlMasterXbar__monitor_1__stopEn3  |  tlMasterXbar__monitor_1__stopEn4  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or16  =  tlMasterXbar__monitor_1__stopEn2  |  tlMasterXbar__monitor_1__TLMonitor_24_or34  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or7  =  tlMasterXbar__monitor_1__TLMonitor_24_or15  |  tlMasterXbar__monitor_1__TLMonitor_24_or16  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or17  =  tlMasterXbar__monitor_1__stopEn5  |  tlMasterXbar__monitor_1__stopEn6  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or38  =  tlMasterXbar__monitor_1__stopEn8  |  tlMasterXbar__monitor_1__stopEn9  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or18  =  tlMasterXbar__monitor_1__stopEn7  |  tlMasterXbar__monitor_1__TLMonitor_24_or38  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or8  =  tlMasterXbar__monitor_1__TLMonitor_24_or17  |  tlMasterXbar__monitor_1__TLMonitor_24_or18  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or3  =  tlMasterXbar__monitor_1__TLMonitor_24_or7  |  tlMasterXbar__monitor_1__TLMonitor_24_or8  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or19  =  tlMasterXbar__monitor_1__stopEn10  |  tlMasterXbar__monitor_1__stopEn11  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or42  =  tlMasterXbar__monitor_1__stopEn13  |  tlMasterXbar__monitor_1__stopEn14  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or20  =  tlMasterXbar__monitor_1__stopEn12  |  tlMasterXbar__monitor_1__TLMonitor_24_or42  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or9  =  tlMasterXbar__monitor_1__TLMonitor_24_or19  |  tlMasterXbar__monitor_1__TLMonitor_24_or20  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or44  =  tlMasterXbar__monitor_1__stopEn16  |  tlMasterXbar__monitor_1__stopEn17  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or21  =  tlMasterXbar__monitor_1__stopEn15  |  tlMasterXbar__monitor_1__TLMonitor_24_or44  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or46  =  tlMasterXbar__monitor_1__stopEn19  |  tlMasterXbar__monitor_1__stopEn20  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or22  =  tlMasterXbar__monitor_1__stopEn18  |  tlMasterXbar__monitor_1__TLMonitor_24_or46  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or10  =  tlMasterXbar__monitor_1__TLMonitor_24_or21  |  tlMasterXbar__monitor_1__TLMonitor_24_or22  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or4  =  tlMasterXbar__monitor_1__TLMonitor_24_or9  |  tlMasterXbar__monitor_1__TLMonitor_24_or10  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or1  =  tlMasterXbar__monitor_1__TLMonitor_24_or3  |  tlMasterXbar__monitor_1__TLMonitor_24_or4  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or23  =  tlMasterXbar__monitor_1__stopEn21  |  tlMasterXbar__monitor_1__stopEn22  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or50  =  tlMasterXbar__monitor_1__stopEn24  |  tlMasterXbar__monitor_1__stopEn25  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or24  =  tlMasterXbar__monitor_1__stopEn23  |  tlMasterXbar__monitor_1__TLMonitor_24_or50  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or11  =  tlMasterXbar__monitor_1__TLMonitor_24_or23  |  tlMasterXbar__monitor_1__TLMonitor_24_or24  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or25  =  tlMasterXbar__monitor_1__stopEn26  |  tlMasterXbar__monitor_1__stopEn27  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or54  =  tlMasterXbar__monitor_1__stopEn29  |  tlMasterXbar__monitor_1__stopEn30  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or26  =  tlMasterXbar__monitor_1__stopEn28  |  tlMasterXbar__monitor_1__TLMonitor_24_or54  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or12  =  tlMasterXbar__monitor_1__TLMonitor_24_or25  |  tlMasterXbar__monitor_1__TLMonitor_24_or26  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or5  =  tlMasterXbar__monitor_1__TLMonitor_24_or11  |  tlMasterXbar__monitor_1__TLMonitor_24_or12  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or27  =  tlMasterXbar__monitor_1__stopEn31  |  tlMasterXbar__monitor_1__stopEn32  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or58  =  tlMasterXbar__monitor_1__stopEn34  |  tlMasterXbar__monitor_1__stopEn35  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or28  =  tlMasterXbar__monitor_1__stopEn33  |  tlMasterXbar__monitor_1__TLMonitor_24_or58  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or13  =  tlMasterXbar__monitor_1__TLMonitor_24_or27  |  tlMasterXbar__monitor_1__TLMonitor_24_or28  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or60  =  tlMasterXbar__monitor_1__stopEn37  |  tlMasterXbar__monitor_1__stopEn38  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or29  =  tlMasterXbar__monitor_1__stopEn36  |  tlMasterXbar__monitor_1__TLMonitor_24_or60  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or62  =  tlMasterXbar__monitor_1__plusarg_reader_metaAssert_wire  |  tlMasterXbar__monitor_1__plusarg_reader_1_metaAssert_wire  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or30  =  tlMasterXbar__monitor_1__stopEn39  |  tlMasterXbar__monitor_1__TLMonitor_24_or62  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or14  =  tlMasterXbar__monitor_1__TLMonitor_24_or29  |  tlMasterXbar__monitor_1__TLMonitor_24_or30  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or6  =  tlMasterXbar__monitor_1__TLMonitor_24_or13  |  tlMasterXbar__monitor_1__TLMonitor_24_or14  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or2  =  tlMasterXbar__monitor_1__TLMonitor_24_or5  |  tlMasterXbar__monitor_1__TLMonitor_24_or6  ; 
  assign   tlMasterXbar__monitor_1__TLMonitor_24_or0  =  tlMasterXbar__monitor_1__TLMonitor_24_or1  |  tlMasterXbar__monitor_1__TLMonitor_24_or2  ; 
  assign   tlMasterXbar__monitor_1__metaAssert  =  tlMasterXbar__monitor_1__TLMonitor_24_metaAssert  ; initial
    begin 
    end  
  always @( posedge   tlMasterXbar__monitor_1__clock  )
       begin 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__a_first_counter   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__a_first_counter   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor_1__a_first_done  )
                  begin 
                    if (  tlMasterXbar__monitor_1__a_first  )
                       begin  
                          tlMasterXbar__monitor_1__a_first_counter   <=9'h0;
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor_1__a_first_counter   <=  tlMasterXbar__monitor_1__a_first_counter1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__address   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1___T_934  )
               begin  
                  tlMasterXbar__monitor_1__address   <=  tlMasterXbar__monitor_1__io_in_a_bits_address  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__d_first_counter   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__d_first_counter   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor_1__io_in_d_valid  )
                  begin 
                    if (  tlMasterXbar__monitor_1__d_first  )
                       begin 
                         if (  tlMasterXbar__monitor_1__d_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor_1__d_first_counter   <=  tlMasterXbar__monitor_1__d_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor_1__d_first_counter   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor_1__d_first_counter   <=  tlMasterXbar__monitor_1__d_first_counter1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__opcode_1   <=3'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1___T_962  )
               begin  
                  tlMasterXbar__monitor_1__opcode_1   <=  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__param_1   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1___T_962  )
               begin  
                  tlMasterXbar__monitor_1__param_1   <=  tlMasterXbar__monitor_1__io_in_d_bits_param  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__size_1   <=4'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1___T_962  )
               begin  
                  tlMasterXbar__monitor_1__size_1   <=  tlMasterXbar__monitor_1__io_in_d_bits_size  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__sink   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1___T_962  )
               begin  
                  tlMasterXbar__monitor_1__sink   <=  tlMasterXbar__monitor_1__io_in_d_bits_sink  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__denied   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1___T_962  )
               begin  
                  tlMasterXbar__monitor_1__denied   <=  tlMasterXbar__monitor_1__io_in_d_bits_denied  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__inflight   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__inflight   <=1'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor_1__inflight   <=  tlMasterXbar__monitor_1___inflight_T_2  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__inflight_opcodes   <=4'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__inflight_opcodes   <=4'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor_1__inflight_opcodes   <=  tlMasterXbar__monitor_1___inflight_opcodes_T_2  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__inflight_sizes   <=8'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__inflight_sizes   <=8'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor_1__inflight_sizes   <=  tlMasterXbar__monitor_1___inflight_sizes_T_2  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__a_first_counter_1   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__a_first_counter_1   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor_1__a_first_done  )
                  begin 
                    if (  tlMasterXbar__monitor_1__a_first_1  )
                       begin  
                          tlMasterXbar__monitor_1__a_first_counter_1   <=9'h0;
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor_1__a_first_counter_1   <=  tlMasterXbar__monitor_1__a_first_counter1_1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__d_first_counter_1   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__d_first_counter_1   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor_1__io_in_d_valid  )
                  begin 
                    if (  tlMasterXbar__monitor_1__d_first_1  )
                       begin 
                         if (  tlMasterXbar__monitor_1__d_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor_1__d_first_counter_1   <=  tlMasterXbar__monitor_1__d_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor_1__d_first_counter_1   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor_1__d_first_counter_1   <=  tlMasterXbar__monitor_1__d_first_counter1_1  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__watchdog   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__watchdog   <=32'h0;
               end 
             else 
               if (  tlMasterXbar__monitor_1___T_1045  )
                  begin  
                     tlMasterXbar__monitor_1__watchdog   <=32'h0;
                  end 
                else 
                  begin  
                     tlMasterXbar__monitor_1__watchdog   <=  tlMasterXbar__monitor_1___watchdog_T_1  ;
                  end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__inflight_1   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__inflight_1   <=1'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor_1__inflight_1   <=  tlMasterXbar__monitor_1___inflight_T_5  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__inflight_sizes_1   <=8'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__inflight_sizes_1   <=8'h0;
               end 
             else 
               begin  
                  tlMasterXbar__monitor_1__inflight_sizes_1   <=  tlMasterXbar__monitor_1___inflight_sizes_T_5  ;
               end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__d_first_counter_2   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__d_first_counter_2   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__monitor_1__io_in_d_valid  )
                  begin 
                    if (  tlMasterXbar__monitor_1__d_first_2  )
                       begin 
                         if (  tlMasterXbar__monitor_1__d_first_beats1_opdata  )
                            begin  
                               tlMasterXbar__monitor_1__d_first_counter_2   <=  tlMasterXbar__monitor_1__d_first_beats1_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__monitor_1__d_first_counter_2   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__monitor_1__d_first_counter_2   <=  tlMasterXbar__monitor_1__d_first_counter1_2  ;
                       end 
                  end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__watchdog_1   <=32'h0;
            end 
          else 
            if (  tlMasterXbar__monitor_1__reset  )
               begin  
                  tlMasterXbar__monitor_1__watchdog_1   <=32'h0;
               end 
             else 
               if (  tlMasterXbar__monitor_1__io_in_d_valid  )
                  begin  
                     tlMasterXbar__monitor_1__watchdog_1   <=32'h0;
                  end 
                else 
                  begin  
                     tlMasterXbar__monitor_1__watchdog_1   <=  tlMasterXbar__monitor_1___watchdog_T_3  ;
                  end 
         if (  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1___T_350  )
            begin $display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1___T_350  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1___T_134  )
            begin $display("Assertion failed: 'A' channel Get address not aligned to size (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1___T_134  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1__io_in_d_valid  &~  tlMasterXbar__monitor_1___T_768  )
            begin $display("Assertion failed: 'D' channel has invalid opcode (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1__io_in_d_valid  &~  tlMasterXbar__monitor_1___T_768  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_776  )
            begin $display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_776  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_788  )
            begin $display("Assertion failed: 'D' channel ReleaseAck is denied (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_81  &~  tlMasterXbar__monitor_1___T_788  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_776  )
            begin $display("Assertion failed: 'D' channel Grant smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_776  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_803  )
            begin $display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_803  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_807  )
            begin $display("Assertion failed: 'D' channel Grant carries toN param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_807  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("Assertion failed: 'D' channel Grant is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_89  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_776  )
            begin $display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_776  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_803  )
            begin $display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_803  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_807  )
            begin $display("Assertion failed: 'D' channel GrantData carries toN param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_807  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_840  )
            begin $display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_97  &~  tlMasterXbar__monitor_1___T_840  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_105  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_105  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_105  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("Assertion failed: 'D' channel AccessAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_105  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_109  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_109  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_109  &~  tlMasterXbar__monitor_1___T_840  )
            begin $display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_109  &~  tlMasterXbar__monitor_1___T_840  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_113  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("Assertion failed: 'D' channel HintAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_113  &~  tlMasterXbar__monitor_1___T_780  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_113  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("Assertion failed: 'D' channel HintAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_113  &~  tlMasterXbar__monitor_1___T_784  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_912  &~  tlMasterXbar__monitor_1___T_931  )
            begin $display("Assertion failed: 'A' channel address changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_912  &~  tlMasterXbar__monitor_1___T_931  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_939  )
            begin $display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_939  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_943  )
            begin $display("Assertion failed: 'D' channel param changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_943  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_947  )
            begin $display("Assertion failed: 'D' channel size changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_947  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_955  )
            begin $display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_955  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_959  )
            begin $display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_936  &~  tlMasterXbar__monitor_1___T_959  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_966  &~  tlMasterXbar__monitor_1___T_972  )
            begin $display("Assertion failed: 'A' channel re-used a source ID (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_966  &~  tlMasterXbar__monitor_1___T_972  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_977  &~  tlMasterXbar__monitor_1___T_991  )
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_977  &~  tlMasterXbar__monitor_1___T_991  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_117  &~  tlMasterXbar__monitor_1___T_997  )
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_117  &~  tlMasterXbar__monitor_1___T_997  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_117  &~  tlMasterXbar__monitor_1___T_1001  )
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_117  &~  tlMasterXbar__monitor_1___T_1001  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_122  &~  tlMasterXbar__monitor_1___T_1009  )
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_122  &~  tlMasterXbar__monitor_1___T_1009  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___GEN_122  &~  tlMasterXbar__monitor_1___T_1013  )
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___GEN_122  &~  tlMasterXbar__monitor_1___T_1013  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_1021  &~  tlMasterXbar__monitor_1___T_1025  )
            begin $display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_1021  &~  tlMasterXbar__monitor_1___T_1025  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar__monitor_1___T_1032  )
            begin $display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (~  tlMasterXbar__monitor_1___T_1032  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar__monitor_1___T_1041  )
            begin $display("Assertion failed: TileLink timeout expired (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~  tlMasterXbar__monitor_1___T_1041  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_1065  &~  tlMasterXbar__monitor_1___T_1077  )
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_1065  &~  tlMasterXbar__monitor_1___T_1077  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_1065  &~  tlMasterXbar__monitor_1___T_1085  )
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_1065  &~  tlMasterXbar__monitor_1___T_1085  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1___T_1098  &~  tlMasterXbar__monitor_1___T_1101  )
            begin $display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (  tlMasterXbar__monitor_1___T_1098  &~  tlMasterXbar__monitor_1___T_1101  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar__monitor_1___T_1110  )
            begin $display("Assertion failed: TileLink timeout expired (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~  tlMasterXbar__monitor_1___T_1110  )
            begin $display("fatal");
            end 
         if (  tlMasterXbar__monitor_1__metaReset  )
            begin  
               tlMasterXbar__monitor_1__TLMonitor_24_metaAssert   <=1'h0;
            end 
          else 
            begin  
               tlMasterXbar__monitor_1__TLMonitor_24_metaAssert   <=  tlMasterXbar__monitor_1__TLMonitor_24_metaAssert  |  tlMasterXbar__monitor_1__TLMonitor_24_or0  ;
            end 
       end
 
assign tlMasterXbar__monitor_1__clock = tlMasterXbar__monitor_1_clock;
assign tlMasterXbar__monitor_1__reset = tlMasterXbar__monitor_1_reset;
assign tlMasterXbar__monitor_1__io_in_a_ready = tlMasterXbar__monitor_1_io_in_a_ready;
assign tlMasterXbar__monitor_1__io_in_a_valid = tlMasterXbar__monitor_1_io_in_a_valid;
assign tlMasterXbar__monitor_1__io_in_a_bits_address = tlMasterXbar__monitor_1_io_in_a_bits_address;
assign tlMasterXbar__monitor_1__io_in_d_valid = tlMasterXbar__monitor_1_io_in_d_valid;
assign tlMasterXbar__monitor_1__io_in_d_bits_opcode = tlMasterXbar__monitor_1_io_in_d_bits_opcode;
assign tlMasterXbar__monitor_1__io_in_d_bits_param = tlMasterXbar__monitor_1_io_in_d_bits_param;
assign tlMasterXbar__monitor_1__io_in_d_bits_size = tlMasterXbar__monitor_1_io_in_d_bits_size;
assign tlMasterXbar__monitor_1__io_in_d_bits_sink = tlMasterXbar__monitor_1_io_in_d_bits_sink;
assign tlMasterXbar__monitor_1__io_in_d_bits_denied = tlMasterXbar__monitor_1_io_in_d_bits_denied;
assign tlMasterXbar__monitor_1__io_in_d_bits_corrupt = tlMasterXbar__monitor_1_io_in_d_bits_corrupt;
assign tlMasterXbar__monitor_1_io_covSum = tlMasterXbar__monitor_1__io_covSum;
assign tlMasterXbar__monitor_1_metaAssert = tlMasterXbar__monitor_1__metaAssert;
assign tlMasterXbar__monitor_1__metaReset = tlMasterXbar__monitor_1_metaReset;
 
  assign   tlMasterXbar__requestBOI_0_0  =~  tlMasterXbar__auto_out_b_bits_source  [1]; 
  assign   tlMasterXbar__requestDOI_0_0  =~  tlMasterXbar__auto_out_d_bits_source  [1]; 
  assign   tlMasterXbar__requestDOI_0_1  =  tlMasterXbar__auto_out_d_bits_source  ==2'h2; 
  assign   tlMasterXbar___beatsAI_decode_T_1  =27'hfff<<  tlMasterXbar__auto_in_0_a_bits_size  ; 
  assign   tlMasterXbar__beatsAI_decode  =~  tlMasterXbar___beatsAI_decode_T_1  [11:3]; 
  assign   tlMasterXbar__beatsAI_opdata  =~  tlMasterXbar__auto_in_0_a_bits_opcode  [2]; 
  assign   tlMasterXbar___portsDIO_out_0_d_ready_T  =  tlMasterXbar__requestDOI_0_0  &  tlMasterXbar__auto_in_0_d_ready  ; 
  assign   tlMasterXbar__idle  =  tlMasterXbar__beatsLeft  ==9'h0; 
  assign   tlMasterXbar__latch  =  tlMasterXbar__idle  &  tlMasterXbar__auto_out_a_ready  ; 
  assign   tlMasterXbar__readys_filter_lo  ={  tlMasterXbar__auto_in_1_a_valid  ,  tlMasterXbar__auto_in_0_a_valid  }; 
  assign   tlMasterXbar___readys_T_1  =  tlMasterXbar__readys_filter_lo  ==  tlMasterXbar__readys_filter_lo  ; 
  assign   tlMasterXbar___readys_T_3  =  tlMasterXbar___readys_T_1  |  tlMasterXbar__reset  ; 
  assign   tlMasterXbar__readys_filter_hi  =  tlMasterXbar__readys_filter_lo  &~  tlMasterXbar__readys_mask  ; 
  assign   tlMasterXbar__readys_filter  ={  tlMasterXbar__readys_filter_hi  ,  tlMasterXbar__auto_in_1_a_valid  ,  tlMasterXbar__auto_in_0_a_valid  }; 
  assign   tlMasterXbar___GEN_1  ={1'b0,  tlMasterXbar__readys_filter  [3:1]}; 
  assign   tlMasterXbar___readys_unready_T_1  =  tlMasterXbar__readys_filter  |  tlMasterXbar___GEN_1  ; 
  assign   tlMasterXbar___readys_unready_T_4  ={  tlMasterXbar__readys_mask  ,2'h0}; 
  assign   tlMasterXbar___GEN_2  ={1'b0,  tlMasterXbar___readys_unready_T_1  [3:1]}; 
  assign   tlMasterXbar__readys_unready  =  tlMasterXbar___GEN_2  |  tlMasterXbar___readys_unready_T_4  ; 
  assign   tlMasterXbar___readys_readys_T_2  =  tlMasterXbar__readys_unready  [3:2]&  tlMasterXbar__readys_unready  [1:0]; 
  assign   tlMasterXbar__readys_readys  =~  tlMasterXbar___readys_readys_T_2  ; 
  assign   tlMasterXbar___readys_T_5  =|  tlMasterXbar__readys_filter_lo  ; 
  assign   tlMasterXbar___readys_T_6  =  tlMasterXbar__latch  &  tlMasterXbar___readys_T_5  ; 
  assign   tlMasterXbar___readys_mask_T  =  tlMasterXbar__readys_readys  &  tlMasterXbar__readys_filter_lo  ; 
  assign   tlMasterXbar___readys_mask_T_1  ={  tlMasterXbar___readys_mask_T  ,1'h0}; 
  assign   tlMasterXbar___readys_mask_T_3  =  tlMasterXbar___readys_mask_T  |  tlMasterXbar___readys_mask_T_1  [1:0]; 
  assign   tlMasterXbar__readys_0  =  tlMasterXbar__readys_readys  [0]; 
  assign   tlMasterXbar__readys_1  =  tlMasterXbar__readys_readys  [1]; 
  assign   tlMasterXbar__earlyWinner_0  =  tlMasterXbar__readys_0  &  tlMasterXbar__auto_in_0_a_valid  ; 
  assign   tlMasterXbar__earlyWinner_1  =  tlMasterXbar__readys_1  &  tlMasterXbar__auto_in_1_a_valid  ; 
  assign   tlMasterXbar___prefixOR_T  =  tlMasterXbar__earlyWinner_0  |  tlMasterXbar__earlyWinner_1  ; 
  assign   tlMasterXbar___T_6  =~  tlMasterXbar__earlyWinner_0  |~  tlMasterXbar__earlyWinner_1  ; 
  assign   tlMasterXbar___T_9  =  tlMasterXbar___T_6  |  tlMasterXbar__reset  ; 
  assign   tlMasterXbar___T_11  =  tlMasterXbar__auto_in_0_a_valid  |  tlMasterXbar__auto_in_1_a_valid  ; 
  assign   tlMasterXbar___T_14  =~  tlMasterXbar___T_11  |  tlMasterXbar___prefixOR_T  ; 
  assign   tlMasterXbar___T_16  =  tlMasterXbar___T_14  |  tlMasterXbar__reset  ; 
  assign   tlMasterXbar___T_21  =~  tlMasterXbar___T_11  |  tlMasterXbar___T_11  ; 
  assign   tlMasterXbar___T_23  =  tlMasterXbar___T_21  |  tlMasterXbar__reset  ; 
  assign   tlMasterXbar__muxStateEarly_0  =  tlMasterXbar__idle   ?   tlMasterXbar__earlyWinner_0  :  tlMasterXbar__state_0  ; 
  assign   tlMasterXbar__muxStateEarly_1  =  tlMasterXbar__idle   ?   tlMasterXbar__earlyWinner_1  :  tlMasterXbar__state_1  ; 
  assign   tlMasterXbar___out_0_a_earlyValid_T_1  =  tlMasterXbar__state_0  &  tlMasterXbar__auto_in_0_a_valid  ; 
  assign   tlMasterXbar___out_0_a_earlyValid_T_2  =  tlMasterXbar__state_1  &  tlMasterXbar__auto_in_1_a_valid  ; 
  assign   tlMasterXbar___out_0_a_earlyValid_T_3  =  tlMasterXbar___out_0_a_earlyValid_T_1  |  tlMasterXbar___out_0_a_earlyValid_T_2  ; 
  assign   tlMasterXbar__out_2_0_a_earlyValid  =  tlMasterXbar__idle   ?   tlMasterXbar___T_11  :  tlMasterXbar___out_0_a_earlyValid_T_3  ; 
  assign   tlMasterXbar___beatsLeft_T_2  =  tlMasterXbar__auto_out_a_ready  &  tlMasterXbar__out_2_0_a_earlyValid  ; 
  assign   tlMasterXbar___GEN_3  ={8'b0,  tlMasterXbar___beatsLeft_T_2  }; 
  assign   tlMasterXbar___beatsLeft_T_4  =  tlMasterXbar__beatsLeft  -  tlMasterXbar___GEN_3  ; 
  assign   tlMasterXbar__allowed_0  =  tlMasterXbar__idle   ?   tlMasterXbar__readys_0  :  tlMasterXbar__state_0  ; 
  assign   tlMasterXbar__allowed_1  =  tlMasterXbar__idle   ?   tlMasterXbar__readys_1  :  tlMasterXbar__state_1  ; 
  assign   tlMasterXbar___T_31  =  tlMasterXbar__muxStateEarly_0   ?   tlMasterXbar__auto_in_0_a_bits_mask  :8'h0; 
  assign   tlMasterXbar___T_32  =  tlMasterXbar__muxStateEarly_1   ? 8'hff:8'h0; 
  assign   tlMasterXbar___T_34  =  tlMasterXbar__muxStateEarly_0   ?   tlMasterXbar__auto_in_0_a_bits_address  :32'h0; 
  assign   tlMasterXbar___T_35  =  tlMasterXbar__muxStateEarly_1   ?   tlMasterXbar__auto_in_1_a_bits_address  :32'h0; 
  assign   tlMasterXbar__in_0_a_bits_source  ={1'b0,  tlMasterXbar__auto_in_0_a_bits_source  }; 
  assign   tlMasterXbar___T_37  =  tlMasterXbar__muxStateEarly_0   ?   tlMasterXbar__in_0_a_bits_source  :2'h0; 
  assign   tlMasterXbar___T_38  =  tlMasterXbar__muxStateEarly_1   ? 2'h2:2'h0; 
  assign   tlMasterXbar___T_40  =  tlMasterXbar__muxStateEarly_0   ?   tlMasterXbar__auto_in_0_a_bits_size  :4'h0; 
  assign   tlMasterXbar___T_41  =  tlMasterXbar__muxStateEarly_1   ? 4'h6:4'h0; 
  assign   tlMasterXbar___T_46  =  tlMasterXbar__muxStateEarly_0   ?   tlMasterXbar__auto_in_0_a_bits_opcode  :3'h0; 
  assign   tlMasterXbar___T_47  =  tlMasterXbar__muxStateEarly_1   ? 3'h4:3'h0; 
  assign   tlMasterXbar__auto_in_1_a_ready  =  tlMasterXbar__auto_out_a_ready  &  tlMasterXbar__allowed_1  ; 
  assign   tlMasterXbar__auto_in_1_d_valid  =  tlMasterXbar__auto_out_d_valid  &  tlMasterXbar__requestDOI_0_1  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_opcode  =  tlMasterXbar__auto_out_d_bits_opcode  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_size  =  tlMasterXbar__auto_out_d_bits_size  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_data  =  tlMasterXbar__auto_out_d_bits_data  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_corrupt  =  tlMasterXbar__auto_out_d_bits_corrupt  ; 
  assign   tlMasterXbar__auto_in_0_a_ready  =  tlMasterXbar__auto_out_a_ready  &  tlMasterXbar__allowed_0  ; 
  assign   tlMasterXbar__auto_in_0_b_valid  =  tlMasterXbar__auto_out_b_valid  &  tlMasterXbar__requestBOI_0_0  ; 
  assign   tlMasterXbar__auto_in_0_b_bits_param  =  tlMasterXbar__auto_out_b_bits_param  ; 
  assign   tlMasterXbar__auto_in_0_b_bits_size  =  tlMasterXbar__auto_out_b_bits_size  ; 
  assign   tlMasterXbar__auto_in_0_b_bits_source  =  tlMasterXbar__auto_out_b_bits_source  [0]; 
  assign   tlMasterXbar__auto_in_0_b_bits_address  =  tlMasterXbar__auto_out_b_bits_address  ; 
  assign   tlMasterXbar__auto_in_0_c_ready  =  tlMasterXbar__auto_out_c_ready  ; 
  assign   tlMasterXbar__auto_in_0_d_valid  =  tlMasterXbar__auto_out_d_valid  &  tlMasterXbar__requestDOI_0_0  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_opcode  =  tlMasterXbar__auto_out_d_bits_opcode  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_param  =  tlMasterXbar__auto_out_d_bits_param  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_size  =  tlMasterXbar__auto_out_d_bits_size  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_source  =  tlMasterXbar__auto_out_d_bits_source  [0]; 
  assign   tlMasterXbar__auto_in_0_d_bits_sink  =  tlMasterXbar__auto_out_d_bits_sink  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_denied  =  tlMasterXbar__auto_out_d_bits_denied  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_data  =  tlMasterXbar__auto_out_d_bits_data  ; 
  assign   tlMasterXbar__auto_in_0_e_ready  =  tlMasterXbar__auto_out_e_ready  ; 
  assign   tlMasterXbar__auto_out_a_valid  =  tlMasterXbar__idle   ?   tlMasterXbar___T_11  :  tlMasterXbar___out_0_a_earlyValid_T_3  ; 
  assign   tlMasterXbar__auto_out_a_bits_opcode  =  tlMasterXbar___T_46  |  tlMasterXbar___T_47  ; 
  assign   tlMasterXbar__auto_out_a_bits_param  =  tlMasterXbar__muxStateEarly_0   ?   tlMasterXbar__auto_in_0_a_bits_param  :3'h0; 
  assign   tlMasterXbar__auto_out_a_bits_size  =  tlMasterXbar___T_40  |  tlMasterXbar___T_41  ; 
  assign   tlMasterXbar__auto_out_a_bits_source  =  tlMasterXbar___T_37  |  tlMasterXbar___T_38  ; 
  assign   tlMasterXbar__auto_out_a_bits_address  =  tlMasterXbar___T_34  |  tlMasterXbar___T_35  ; 
  assign   tlMasterXbar__auto_out_a_bits_mask  =  tlMasterXbar___T_31  |  tlMasterXbar___T_32  ; 
  assign   tlMasterXbar__auto_out_a_bits_data  =  tlMasterXbar__muxStateEarly_0   ?   tlMasterXbar__auto_in_0_a_bits_data  :64'h0; 
  assign   tlMasterXbar__auto_out_b_ready  =  tlMasterXbar__requestBOI_0_0  &  tlMasterXbar__auto_in_0_b_ready  ; 
  assign   tlMasterXbar__auto_out_c_valid  =  tlMasterXbar__auto_in_0_c_valid  ; 
  assign   tlMasterXbar__auto_out_c_bits_opcode  =  tlMasterXbar__auto_in_0_c_bits_opcode  ; 
  assign   tlMasterXbar__auto_out_c_bits_param  =  tlMasterXbar__auto_in_0_c_bits_param  ; 
  assign   tlMasterXbar__auto_out_c_bits_size  =  tlMasterXbar__auto_in_0_c_bits_size  ; 
  assign   tlMasterXbar__auto_out_c_bits_source  ={1'b0,  tlMasterXbar__auto_in_0_c_bits_source  }; 
  assign   tlMasterXbar__auto_out_c_bits_address  =  tlMasterXbar__auto_in_0_c_bits_address  ; 
  assign   tlMasterXbar__auto_out_c_bits_data  =  tlMasterXbar__auto_in_0_c_bits_data  ; 
  assign   tlMasterXbar__auto_out_d_ready  =  tlMasterXbar___portsDIO_out_0_d_ready_T  |  tlMasterXbar__requestDOI_0_1  ; 
  assign   tlMasterXbar__auto_out_e_valid  =  tlMasterXbar__auto_in_0_e_valid  ; 
  assign   tlMasterXbar__auto_out_e_bits_sink  =  tlMasterXbar__auto_in_0_e_bits_sink  ; 
  assign   tlMasterXbar__monitor_clock  =  tlMasterXbar__clock  ; 
  assign   tlMasterXbar__monitor_reset  =  tlMasterXbar__reset  ; 
  assign   tlMasterXbar__monitor_io_in_a_ready  =  tlMasterXbar__auto_out_a_ready  &  tlMasterXbar__allowed_0  ; 
  assign   tlMasterXbar__monitor_io_in_a_valid  =  tlMasterXbar__auto_in_0_a_valid  ; 
  assign   tlMasterXbar__monitor_io_in_a_bits_opcode  =  tlMasterXbar__auto_in_0_a_bits_opcode  ; 
  assign   tlMasterXbar__monitor_io_in_a_bits_param  =  tlMasterXbar__auto_in_0_a_bits_param  ; 
  assign   tlMasterXbar__monitor_io_in_a_bits_size  =  tlMasterXbar__auto_in_0_a_bits_size  ; 
  assign   tlMasterXbar__monitor_io_in_a_bits_source  =  tlMasterXbar__auto_in_0_a_bits_source  ; 
  assign   tlMasterXbar__monitor_io_in_a_bits_address  =  tlMasterXbar__auto_in_0_a_bits_address  ; 
  assign   tlMasterXbar__monitor_io_in_a_bits_mask  =  tlMasterXbar__auto_in_0_a_bits_mask  ; 
  assign   tlMasterXbar__monitor_io_in_b_ready  =  tlMasterXbar__auto_in_0_b_ready  ; 
  assign   tlMasterXbar__monitor_io_in_b_valid  =  tlMasterXbar__auto_out_b_valid  &  tlMasterXbar__requestBOI_0_0  ; 
  assign   tlMasterXbar__monitor_io_in_b_bits_opcode  =  tlMasterXbar__auto_out_b_bits_opcode  ; 
  assign   tlMasterXbar__monitor_io_in_b_bits_param  =  tlMasterXbar__auto_out_b_bits_param  ; 
  assign   tlMasterXbar__monitor_io_in_b_bits_size  =  tlMasterXbar__auto_out_b_bits_size  ; 
  assign   tlMasterXbar__monitor_io_in_b_bits_source  =  tlMasterXbar__auto_out_b_bits_source  [0]; 
  assign   tlMasterXbar__monitor_io_in_b_bits_address  =  tlMasterXbar__auto_out_b_bits_address  ; 
  assign   tlMasterXbar__monitor_io_in_b_bits_mask  =  tlMasterXbar__auto_out_b_bits_mask  ; 
  assign   tlMasterXbar__monitor_io_in_b_bits_corrupt  =  tlMasterXbar__auto_out_b_bits_corrupt  ; 
  assign   tlMasterXbar__monitor_io_in_c_ready  =  tlMasterXbar__auto_out_c_ready  ; 
  assign   tlMasterXbar__monitor_io_in_c_valid  =  tlMasterXbar__auto_in_0_c_valid  ; 
  assign   tlMasterXbar__monitor_io_in_c_bits_opcode  =  tlMasterXbar__auto_in_0_c_bits_opcode  ; 
  assign   tlMasterXbar__monitor_io_in_c_bits_param  =  tlMasterXbar__auto_in_0_c_bits_param  ; 
  assign   tlMasterXbar__monitor_io_in_c_bits_size  =  tlMasterXbar__auto_in_0_c_bits_size  ; 
  assign   tlMasterXbar__monitor_io_in_c_bits_source  =  tlMasterXbar__auto_in_0_c_bits_source  ; 
  assign   tlMasterXbar__monitor_io_in_c_bits_address  =  tlMasterXbar__auto_in_0_c_bits_address  ; 
  assign   tlMasterXbar__monitor_io_in_d_ready  =  tlMasterXbar__auto_in_0_d_ready  ; 
  assign   tlMasterXbar__monitor_io_in_d_valid  =  tlMasterXbar__auto_out_d_valid  &  tlMasterXbar__requestDOI_0_0  ; 
  assign   tlMasterXbar__monitor_io_in_d_bits_opcode  =  tlMasterXbar__auto_out_d_bits_opcode  ; 
  assign   tlMasterXbar__monitor_io_in_d_bits_param  =  tlMasterXbar__auto_out_d_bits_param  ; 
  assign   tlMasterXbar__monitor_io_in_d_bits_size  =  tlMasterXbar__auto_out_d_bits_size  ; 
  assign   tlMasterXbar__monitor_io_in_d_bits_source  =  tlMasterXbar__auto_out_d_bits_source  [0]; 
  assign   tlMasterXbar__monitor_io_in_d_bits_sink  =  tlMasterXbar__auto_out_d_bits_sink  ; 
  assign   tlMasterXbar__monitor_io_in_d_bits_denied  =  tlMasterXbar__auto_out_d_bits_denied  ; 
  assign   tlMasterXbar__monitor_io_in_d_bits_corrupt  =  tlMasterXbar__auto_out_d_bits_corrupt  ; 
  assign   tlMasterXbar__monitor_io_in_e_ready  =  tlMasterXbar__auto_out_e_ready  ; 
  assign   tlMasterXbar__monitor_io_in_e_valid  =  tlMasterXbar__auto_in_0_e_valid  ; 
  assign   tlMasterXbar__monitor_io_in_e_bits_sink  =  tlMasterXbar__auto_in_0_e_bits_sink  ; 
  assign   tlMasterXbar__monitor_1_clock  =  tlMasterXbar__clock  ; 
  assign   tlMasterXbar__monitor_1_reset  =  tlMasterXbar__reset  ; 
  assign   tlMasterXbar__monitor_1_io_in_a_ready  =  tlMasterXbar__auto_out_a_ready  &  tlMasterXbar__allowed_1  ; 
  assign   tlMasterXbar__monitor_1_io_in_a_valid  =  tlMasterXbar__auto_in_1_a_valid  ; 
  assign   tlMasterXbar__monitor_1_io_in_a_bits_address  =  tlMasterXbar__auto_in_1_a_bits_address  ; 
  assign   tlMasterXbar__monitor_1_io_in_d_valid  =  tlMasterXbar__auto_out_d_valid  &  tlMasterXbar__requestDOI_0_1  ; 
  assign   tlMasterXbar__monitor_1_io_in_d_bits_opcode  =  tlMasterXbar__auto_out_d_bits_opcode  ; 
  assign   tlMasterXbar__monitor_1_io_in_d_bits_param  =  tlMasterXbar__auto_out_d_bits_param  ; 
  assign   tlMasterXbar__monitor_1_io_in_d_bits_size  =  tlMasterXbar__auto_out_d_bits_size  ; 
  assign   tlMasterXbar__monitor_1_io_in_d_bits_sink  =  tlMasterXbar__auto_out_d_bits_sink  ; 
  assign   tlMasterXbar__monitor_1_io_in_d_bits_denied  =  tlMasterXbar__auto_out_d_bits_denied  ; 
  assign   tlMasterXbar__monitor_1_io_in_d_bits_corrupt  =  tlMasterXbar__auto_out_d_bits_corrupt  ; 
  assign   tlMasterXbar__TLXbar_7_cov_read_addr  =  tlMasterXbar__TLXbar_7_state  ; 
  assign   tlMasterXbar__TLXbar_7_cov_read_data  =  tlMasterXbar__TLXbar_7_cov  [  tlMasterXbar__TLXbar_7_cov_read_addr  ]; 
  assign   tlMasterXbar__TLXbar_7_cov_write_data  =1'h1; 
  assign   tlMasterXbar__TLXbar_7_cov_write_addr  =  tlMasterXbar__TLXbar_7_state  ; 
  assign   tlMasterXbar__TLXbar_7_cov_write_mask  =1'h1; 
  assign   tlMasterXbar__TLXbar_7_cov_write_en  =1'h1; 
  assign   tlMasterXbar__readys_mask_shl  =  tlMasterXbar__readys_mask  ; 
  assign   tlMasterXbar__readys_mask_pad  ={1'h0,  tlMasterXbar__readys_mask_shl  }; 
  assign   tlMasterXbar__state_0_shl  ={  tlMasterXbar__state_0  ,2'h0}; 
  assign   tlMasterXbar__state_0_pad  =  tlMasterXbar__state_0_shl  ; 
  assign   tlMasterXbar__state_1_shl  ={  tlMasterXbar__state_1  ,2'h0}; 
  assign   tlMasterXbar__state_1_pad  =  tlMasterXbar__state_1_shl  ; 
  assign   tlMasterXbar__TLXbar_7_xor2  =  tlMasterXbar__state_0_pad  ^  tlMasterXbar__state_1_pad  ; 
  assign   tlMasterXbar__TLXbar_7_xor0  =  tlMasterXbar__readys_mask_pad  ^  tlMasterXbar__TLXbar_7_xor2  ; 
  assign   tlMasterXbar__monitor_sum  =  tlMasterXbar__TLXbar_7_covSum  +  tlMasterXbar__monitor_io_covSum  ; 
  assign   tlMasterXbar__monitor_1_sum  =  tlMasterXbar__monitor_sum  +  tlMasterXbar__monitor_1_io_covSum  ; 
  assign   tlMasterXbar__io_covSum  =  tlMasterXbar__monitor_1_sum  ; 
  assign   tlMasterXbar__stopEn0  =~  tlMasterXbar___readys_T_3  ; 
  assign   tlMasterXbar__stopEn1  =~  tlMasterXbar___T_9  ; 
  assign   tlMasterXbar__stopEn2  =~  tlMasterXbar___T_16  ; 
  assign   tlMasterXbar__stopEn3  =~  tlMasterXbar___T_23  ; 
  assign   tlMasterXbar__monitor_metaAssert_wire  =  tlMasterXbar__monitor_metaAssert  ; 
  assign   tlMasterXbar__monitor_1_metaAssert_wire  =  tlMasterXbar__monitor_1_metaAssert  ; 
  assign   tlMasterXbar__TLXbar_7_or4  =  tlMasterXbar__stopEn1  |  tlMasterXbar__stopEn2  ; 
  assign   tlMasterXbar__TLXbar_7_or1  =  tlMasterXbar__stopEn0  |  tlMasterXbar__TLXbar_7_or4  ; 
  assign   tlMasterXbar__TLXbar_7_or6  =  tlMasterXbar__monitor_metaAssert_wire  |  tlMasterXbar__monitor_1_metaAssert_wire  ; 
  assign   tlMasterXbar__TLXbar_7_or2  =  tlMasterXbar__stopEn3  |  tlMasterXbar__TLXbar_7_or6  ; 
  assign   tlMasterXbar__TLXbar_7_or0  =  tlMasterXbar__TLXbar_7_or1  |  tlMasterXbar__TLXbar_7_or2  ; 
  assign   tlMasterXbar__metaAssert  =  tlMasterXbar__TLXbar_7_metaAssert  ; 
  assign   tlMasterXbar__monitor_metaReset  =  tlMasterXbar__metaReset  |  tlMasterXbar__monitor_halt  ; 
  assign   tlMasterXbar__monitor_1_metaReset  =  tlMasterXbar__metaReset  |  tlMasterXbar__monitor_1_halt  ; initial
    begin 
    end  
  always @( posedge   tlMasterXbar__clock  )
       begin 
         if (  tlMasterXbar__metaReset  )
            begin  
               tlMasterXbar__beatsLeft   <=9'h0;
            end 
          else 
            if (  tlMasterXbar__reset  )
               begin  
                  tlMasterXbar__beatsLeft   <=9'h0;
               end 
             else 
               if (  tlMasterXbar__latch  )
                  begin 
                    if (  tlMasterXbar__earlyWinner_0  )
                       begin 
                         if (  tlMasterXbar__beatsAI_opdata  )
                            begin  
                               tlMasterXbar__beatsLeft   <=  tlMasterXbar__beatsAI_decode  ;
                            end 
                          else 
                            begin  
                               tlMasterXbar__beatsLeft   <=9'h0;
                            end 
                       end 
                     else 
                       begin  
                          tlMasterXbar__beatsLeft   <=9'h0;
                       end 
                  end 
                else 
                  begin  
                     tlMasterXbar__beatsLeft   <=  tlMasterXbar___beatsLeft_T_4  ;
                  end 
         if (  tlMasterXbar__metaReset  )
            begin  
               tlMasterXbar__readys_mask   <=2'h0;
            end 
          else 
            if (  tlMasterXbar__reset  )
               begin  
                  tlMasterXbar__readys_mask   <=2'h3;
               end 
             else 
               if (  tlMasterXbar___readys_T_6  )
                  begin  
                     tlMasterXbar__readys_mask   <=  tlMasterXbar___readys_mask_T_3  ;
                  end 
         if (  tlMasterXbar__metaReset  )
            begin  
               tlMasterXbar__state_0   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__reset  )
               begin  
                  tlMasterXbar__state_0   <=1'h0;
               end 
             else 
               if (  tlMasterXbar__idle  )
                  begin  
                     tlMasterXbar__state_0   <=  tlMasterXbar__earlyWinner_0  ;
                  end 
         if (  tlMasterXbar__metaReset  )
            begin  
               tlMasterXbar__state_1   <=1'h0;
            end 
          else 
            if (  tlMasterXbar__reset  )
               begin  
                  tlMasterXbar__state_1   <=1'h0;
               end 
             else 
               if (  tlMasterXbar__idle  )
                  begin  
                     tlMasterXbar__state_1   <=  tlMasterXbar__earlyWinner_1  ;
                  end 
         if (~  tlMasterXbar___readys_T_3  )
            begin $display("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");
            end 
         if (~  tlMasterXbar___readys_T_3  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar___T_9  )
            begin $display("Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
            end 
         if (~  tlMasterXbar___T_9  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar___T_16  )
            begin $display("Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n");
            end 
         if (~  tlMasterXbar___T_16  )
            begin $display("fatal");
            end 
         if (~  tlMasterXbar___T_23  )
            begin $display("Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n");
            end 
         if (~  tlMasterXbar___T_23  )
            begin $display("fatal");
            end  
          tlMasterXbar__TLXbar_7_state   <=  tlMasterXbar__TLXbar_7_xor0  ;
         if (!(  tlMasterXbar__TLXbar_7_cov_read_data  ))
            begin  
               tlMasterXbar__TLXbar_7_covSum   <=  tlMasterXbar__TLXbar_7_covSum  +1'h1;
            end 
         if (  tlMasterXbar__metaReset  )
            begin  
               tlMasterXbar__TLXbar_7_metaAssert   <=1'h0;
            end 
          else 
            begin  
               tlMasterXbar__TLXbar_7_metaAssert   <=  tlMasterXbar__TLXbar_7_metaAssert  |  tlMasterXbar__TLXbar_7_or0  ;
            end 
       end
  
  always @( posedge   tlMasterXbar__clock  )
       begin 
         if (  tlMasterXbar__TLXbar_7_cov_write_en  &  tlMasterXbar__TLXbar_7_cov_write_mask  )
            begin  
               tlMasterXbar__TLXbar_7_cov   [  tlMasterXbar__TLXbar_7_cov_write_addr  ]<=  tlMasterXbar__TLXbar_7_cov_write_data  ;
            end 
       end
 
assign tlMasterXbar__clock = tlMasterXbar_clock;
assign tlMasterXbar__reset = tlMasterXbar_reset;
assign tlMasterXbar_auto_in_1_a_ready = tlMasterXbar__auto_in_1_a_ready;
assign tlMasterXbar__auto_in_1_a_valid = tlMasterXbar_auto_in_1_a_valid;
assign tlMasterXbar__auto_in_1_a_bits_address = tlMasterXbar_auto_in_1_a_bits_address;
assign tlMasterXbar_auto_in_1_d_valid = tlMasterXbar__auto_in_1_d_valid;
assign tlMasterXbar_auto_in_1_d_bits_opcode = tlMasterXbar__auto_in_1_d_bits_opcode;
assign tlMasterXbar_auto_in_1_d_bits_size = tlMasterXbar__auto_in_1_d_bits_size;
assign tlMasterXbar_auto_in_1_d_bits_data = tlMasterXbar__auto_in_1_d_bits_data;
assign tlMasterXbar_auto_in_1_d_bits_corrupt = tlMasterXbar__auto_in_1_d_bits_corrupt;
assign tlMasterXbar_auto_in_0_a_ready = tlMasterXbar__auto_in_0_a_ready;
assign tlMasterXbar__auto_in_0_a_valid = tlMasterXbar_auto_in_0_a_valid;
assign tlMasterXbar__auto_in_0_a_bits_opcode = tlMasterXbar_auto_in_0_a_bits_opcode;
assign tlMasterXbar__auto_in_0_a_bits_param = tlMasterXbar_auto_in_0_a_bits_param;
assign tlMasterXbar__auto_in_0_a_bits_size = tlMasterXbar_auto_in_0_a_bits_size;
assign tlMasterXbar__auto_in_0_a_bits_source = tlMasterXbar_auto_in_0_a_bits_source;
assign tlMasterXbar__auto_in_0_a_bits_address = tlMasterXbar_auto_in_0_a_bits_address;
assign tlMasterXbar__auto_in_0_a_bits_mask = tlMasterXbar_auto_in_0_a_bits_mask;
assign tlMasterXbar__auto_in_0_a_bits_data = tlMasterXbar_auto_in_0_a_bits_data;
assign tlMasterXbar__auto_in_0_b_ready = tlMasterXbar_auto_in_0_b_ready;
assign tlMasterXbar_auto_in_0_b_valid = tlMasterXbar__auto_in_0_b_valid;
assign tlMasterXbar_auto_in_0_b_bits_param = tlMasterXbar__auto_in_0_b_bits_param;
assign tlMasterXbar_auto_in_0_b_bits_size = tlMasterXbar__auto_in_0_b_bits_size;
assign tlMasterXbar_auto_in_0_b_bits_source = tlMasterXbar__auto_in_0_b_bits_source;
assign tlMasterXbar_auto_in_0_b_bits_address = tlMasterXbar__auto_in_0_b_bits_address;
assign tlMasterXbar_auto_in_0_c_ready = tlMasterXbar__auto_in_0_c_ready;
assign tlMasterXbar__auto_in_0_c_valid = tlMasterXbar_auto_in_0_c_valid;
assign tlMasterXbar__auto_in_0_c_bits_opcode = tlMasterXbar_auto_in_0_c_bits_opcode;
assign tlMasterXbar__auto_in_0_c_bits_param = tlMasterXbar_auto_in_0_c_bits_param;
assign tlMasterXbar__auto_in_0_c_bits_size = tlMasterXbar_auto_in_0_c_bits_size;
assign tlMasterXbar__auto_in_0_c_bits_source = tlMasterXbar_auto_in_0_c_bits_source;
assign tlMasterXbar__auto_in_0_c_bits_address = tlMasterXbar_auto_in_0_c_bits_address;
assign tlMasterXbar__auto_in_0_c_bits_data = tlMasterXbar_auto_in_0_c_bits_data;
assign tlMasterXbar__auto_in_0_d_ready = tlMasterXbar_auto_in_0_d_ready;
assign tlMasterXbar_auto_in_0_d_valid = tlMasterXbar__auto_in_0_d_valid;
assign tlMasterXbar_auto_in_0_d_bits_opcode = tlMasterXbar__auto_in_0_d_bits_opcode;
assign tlMasterXbar_auto_in_0_d_bits_param = tlMasterXbar__auto_in_0_d_bits_param;
assign tlMasterXbar_auto_in_0_d_bits_size = tlMasterXbar__auto_in_0_d_bits_size;
assign tlMasterXbar_auto_in_0_d_bits_source = tlMasterXbar__auto_in_0_d_bits_source;
assign tlMasterXbar_auto_in_0_d_bits_sink = tlMasterXbar__auto_in_0_d_bits_sink;
assign tlMasterXbar_auto_in_0_d_bits_denied = tlMasterXbar__auto_in_0_d_bits_denied;
assign tlMasterXbar_auto_in_0_d_bits_data = tlMasterXbar__auto_in_0_d_bits_data;
assign tlMasterXbar_auto_in_0_e_ready = tlMasterXbar__auto_in_0_e_ready;
assign tlMasterXbar__auto_in_0_e_valid = tlMasterXbar_auto_in_0_e_valid;
assign tlMasterXbar__auto_in_0_e_bits_sink = tlMasterXbar_auto_in_0_e_bits_sink;
assign tlMasterXbar__auto_out_a_ready = tlMasterXbar_auto_out_a_ready;
assign tlMasterXbar_auto_out_a_valid = tlMasterXbar__auto_out_a_valid;
assign tlMasterXbar_auto_out_a_bits_opcode = tlMasterXbar__auto_out_a_bits_opcode;
assign tlMasterXbar_auto_out_a_bits_param = tlMasterXbar__auto_out_a_bits_param;
assign tlMasterXbar_auto_out_a_bits_size = tlMasterXbar__auto_out_a_bits_size;
assign tlMasterXbar_auto_out_a_bits_source = tlMasterXbar__auto_out_a_bits_source;
assign tlMasterXbar_auto_out_a_bits_address = tlMasterXbar__auto_out_a_bits_address;
assign tlMasterXbar_auto_out_a_bits_mask = tlMasterXbar__auto_out_a_bits_mask;
assign tlMasterXbar_auto_out_a_bits_data = tlMasterXbar__auto_out_a_bits_data;
assign tlMasterXbar_auto_out_b_ready = tlMasterXbar__auto_out_b_ready;
assign tlMasterXbar__auto_out_b_valid = tlMasterXbar_auto_out_b_valid;
assign tlMasterXbar__auto_out_b_bits_opcode = tlMasterXbar_auto_out_b_bits_opcode;
assign tlMasterXbar__auto_out_b_bits_param = tlMasterXbar_auto_out_b_bits_param;
assign tlMasterXbar__auto_out_b_bits_size = tlMasterXbar_auto_out_b_bits_size;
assign tlMasterXbar__auto_out_b_bits_source = tlMasterXbar_auto_out_b_bits_source;
assign tlMasterXbar__auto_out_b_bits_address = tlMasterXbar_auto_out_b_bits_address;
assign tlMasterXbar__auto_out_b_bits_mask = tlMasterXbar_auto_out_b_bits_mask;
assign tlMasterXbar__auto_out_b_bits_corrupt = tlMasterXbar_auto_out_b_bits_corrupt;
assign tlMasterXbar__auto_out_c_ready = tlMasterXbar_auto_out_c_ready;
assign tlMasterXbar_auto_out_c_valid = tlMasterXbar__auto_out_c_valid;
assign tlMasterXbar_auto_out_c_bits_opcode = tlMasterXbar__auto_out_c_bits_opcode;
assign tlMasterXbar_auto_out_c_bits_param = tlMasterXbar__auto_out_c_bits_param;
assign tlMasterXbar_auto_out_c_bits_size = tlMasterXbar__auto_out_c_bits_size;
assign tlMasterXbar_auto_out_c_bits_source = tlMasterXbar__auto_out_c_bits_source;
assign tlMasterXbar_auto_out_c_bits_address = tlMasterXbar__auto_out_c_bits_address;
assign tlMasterXbar_auto_out_c_bits_data = tlMasterXbar__auto_out_c_bits_data;
assign tlMasterXbar_auto_out_d_ready = tlMasterXbar__auto_out_d_ready;
assign tlMasterXbar__auto_out_d_valid = tlMasterXbar_auto_out_d_valid;
assign tlMasterXbar__auto_out_d_bits_opcode = tlMasterXbar_auto_out_d_bits_opcode;
assign tlMasterXbar__auto_out_d_bits_param = tlMasterXbar_auto_out_d_bits_param;
assign tlMasterXbar__auto_out_d_bits_size = tlMasterXbar_auto_out_d_bits_size;
assign tlMasterXbar__auto_out_d_bits_source = tlMasterXbar_auto_out_d_bits_source;
assign tlMasterXbar__auto_out_d_bits_sink = tlMasterXbar_auto_out_d_bits_sink;
assign tlMasterXbar__auto_out_d_bits_denied = tlMasterXbar_auto_out_d_bits_denied;
assign tlMasterXbar__auto_out_d_bits_data = tlMasterXbar_auto_out_d_bits_data;
assign tlMasterXbar__auto_out_d_bits_corrupt = tlMasterXbar_auto_out_d_bits_corrupt;
assign tlMasterXbar__auto_out_e_ready = tlMasterXbar_auto_out_e_ready;
assign tlMasterXbar_auto_out_e_valid = tlMasterXbar__auto_out_e_valid;
assign tlMasterXbar_auto_out_e_bits_sink = tlMasterXbar__auto_out_e_bits_sink;
assign tlMasterXbar_io_covSum = tlMasterXbar__io_covSum;
assign tlMasterXbar_metaAssert = tlMasterXbar__metaAssert;
assign tlMasterXbar__metaReset = tlMasterXbar_metaReset;
assign tlMasterXbar__monitor_halt = tlMasterXbar_monitor_halt;
assign tlMasterXbar__monitor_1_halt = tlMasterXbar_monitor_1_halt;
 
  
wire  intXbar__auto_int_in_3_0;
wire  intXbar__auto_int_in_2_0;
wire  intXbar__auto_int_in_1_0;
wire  intXbar__auto_int_in_1_1;
wire  intXbar__auto_int_in_0_0;
wire  intXbar__auto_int_out_0;
wire  intXbar__auto_int_out_1;
wire  intXbar__auto_int_out_2;
wire  intXbar__auto_int_out_3;
wire  intXbar__auto_int_out_4;
wire [29:0] intXbar__io_covSum;
wire  intXbar__metaAssert;
 
   wire[29:0]  intXbar__IntXbar_1_covSum  ; 
  assign   intXbar__auto_int_out_0  =  intXbar__auto_int_in_0_0  ; 
  assign   intXbar__auto_int_out_1  =  intXbar__auto_int_in_1_0  ; 
  assign   intXbar__auto_int_out_2  =  intXbar__auto_int_in_1_1  ; 
  assign   intXbar__auto_int_out_3  =  intXbar__auto_int_in_2_0  ; 
  assign   intXbar__auto_int_out_4  =  intXbar__auto_int_in_3_0  ; 
  assign   intXbar__IntXbar_1_covSum  =30'h0; 
  assign   intXbar__io_covSum  =  intXbar__IntXbar_1_covSum  ; 
  assign   intXbar__metaAssert  =1'h0;
assign intXbar__auto_int_in_3_0 = intXbar_auto_int_in_3_0;
assign intXbar__auto_int_in_2_0 = intXbar_auto_int_in_2_0;
assign intXbar__auto_int_in_1_0 = intXbar_auto_int_in_1_0;
assign intXbar__auto_int_in_1_1 = intXbar_auto_int_in_1_1;
assign intXbar__auto_int_in_0_0 = intXbar_auto_int_in_0_0;
assign intXbar_auto_int_out_0 = intXbar__auto_int_out_0;
assign intXbar_auto_int_out_1 = intXbar__auto_int_out_1;
assign intXbar_auto_int_out_2 = intXbar__auto_int_out_2;
assign intXbar_auto_int_out_3 = intXbar__auto_int_out_3;
assign intXbar_auto_int_out_4 = intXbar__auto_int_out_4;
assign intXbar_io_covSum = intXbar__io_covSum;
assign intXbar_metaAssert = intXbar__metaAssert;
 
  BundleBridgeNexus_6 broadcast(.auto_in(broadcast_auto_in),.auto_out(broadcast_auto_out),.io_covSum(broadcast_io_covSum),.metaAssert(broadcast_metaAssert)); 
  BundleBridgeNexus_7 broadcast_1(.auto_in(broadcast_1_auto_in),.auto_out_1(broadcast_1_auto_out_1),.io_covSum(broadcast_1_io_covSum),.metaAssert(broadcast_1_metaAssert)); 
  BundleBridgeNexus_10 broadcast_3(.auto_in_0_valid(broadcast_3_auto_in_0_valid),.auto_in_0_iaddr(broadcast_3_auto_in_0_iaddr),.auto_in_0_insn(broadcast_3_auto_in_0_insn),.auto_in_0_priv(broadcast_3_auto_in_0_priv),.auto_in_0_exception(broadcast_3_auto_in_0_exception),.auto_in_0_interrupt(broadcast_3_auto_in_0_interrupt),.auto_in_0_cause(broadcast_3_auto_in_0_cause),.auto_in_0_tval(broadcast_3_auto_in_0_tval),.auto_out_0_valid(broadcast_3_auto_out_0_valid),.auto_out_0_iaddr(broadcast_3_auto_out_0_iaddr),.auto_out_0_insn(broadcast_3_auto_out_0_insn),.auto_out_0_priv(broadcast_3_auto_out_0_priv),.auto_out_0_exception(broadcast_3_auto_out_0_exception),.auto_out_0_interrupt(broadcast_3_auto_out_0_interrupt),.auto_out_0_cause(broadcast_3_auto_out_0_cause),.auto_out_0_tval(broadcast_3_auto_out_0_tval),.io_covSum(broadcast_3_io_covSum),.metaAssert(broadcast_3_metaAssert)); 
  DCache dcache(.gated_clock(dcache_gated_clock),.reset(dcache_reset),.auto_out_a_ready(dcache_auto_out_a_ready),.auto_out_a_valid(dcache_auto_out_a_valid),.auto_out_a_bits_opcode(dcache_auto_out_a_bits_opcode),.auto_out_a_bits_param(dcache_auto_out_a_bits_param),.auto_out_a_bits_size(dcache_auto_out_a_bits_size),.auto_out_a_bits_source(dcache_auto_out_a_bits_source),.auto_out_a_bits_address(dcache_auto_out_a_bits_address),.auto_out_a_bits_mask(dcache_auto_out_a_bits_mask),.auto_out_a_bits_data(dcache_auto_out_a_bits_data),.auto_out_b_ready(dcache_auto_out_b_ready),.auto_out_b_valid(dcache_auto_out_b_valid),.auto_out_b_bits_param(dcache_auto_out_b_bits_param),.auto_out_b_bits_size(dcache_auto_out_b_bits_size),.auto_out_b_bits_source(dcache_auto_out_b_bits_source),.auto_out_b_bits_address(dcache_auto_out_b_bits_address),.auto_out_c_ready(dcache_auto_out_c_ready),.auto_out_c_valid(dcache_auto_out_c_valid),.auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),.auto_out_c_bits_param(dcache_auto_out_c_bits_param),.auto_out_c_bits_size(dcache_auto_out_c_bits_size),.auto_out_c_bits_source(dcache_auto_out_c_bits_source),.auto_out_c_bits_address(dcache_auto_out_c_bits_address),.auto_out_c_bits_data(dcache_auto_out_c_bits_data),.auto_out_d_ready(dcache_auto_out_d_ready),.auto_out_d_valid(dcache_auto_out_d_valid),.auto_out_d_bits_opcode(dcache_auto_out_d_bits_opcode),.auto_out_d_bits_param(dcache_auto_out_d_bits_param),.auto_out_d_bits_size(dcache_auto_out_d_bits_size),.auto_out_d_bits_source(dcache_auto_out_d_bits_source),.auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),.auto_out_d_bits_denied(dcache_auto_out_d_bits_denied),.auto_out_d_bits_data(dcache_auto_out_d_bits_data),.auto_out_e_ready(dcache_auto_out_e_ready),.auto_out_e_valid(dcache_auto_out_e_valid),.auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),.io_cpu_req_ready(dcache_io_cpu_req_ready),.io_cpu_req_valid(dcache_io_cpu_req_valid),.io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),.io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),.io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),.io_cpu_req_bits_size(dcache_io_cpu_req_bits_size),.io_cpu_req_bits_signed(dcache_io_cpu_req_bits_signed),.io_cpu_req_bits_phys(dcache_io_cpu_req_bits_phys),.io_cpu_s1_kill(dcache_io_cpu_s1_kill),.io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),.io_cpu_s2_nack(dcache_io_cpu_s2_nack),.io_cpu_resp_valid(dcache_io_cpu_resp_valid),.io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),.io_cpu_resp_bits_size(dcache_io_cpu_resp_bits_size),.io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),.io_cpu_resp_bits_replay(dcache_io_cpu_resp_bits_replay),.io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),.io_cpu_resp_bits_data_word_bypass(dcache_io_cpu_resp_bits_data_word_bypass),.io_cpu_replay_next(dcache_io_cpu_replay_next),.io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),.io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),.io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),.io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),.io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),.io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),.io_cpu_ordered(dcache_io_cpu_ordered),.io_cpu_perf_release(dcache_io_cpu_perf_release),.io_cpu_perf_grant(dcache_io_cpu_perf_grant),.io_ptw_req_ready(dcache_io_ptw_req_ready),.io_ptw_req_valid(dcache_io_ptw_req_valid),.io_ptw_req_bits_bits_addr(dcache_io_ptw_req_bits_bits_addr),.io_ptw_resp_valid(dcache_io_ptw_resp_valid),.io_ptw_resp_bits_ae(dcache_io_ptw_resp_bits_ae),.io_ptw_resp_bits_pte_ppn(dcache_io_ptw_resp_bits_pte_ppn),.io_ptw_resp_bits_pte_d(dcache_io_ptw_resp_bits_pte_d),.io_ptw_resp_bits_pte_a(dcache_io_ptw_resp_bits_pte_a),.io_ptw_resp_bits_pte_g(dcache_io_ptw_resp_bits_pte_g),.io_ptw_resp_bits_pte_u(dcache_io_ptw_resp_bits_pte_u),.io_ptw_resp_bits_pte_x(dcache_io_ptw_resp_bits_pte_x),.io_ptw_resp_bits_pte_w(dcache_io_ptw_resp_bits_pte_w),.io_ptw_resp_bits_pte_r(dcache_io_ptw_resp_bits_pte_r),.io_ptw_resp_bits_pte_v(dcache_io_ptw_resp_bits_pte_v),.io_ptw_resp_bits_level(dcache_io_ptw_resp_bits_level),.io_ptw_resp_bits_homogeneous(dcache_io_ptw_resp_bits_homogeneous),.io_ptw_ptbr_mode(dcache_io_ptw_ptbr_mode),.io_ptw_status_debug(dcache_io_ptw_status_debug),.io_ptw_status_dprv(dcache_io_ptw_status_dprv),.io_ptw_status_mxr(dcache_io_ptw_status_mxr),.io_ptw_status_sum(dcache_io_ptw_status_sum),.io_ptw_pmp_0_cfg_l(dcache_io_ptw_pmp_0_cfg_l),.io_ptw_pmp_0_cfg_a(dcache_io_ptw_pmp_0_cfg_a),.io_ptw_pmp_0_cfg_x(dcache_io_ptw_pmp_0_cfg_x),.io_ptw_pmp_0_cfg_w(dcache_io_ptw_pmp_0_cfg_w),.io_ptw_pmp_0_cfg_r(dcache_io_ptw_pmp_0_cfg_r),.io_ptw_pmp_0_addr(dcache_io_ptw_pmp_0_addr),.io_ptw_pmp_0_mask(dcache_io_ptw_pmp_0_mask),.io_ptw_pmp_1_cfg_l(dcache_io_ptw_pmp_1_cfg_l),.io_ptw_pmp_1_cfg_a(dcache_io_ptw_pmp_1_cfg_a),.io_ptw_pmp_1_cfg_x(dcache_io_ptw_pmp_1_cfg_x),.io_ptw_pmp_1_cfg_w(dcache_io_ptw_pmp_1_cfg_w),.io_ptw_pmp_1_cfg_r(dcache_io_ptw_pmp_1_cfg_r),.io_ptw_pmp_1_addr(dcache_io_ptw_pmp_1_addr),.io_ptw_pmp_1_mask(dcache_io_ptw_pmp_1_mask),.io_ptw_pmp_2_cfg_l(dcache_io_ptw_pmp_2_cfg_l),.io_ptw_pmp_2_cfg_a(dcache_io_ptw_pmp_2_cfg_a),.io_ptw_pmp_2_cfg_x(dcache_io_ptw_pmp_2_cfg_x),.io_ptw_pmp_2_cfg_w(dcache_io_ptw_pmp_2_cfg_w),.io_ptw_pmp_2_cfg_r(dcache_io_ptw_pmp_2_cfg_r),.io_ptw_pmp_2_addr(dcache_io_ptw_pmp_2_addr),.io_ptw_pmp_2_mask(dcache_io_ptw_pmp_2_mask),.io_ptw_pmp_3_cfg_l(dcache_io_ptw_pmp_3_cfg_l),.io_ptw_pmp_3_cfg_a(dcache_io_ptw_pmp_3_cfg_a),.io_ptw_pmp_3_cfg_x(dcache_io_ptw_pmp_3_cfg_x),.io_ptw_pmp_3_cfg_w(dcache_io_ptw_pmp_3_cfg_w),.io_ptw_pmp_3_cfg_r(dcache_io_ptw_pmp_3_cfg_r),.io_ptw_pmp_3_addr(dcache_io_ptw_pmp_3_addr),.io_ptw_pmp_3_mask(dcache_io_ptw_pmp_3_mask),.io_ptw_pmp_4_cfg_l(dcache_io_ptw_pmp_4_cfg_l),.io_ptw_pmp_4_cfg_a(dcache_io_ptw_pmp_4_cfg_a),.io_ptw_pmp_4_cfg_x(dcache_io_ptw_pmp_4_cfg_x),.io_ptw_pmp_4_cfg_w(dcache_io_ptw_pmp_4_cfg_w),.io_ptw_pmp_4_cfg_r(dcache_io_ptw_pmp_4_cfg_r),.io_ptw_pmp_4_addr(dcache_io_ptw_pmp_4_addr),.io_ptw_pmp_4_mask(dcache_io_ptw_pmp_4_mask),.io_ptw_pmp_5_cfg_l(dcache_io_ptw_pmp_5_cfg_l),.io_ptw_pmp_5_cfg_a(dcache_io_ptw_pmp_5_cfg_a),.io_ptw_pmp_5_cfg_x(dcache_io_ptw_pmp_5_cfg_x),.io_ptw_pmp_5_cfg_w(dcache_io_ptw_pmp_5_cfg_w),.io_ptw_pmp_5_cfg_r(dcache_io_ptw_pmp_5_cfg_r),.io_ptw_pmp_5_addr(dcache_io_ptw_pmp_5_addr),.io_ptw_pmp_5_mask(dcache_io_ptw_pmp_5_mask),.io_ptw_pmp_6_cfg_l(dcache_io_ptw_pmp_6_cfg_l),.io_ptw_pmp_6_cfg_a(dcache_io_ptw_pmp_6_cfg_a),.io_ptw_pmp_6_cfg_x(dcache_io_ptw_pmp_6_cfg_x),.io_ptw_pmp_6_cfg_w(dcache_io_ptw_pmp_6_cfg_w),.io_ptw_pmp_6_cfg_r(dcache_io_ptw_pmp_6_cfg_r),.io_ptw_pmp_6_addr(dcache_io_ptw_pmp_6_addr),.io_ptw_pmp_6_mask(dcache_io_ptw_pmp_6_mask),.io_ptw_pmp_7_cfg_l(dcache_io_ptw_pmp_7_cfg_l),.io_ptw_pmp_7_cfg_a(dcache_io_ptw_pmp_7_cfg_a),.io_ptw_pmp_7_cfg_x(dcache_io_ptw_pmp_7_cfg_x),.io_ptw_pmp_7_cfg_w(dcache_io_ptw_pmp_7_cfg_w),.io_ptw_pmp_7_cfg_r(dcache_io_ptw_pmp_7_cfg_r),.io_ptw_pmp_7_addr(dcache_io_ptw_pmp_7_addr),.io_ptw_pmp_7_mask(dcache_io_ptw_pmp_7_mask),.io_covSum(dcache_io_covSum),.metaAssert(dcache_metaAssert),.metaReset(dcache_metaReset),.data_halt(dcache_data_halt),.tlb_halt(dcache_tlb_halt),.pma_checker_halt(dcache_pma_checker_halt),.lfsr_prng_halt(dcache_lfsr_prng_halt)); 
  Frontend frontend(.gated_clock(frontend_gated_clock),.reset(frontend_reset),.auto_icache_master_out_a_ready(frontend_auto_icache_master_out_a_ready),.auto_icache_master_out_a_valid(frontend_auto_icache_master_out_a_valid),.auto_icache_master_out_a_bits_address(frontend_auto_icache_master_out_a_bits_address),.auto_icache_master_out_d_valid(frontend_auto_icache_master_out_d_valid),.auto_icache_master_out_d_bits_opcode(frontend_auto_icache_master_out_d_bits_opcode),.auto_icache_master_out_d_bits_size(frontend_auto_icache_master_out_d_bits_size),.auto_icache_master_out_d_bits_data(frontend_auto_icache_master_out_d_bits_data),.auto_icache_master_out_d_bits_corrupt(frontend_auto_icache_master_out_d_bits_corrupt),.auto_reset_vector_sink_in(frontend_auto_reset_vector_sink_in),.io_cpu_might_request(frontend_io_cpu_might_request),.io_cpu_req_valid(frontend_io_cpu_req_valid),.io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),.io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),.io_cpu_sfence_valid(frontend_io_cpu_sfence_valid),.io_cpu_sfence_bits_rs1(frontend_io_cpu_sfence_bits_rs1),.io_cpu_sfence_bits_rs2(frontend_io_cpu_sfence_bits_rs2),.io_cpu_sfence_bits_addr(frontend_io_cpu_sfence_bits_addr),.io_cpu_resp_ready(frontend_io_cpu_resp_ready),.io_cpu_resp_valid(frontend_io_cpu_resp_valid),.io_cpu_resp_bits_btb_taken(frontend_io_cpu_resp_bits_btb_taken),.io_cpu_resp_bits_btb_bridx(frontend_io_cpu_resp_bits_btb_bridx),.io_cpu_resp_bits_btb_entry(frontend_io_cpu_resp_bits_btb_entry),.io_cpu_resp_bits_btb_bht_history(frontend_io_cpu_resp_bits_btb_bht_history),.io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),.io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),.io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),.io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),.io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),.io_cpu_btb_update_valid(frontend_io_cpu_btb_update_valid),.io_cpu_btb_update_bits_prediction_entry(frontend_io_cpu_btb_update_bits_prediction_entry),.io_cpu_btb_update_bits_pc(frontend_io_cpu_btb_update_bits_pc),.io_cpu_btb_update_bits_isValid(frontend_io_cpu_btb_update_bits_isValid),.io_cpu_btb_update_bits_br_pc(frontend_io_cpu_btb_update_bits_br_pc),.io_cpu_btb_update_bits_cfiType(frontend_io_cpu_btb_update_bits_cfiType),.io_cpu_bht_update_valid(frontend_io_cpu_bht_update_valid),.io_cpu_bht_update_bits_prediction_history(frontend_io_cpu_bht_update_bits_prediction_history),.io_cpu_bht_update_bits_pc(frontend_io_cpu_bht_update_bits_pc),.io_cpu_bht_update_bits_branch(frontend_io_cpu_bht_update_bits_branch),.io_cpu_bht_update_bits_taken(frontend_io_cpu_bht_update_bits_taken),.io_cpu_bht_update_bits_mispredict(frontend_io_cpu_bht_update_bits_mispredict),.io_cpu_flush_icache(frontend_io_cpu_flush_icache),.io_cpu_npc(frontend_io_cpu_npc),.io_ptw_req_ready(frontend_io_ptw_req_ready),.io_ptw_req_valid(frontend_io_ptw_req_valid),.io_ptw_req_bits_valid(frontend_io_ptw_req_bits_valid),.io_ptw_req_bits_bits_addr(frontend_io_ptw_req_bits_bits_addr),.io_ptw_resp_valid(frontend_io_ptw_resp_valid),.io_ptw_resp_bits_ae(frontend_io_ptw_resp_bits_ae),.io_ptw_resp_bits_pte_ppn(frontend_io_ptw_resp_bits_pte_ppn),.io_ptw_resp_bits_pte_d(frontend_io_ptw_resp_bits_pte_d),.io_ptw_resp_bits_pte_a(frontend_io_ptw_resp_bits_pte_a),.io_ptw_resp_bits_pte_g(frontend_io_ptw_resp_bits_pte_g),.io_ptw_resp_bits_pte_u(frontend_io_ptw_resp_bits_pte_u),.io_ptw_resp_bits_pte_x(frontend_io_ptw_resp_bits_pte_x),.io_ptw_resp_bits_pte_w(frontend_io_ptw_resp_bits_pte_w),.io_ptw_resp_bits_pte_r(frontend_io_ptw_resp_bits_pte_r),.io_ptw_resp_bits_pte_v(frontend_io_ptw_resp_bits_pte_v),.io_ptw_resp_bits_level(frontend_io_ptw_resp_bits_level),.io_ptw_resp_bits_homogeneous(frontend_io_ptw_resp_bits_homogeneous),.io_ptw_ptbr_mode(frontend_io_ptw_ptbr_mode),.io_ptw_status_debug(frontend_io_ptw_status_debug),.io_ptw_status_prv(frontend_io_ptw_status_prv),.io_ptw_pmp_0_cfg_l(frontend_io_ptw_pmp_0_cfg_l),.io_ptw_pmp_0_cfg_a(frontend_io_ptw_pmp_0_cfg_a),.io_ptw_pmp_0_cfg_x(frontend_io_ptw_pmp_0_cfg_x),.io_ptw_pmp_0_cfg_w(frontend_io_ptw_pmp_0_cfg_w),.io_ptw_pmp_0_cfg_r(frontend_io_ptw_pmp_0_cfg_r),.io_ptw_pmp_0_addr(frontend_io_ptw_pmp_0_addr),.io_ptw_pmp_0_mask(frontend_io_ptw_pmp_0_mask),.io_ptw_pmp_1_cfg_l(frontend_io_ptw_pmp_1_cfg_l),.io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),.io_ptw_pmp_1_cfg_x(frontend_io_ptw_pmp_1_cfg_x),.io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),.io_ptw_pmp_1_cfg_r(frontend_io_ptw_pmp_1_cfg_r),.io_ptw_pmp_1_addr(frontend_io_ptw_pmp_1_addr),.io_ptw_pmp_1_mask(frontend_io_ptw_pmp_1_mask),.io_ptw_pmp_2_cfg_l(frontend_io_ptw_pmp_2_cfg_l),.io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),.io_ptw_pmp_2_cfg_x(frontend_io_ptw_pmp_2_cfg_x),.io_ptw_pmp_2_cfg_w(frontend_io_ptw_pmp_2_cfg_w),.io_ptw_pmp_2_cfg_r(frontend_io_ptw_pmp_2_cfg_r),.io_ptw_pmp_2_addr(frontend_io_ptw_pmp_2_addr),.io_ptw_pmp_2_mask(frontend_io_ptw_pmp_2_mask),.io_ptw_pmp_3_cfg_l(frontend_io_ptw_pmp_3_cfg_l),.io_ptw_pmp_3_cfg_a(frontend_io_ptw_pmp_3_cfg_a),.io_ptw_pmp_3_cfg_x(frontend_io_ptw_pmp_3_cfg_x),.io_ptw_pmp_3_cfg_w(frontend_io_ptw_pmp_3_cfg_w),.io_ptw_pmp_3_cfg_r(frontend_io_ptw_pmp_3_cfg_r),.io_ptw_pmp_3_addr(frontend_io_ptw_pmp_3_addr),.io_ptw_pmp_3_mask(frontend_io_ptw_pmp_3_mask),.io_ptw_pmp_4_cfg_l(frontend_io_ptw_pmp_4_cfg_l),.io_ptw_pmp_4_cfg_a(frontend_io_ptw_pmp_4_cfg_a),.io_ptw_pmp_4_cfg_x(frontend_io_ptw_pmp_4_cfg_x),.io_ptw_pmp_4_cfg_w(frontend_io_ptw_pmp_4_cfg_w),.io_ptw_pmp_4_cfg_r(frontend_io_ptw_pmp_4_cfg_r),.io_ptw_pmp_4_addr(frontend_io_ptw_pmp_4_addr),.io_ptw_pmp_4_mask(frontend_io_ptw_pmp_4_mask),.io_ptw_pmp_5_cfg_l(frontend_io_ptw_pmp_5_cfg_l),.io_ptw_pmp_5_cfg_a(frontend_io_ptw_pmp_5_cfg_a),.io_ptw_pmp_5_cfg_x(frontend_io_ptw_pmp_5_cfg_x),.io_ptw_pmp_5_cfg_w(frontend_io_ptw_pmp_5_cfg_w),.io_ptw_pmp_5_cfg_r(frontend_io_ptw_pmp_5_cfg_r),.io_ptw_pmp_5_addr(frontend_io_ptw_pmp_5_addr),.io_ptw_pmp_5_mask(frontend_io_ptw_pmp_5_mask),.io_ptw_pmp_6_cfg_l(frontend_io_ptw_pmp_6_cfg_l),.io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),.io_ptw_pmp_6_cfg_x(frontend_io_ptw_pmp_6_cfg_x),.io_ptw_pmp_6_cfg_w(frontend_io_ptw_pmp_6_cfg_w),.io_ptw_pmp_6_cfg_r(frontend_io_ptw_pmp_6_cfg_r),.io_ptw_pmp_6_addr(frontend_io_ptw_pmp_6_addr),.io_ptw_pmp_6_mask(frontend_io_ptw_pmp_6_mask),.io_ptw_pmp_7_cfg_l(frontend_io_ptw_pmp_7_cfg_l),.io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),.io_ptw_pmp_7_cfg_x(frontend_io_ptw_pmp_7_cfg_x),.io_ptw_pmp_7_cfg_w(frontend_io_ptw_pmp_7_cfg_w),.io_ptw_pmp_7_cfg_r(frontend_io_ptw_pmp_7_cfg_r),.io_ptw_pmp_7_addr(frontend_io_ptw_pmp_7_addr),.io_ptw_pmp_7_mask(frontend_io_ptw_pmp_7_mask),.io_ptw_customCSRs_csrs_0_value(frontend_io_ptw_customCSRs_csrs_0_value),.io_covSum(frontend_io_covSum),.metaAssert(frontend_metaAssert),.metaReset(frontend_metaReset),.icache_halt(frontend_icache_halt),.fq_halt(frontend_fq_halt),.tlb_halt(frontend_tlb_halt),.btb_halt(frontend_btb_halt)); 
  FPU fpuOpt(.clock(fpuOpt_clock),.reset(fpuOpt_reset),.io_inst(fpuOpt_io_inst),.io_fromint_data(fpuOpt_io_fromint_data),.io_fcsr_rm(fpuOpt_io_fcsr_rm),.io_fcsr_flags_valid(fpuOpt_io_fcsr_flags_valid),.io_fcsr_flags_bits(fpuOpt_io_fcsr_flags_bits),.io_store_data(fpuOpt_io_store_data),.io_toint_data(fpuOpt_io_toint_data),.io_dmem_resp_val(fpuOpt_io_dmem_resp_val),.io_dmem_resp_type(fpuOpt_io_dmem_resp_type),.io_dmem_resp_tag(fpuOpt_io_dmem_resp_tag),.io_dmem_resp_data(fpuOpt_io_dmem_resp_data),.io_valid(fpuOpt_io_valid),.io_fcsr_rdy(fpuOpt_io_fcsr_rdy),.io_nack_mem(fpuOpt_io_nack_mem),.io_illegal_rm(fpuOpt_io_illegal_rm),.io_killx(fpuOpt_io_killx),.io_killm(fpuOpt_io_killm),.io_dec_wen(fpuOpt_io_dec_wen),.io_dec_ren1(fpuOpt_io_dec_ren1),.io_dec_ren2(fpuOpt_io_dec_ren2),.io_dec_ren3(fpuOpt_io_dec_ren3),.io_sboard_set(fpuOpt_io_sboard_set),.io_sboard_clr(fpuOpt_io_sboard_clr),.io_sboard_clra(fpuOpt_io_sboard_clra),.io_covSum(fpuOpt_io_covSum),.metaAssert(fpuOpt_metaAssert),.metaReset(fpuOpt_metaReset),.fpiu_halt(fpuOpt_fpiu_halt),.ifpu_halt(fpuOpt_ifpu_halt),.sfma_halt(fpuOpt_sfma_halt),.fpmu_halt(fpuOpt_fpmu_halt),.divSqrt_1_halt(fpuOpt_divSqrt_1_halt),.dfma_halt(fpuOpt_dfma_halt),.divSqrt_halt(fpuOpt_divSqrt_halt)); 
  HellaCacheArbiter dcacheArb(.clock(dcacheArb_clock),.io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),.io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),.io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),.io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),.io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),.io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),.io_requestor_0_resp_bits_data(dcacheArb_io_requestor_0_resp_bits_data),.io_requestor_0_s2_xcpt_ae_ld(dcacheArb_io_requestor_0_s2_xcpt_ae_ld),.io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),.io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),.io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),.io_requestor_1_req_bits_tag(dcacheArb_io_requestor_1_req_bits_tag),.io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),.io_requestor_1_req_bits_size(dcacheArb_io_requestor_1_req_bits_size),.io_requestor_1_req_bits_signed(dcacheArb_io_requestor_1_req_bits_signed),.io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),.io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),.io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),.io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),.io_requestor_1_resp_bits_tag(dcacheArb_io_requestor_1_resp_bits_tag),.io_requestor_1_resp_bits_size(dcacheArb_io_requestor_1_resp_bits_size),.io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),.io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),.io_requestor_1_resp_bits_has_data(dcacheArb_io_requestor_1_resp_bits_has_data),.io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),.io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),.io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),.io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),.io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),.io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),.io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),.io_requestor_1_s2_xcpt_ae_st(dcacheArb_io_requestor_1_s2_xcpt_ae_st),.io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),.io_requestor_1_perf_release(dcacheArb_io_requestor_1_perf_release),.io_requestor_1_perf_grant(dcacheArb_io_requestor_1_perf_grant),.io_mem_req_ready(dcacheArb_io_mem_req_ready),.io_mem_req_valid(dcacheArb_io_mem_req_valid),.io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),.io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),.io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),.io_mem_req_bits_size(dcacheArb_io_mem_req_bits_size),.io_mem_req_bits_signed(dcacheArb_io_mem_req_bits_signed),.io_mem_req_bits_phys(dcacheArb_io_mem_req_bits_phys),.io_mem_s1_kill(dcacheArb_io_mem_s1_kill),.io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),.io_mem_s2_nack(dcacheArb_io_mem_s2_nack),.io_mem_resp_valid(dcacheArb_io_mem_resp_valid),.io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),.io_mem_resp_bits_size(dcacheArb_io_mem_resp_bits_size),.io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),.io_mem_resp_bits_replay(dcacheArb_io_mem_resp_bits_replay),.io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),.io_mem_resp_bits_data_word_bypass(dcacheArb_io_mem_resp_bits_data_word_bypass),.io_mem_replay_next(dcacheArb_io_mem_replay_next),.io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),.io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),.io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),.io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),.io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),.io_mem_s2_xcpt_ae_st(dcacheArb_io_mem_s2_xcpt_ae_st),.io_mem_ordered(dcacheArb_io_mem_ordered),.io_mem_perf_release(dcacheArb_io_mem_perf_release),.io_mem_perf_grant(dcacheArb_io_mem_perf_grant),.io_covSum(dcacheArb_io_covSum),.metaAssert(dcacheArb_metaAssert),.metaReset(dcacheArb_metaReset)); 
  PTW ptw(.clock(ptw_clock),.reset(ptw_reset),.io_requestor_0_req_ready(ptw_io_requestor_0_req_ready),.io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),.io_requestor_0_req_bits_bits_addr(ptw_io_requestor_0_req_bits_bits_addr),.io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),.io_requestor_0_resp_bits_ae(ptw_io_requestor_0_resp_bits_ae),.io_requestor_0_resp_bits_pte_ppn(ptw_io_requestor_0_resp_bits_pte_ppn),.io_requestor_0_resp_bits_pte_d(ptw_io_requestor_0_resp_bits_pte_d),.io_requestor_0_resp_bits_pte_a(ptw_io_requestor_0_resp_bits_pte_a),.io_requestor_0_resp_bits_pte_g(ptw_io_requestor_0_resp_bits_pte_g),.io_requestor_0_resp_bits_pte_u(ptw_io_requestor_0_resp_bits_pte_u),.io_requestor_0_resp_bits_pte_x(ptw_io_requestor_0_resp_bits_pte_x),.io_requestor_0_resp_bits_pte_w(ptw_io_requestor_0_resp_bits_pte_w),.io_requestor_0_resp_bits_pte_r(ptw_io_requestor_0_resp_bits_pte_r),.io_requestor_0_resp_bits_pte_v(ptw_io_requestor_0_resp_bits_pte_v),.io_requestor_0_resp_bits_level(ptw_io_requestor_0_resp_bits_level),.io_requestor_0_resp_bits_homogeneous(ptw_io_requestor_0_resp_bits_homogeneous),.io_requestor_0_ptbr_mode(ptw_io_requestor_0_ptbr_mode),.io_requestor_0_status_debug(ptw_io_requestor_0_status_debug),.io_requestor_0_status_dprv(ptw_io_requestor_0_status_dprv),.io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),.io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),.io_requestor_0_pmp_0_cfg_l(ptw_io_requestor_0_pmp_0_cfg_l),.io_requestor_0_pmp_0_cfg_a(ptw_io_requestor_0_pmp_0_cfg_a),.io_requestor_0_pmp_0_cfg_x(ptw_io_requestor_0_pmp_0_cfg_x),.io_requestor_0_pmp_0_cfg_w(ptw_io_requestor_0_pmp_0_cfg_w),.io_requestor_0_pmp_0_cfg_r(ptw_io_requestor_0_pmp_0_cfg_r),.io_requestor_0_pmp_0_addr(ptw_io_requestor_0_pmp_0_addr),.io_requestor_0_pmp_0_mask(ptw_io_requestor_0_pmp_0_mask),.io_requestor_0_pmp_1_cfg_l(ptw_io_requestor_0_pmp_1_cfg_l),.io_requestor_0_pmp_1_cfg_a(ptw_io_requestor_0_pmp_1_cfg_a),.io_requestor_0_pmp_1_cfg_x(ptw_io_requestor_0_pmp_1_cfg_x),.io_requestor_0_pmp_1_cfg_w(ptw_io_requestor_0_pmp_1_cfg_w),.io_requestor_0_pmp_1_cfg_r(ptw_io_requestor_0_pmp_1_cfg_r),.io_requestor_0_pmp_1_addr(ptw_io_requestor_0_pmp_1_addr),.io_requestor_0_pmp_1_mask(ptw_io_requestor_0_pmp_1_mask),.io_requestor_0_pmp_2_cfg_l(ptw_io_requestor_0_pmp_2_cfg_l),.io_requestor_0_pmp_2_cfg_a(ptw_io_requestor_0_pmp_2_cfg_a),.io_requestor_0_pmp_2_cfg_x(ptw_io_requestor_0_pmp_2_cfg_x),.io_requestor_0_pmp_2_cfg_w(ptw_io_requestor_0_pmp_2_cfg_w),.io_requestor_0_pmp_2_cfg_r(ptw_io_requestor_0_pmp_2_cfg_r),.io_requestor_0_pmp_2_addr(ptw_io_requestor_0_pmp_2_addr),.io_requestor_0_pmp_2_mask(ptw_io_requestor_0_pmp_2_mask),.io_requestor_0_pmp_3_cfg_l(ptw_io_requestor_0_pmp_3_cfg_l),.io_requestor_0_pmp_3_cfg_a(ptw_io_requestor_0_pmp_3_cfg_a),.io_requestor_0_pmp_3_cfg_x(ptw_io_requestor_0_pmp_3_cfg_x),.io_requestor_0_pmp_3_cfg_w(ptw_io_requestor_0_pmp_3_cfg_w),.io_requestor_0_pmp_3_cfg_r(ptw_io_requestor_0_pmp_3_cfg_r),.io_requestor_0_pmp_3_addr(ptw_io_requestor_0_pmp_3_addr),.io_requestor_0_pmp_3_mask(ptw_io_requestor_0_pmp_3_mask),.io_requestor_0_pmp_4_cfg_l(ptw_io_requestor_0_pmp_4_cfg_l),.io_requestor_0_pmp_4_cfg_a(ptw_io_requestor_0_pmp_4_cfg_a),.io_requestor_0_pmp_4_cfg_x(ptw_io_requestor_0_pmp_4_cfg_x),.io_requestor_0_pmp_4_cfg_w(ptw_io_requestor_0_pmp_4_cfg_w),.io_requestor_0_pmp_4_cfg_r(ptw_io_requestor_0_pmp_4_cfg_r),.io_requestor_0_pmp_4_addr(ptw_io_requestor_0_pmp_4_addr),.io_requestor_0_pmp_4_mask(ptw_io_requestor_0_pmp_4_mask),.io_requestor_0_pmp_5_cfg_l(ptw_io_requestor_0_pmp_5_cfg_l),.io_requestor_0_pmp_5_cfg_a(ptw_io_requestor_0_pmp_5_cfg_a),.io_requestor_0_pmp_5_cfg_x(ptw_io_requestor_0_pmp_5_cfg_x),.io_requestor_0_pmp_5_cfg_w(ptw_io_requestor_0_pmp_5_cfg_w),.io_requestor_0_pmp_5_cfg_r(ptw_io_requestor_0_pmp_5_cfg_r),.io_requestor_0_pmp_5_addr(ptw_io_requestor_0_pmp_5_addr),.io_requestor_0_pmp_5_mask(ptw_io_requestor_0_pmp_5_mask),.io_requestor_0_pmp_6_cfg_l(ptw_io_requestor_0_pmp_6_cfg_l),.io_requestor_0_pmp_6_cfg_a(ptw_io_requestor_0_pmp_6_cfg_a),.io_requestor_0_pmp_6_cfg_x(ptw_io_requestor_0_pmp_6_cfg_x),.io_requestor_0_pmp_6_cfg_w(ptw_io_requestor_0_pmp_6_cfg_w),.io_requestor_0_pmp_6_cfg_r(ptw_io_requestor_0_pmp_6_cfg_r),.io_requestor_0_pmp_6_addr(ptw_io_requestor_0_pmp_6_addr),.io_requestor_0_pmp_6_mask(ptw_io_requestor_0_pmp_6_mask),.io_requestor_0_pmp_7_cfg_l(ptw_io_requestor_0_pmp_7_cfg_l),.io_requestor_0_pmp_7_cfg_a(ptw_io_requestor_0_pmp_7_cfg_a),.io_requestor_0_pmp_7_cfg_x(ptw_io_requestor_0_pmp_7_cfg_x),.io_requestor_0_pmp_7_cfg_w(ptw_io_requestor_0_pmp_7_cfg_w),.io_requestor_0_pmp_7_cfg_r(ptw_io_requestor_0_pmp_7_cfg_r),.io_requestor_0_pmp_7_addr(ptw_io_requestor_0_pmp_7_addr),.io_requestor_0_pmp_7_mask(ptw_io_requestor_0_pmp_7_mask),.io_requestor_1_req_ready(ptw_io_requestor_1_req_ready),.io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),.io_requestor_1_req_bits_valid(ptw_io_requestor_1_req_bits_valid),.io_requestor_1_req_bits_bits_addr(ptw_io_requestor_1_req_bits_bits_addr),.io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),.io_requestor_1_resp_bits_ae(ptw_io_requestor_1_resp_bits_ae),.io_requestor_1_resp_bits_pte_ppn(ptw_io_requestor_1_resp_bits_pte_ppn),.io_requestor_1_resp_bits_pte_d(ptw_io_requestor_1_resp_bits_pte_d),.io_requestor_1_resp_bits_pte_a(ptw_io_requestor_1_resp_bits_pte_a),.io_requestor_1_resp_bits_pte_g(ptw_io_requestor_1_resp_bits_pte_g),.io_requestor_1_resp_bits_pte_u(ptw_io_requestor_1_resp_bits_pte_u),.io_requestor_1_resp_bits_pte_x(ptw_io_requestor_1_resp_bits_pte_x),.io_requestor_1_resp_bits_pte_w(ptw_io_requestor_1_resp_bits_pte_w),.io_requestor_1_resp_bits_pte_r(ptw_io_requestor_1_resp_bits_pte_r),.io_requestor_1_resp_bits_pte_v(ptw_io_requestor_1_resp_bits_pte_v),.io_requestor_1_resp_bits_level(ptw_io_requestor_1_resp_bits_level),.io_requestor_1_resp_bits_homogeneous(ptw_io_requestor_1_resp_bits_homogeneous),.io_requestor_1_ptbr_mode(ptw_io_requestor_1_ptbr_mode),.io_requestor_1_status_debug(ptw_io_requestor_1_status_debug),.io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),.io_requestor_1_pmp_0_cfg_l(ptw_io_requestor_1_pmp_0_cfg_l),.io_requestor_1_pmp_0_cfg_a(ptw_io_requestor_1_pmp_0_cfg_a),.io_requestor_1_pmp_0_cfg_x(ptw_io_requestor_1_pmp_0_cfg_x),.io_requestor_1_pmp_0_cfg_w(ptw_io_requestor_1_pmp_0_cfg_w),.io_requestor_1_pmp_0_cfg_r(ptw_io_requestor_1_pmp_0_cfg_r),.io_requestor_1_pmp_0_addr(ptw_io_requestor_1_pmp_0_addr),.io_requestor_1_pmp_0_mask(ptw_io_requestor_1_pmp_0_mask),.io_requestor_1_pmp_1_cfg_l(ptw_io_requestor_1_pmp_1_cfg_l),.io_requestor_1_pmp_1_cfg_a(ptw_io_requestor_1_pmp_1_cfg_a),.io_requestor_1_pmp_1_cfg_x(ptw_io_requestor_1_pmp_1_cfg_x),.io_requestor_1_pmp_1_cfg_w(ptw_io_requestor_1_pmp_1_cfg_w),.io_requestor_1_pmp_1_cfg_r(ptw_io_requestor_1_pmp_1_cfg_r),.io_requestor_1_pmp_1_addr(ptw_io_requestor_1_pmp_1_addr),.io_requestor_1_pmp_1_mask(ptw_io_requestor_1_pmp_1_mask),.io_requestor_1_pmp_2_cfg_l(ptw_io_requestor_1_pmp_2_cfg_l),.io_requestor_1_pmp_2_cfg_a(ptw_io_requestor_1_pmp_2_cfg_a),.io_requestor_1_pmp_2_cfg_x(ptw_io_requestor_1_pmp_2_cfg_x),.io_requestor_1_pmp_2_cfg_w(ptw_io_requestor_1_pmp_2_cfg_w),.io_requestor_1_pmp_2_cfg_r(ptw_io_requestor_1_pmp_2_cfg_r),.io_requestor_1_pmp_2_addr(ptw_io_requestor_1_pmp_2_addr),.io_requestor_1_pmp_2_mask(ptw_io_requestor_1_pmp_2_mask),.io_requestor_1_pmp_3_cfg_l(ptw_io_requestor_1_pmp_3_cfg_l),.io_requestor_1_pmp_3_cfg_a(ptw_io_requestor_1_pmp_3_cfg_a),.io_requestor_1_pmp_3_cfg_x(ptw_io_requestor_1_pmp_3_cfg_x),.io_requestor_1_pmp_3_cfg_w(ptw_io_requestor_1_pmp_3_cfg_w),.io_requestor_1_pmp_3_cfg_r(ptw_io_requestor_1_pmp_3_cfg_r),.io_requestor_1_pmp_3_addr(ptw_io_requestor_1_pmp_3_addr),.io_requestor_1_pmp_3_mask(ptw_io_requestor_1_pmp_3_mask),.io_requestor_1_pmp_4_cfg_l(ptw_io_requestor_1_pmp_4_cfg_l),.io_requestor_1_pmp_4_cfg_a(ptw_io_requestor_1_pmp_4_cfg_a),.io_requestor_1_pmp_4_cfg_x(ptw_io_requestor_1_pmp_4_cfg_x),.io_requestor_1_pmp_4_cfg_w(ptw_io_requestor_1_pmp_4_cfg_w),.io_requestor_1_pmp_4_cfg_r(ptw_io_requestor_1_pmp_4_cfg_r),.io_requestor_1_pmp_4_addr(ptw_io_requestor_1_pmp_4_addr),.io_requestor_1_pmp_4_mask(ptw_io_requestor_1_pmp_4_mask),.io_requestor_1_pmp_5_cfg_l(ptw_io_requestor_1_pmp_5_cfg_l),.io_requestor_1_pmp_5_cfg_a(ptw_io_requestor_1_pmp_5_cfg_a),.io_requestor_1_pmp_5_cfg_x(ptw_io_requestor_1_pmp_5_cfg_x),.io_requestor_1_pmp_5_cfg_w(ptw_io_requestor_1_pmp_5_cfg_w),.io_requestor_1_pmp_5_cfg_r(ptw_io_requestor_1_pmp_5_cfg_r),.io_requestor_1_pmp_5_addr(ptw_io_requestor_1_pmp_5_addr),.io_requestor_1_pmp_5_mask(ptw_io_requestor_1_pmp_5_mask),.io_requestor_1_pmp_6_cfg_l(ptw_io_requestor_1_pmp_6_cfg_l),.io_requestor_1_pmp_6_cfg_a(ptw_io_requestor_1_pmp_6_cfg_a),.io_requestor_1_pmp_6_cfg_x(ptw_io_requestor_1_pmp_6_cfg_x),.io_requestor_1_pmp_6_cfg_w(ptw_io_requestor_1_pmp_6_cfg_w),.io_requestor_1_pmp_6_cfg_r(ptw_io_requestor_1_pmp_6_cfg_r),.io_requestor_1_pmp_6_addr(ptw_io_requestor_1_pmp_6_addr),.io_requestor_1_pmp_6_mask(ptw_io_requestor_1_pmp_6_mask),.io_requestor_1_pmp_7_cfg_l(ptw_io_requestor_1_pmp_7_cfg_l),.io_requestor_1_pmp_7_cfg_a(ptw_io_requestor_1_pmp_7_cfg_a),.io_requestor_1_pmp_7_cfg_x(ptw_io_requestor_1_pmp_7_cfg_x),.io_requestor_1_pmp_7_cfg_w(ptw_io_requestor_1_pmp_7_cfg_w),.io_requestor_1_pmp_7_cfg_r(ptw_io_requestor_1_pmp_7_cfg_r),.io_requestor_1_pmp_7_addr(ptw_io_requestor_1_pmp_7_addr),.io_requestor_1_pmp_7_mask(ptw_io_requestor_1_pmp_7_mask),.io_requestor_1_customCSRs_csrs_0_value(ptw_io_requestor_1_customCSRs_csrs_0_value),.io_mem_req_ready(ptw_io_mem_req_ready),.io_mem_req_valid(ptw_io_mem_req_valid),.io_mem_req_bits_addr(ptw_io_mem_req_bits_addr),.io_mem_s1_kill(ptw_io_mem_s1_kill),.io_mem_s2_nack(ptw_io_mem_s2_nack),.io_mem_resp_valid(ptw_io_mem_resp_valid),.io_mem_resp_bits_data(ptw_io_mem_resp_bits_data),.io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),.io_dpath_ptbr_mode(ptw_io_dpath_ptbr_mode),.io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),.io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),.io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),.io_dpath_status_debug(ptw_io_dpath_status_debug),.io_dpath_status_dprv(ptw_io_dpath_status_dprv),.io_dpath_status_prv(ptw_io_dpath_status_prv),.io_dpath_status_mxr(ptw_io_dpath_status_mxr),.io_dpath_status_sum(ptw_io_dpath_status_sum),.io_dpath_pmp_0_cfg_l(ptw_io_dpath_pmp_0_cfg_l),.io_dpath_pmp_0_cfg_a(ptw_io_dpath_pmp_0_cfg_a),.io_dpath_pmp_0_cfg_x(ptw_io_dpath_pmp_0_cfg_x),.io_dpath_pmp_0_cfg_w(ptw_io_dpath_pmp_0_cfg_w),.io_dpath_pmp_0_cfg_r(ptw_io_dpath_pmp_0_cfg_r),.io_dpath_pmp_0_addr(ptw_io_dpath_pmp_0_addr),.io_dpath_pmp_0_mask(ptw_io_dpath_pmp_0_mask),.io_dpath_pmp_1_cfg_l(ptw_io_dpath_pmp_1_cfg_l),.io_dpath_pmp_1_cfg_a(ptw_io_dpath_pmp_1_cfg_a),.io_dpath_pmp_1_cfg_x(ptw_io_dpath_pmp_1_cfg_x),.io_dpath_pmp_1_cfg_w(ptw_io_dpath_pmp_1_cfg_w),.io_dpath_pmp_1_cfg_r(ptw_io_dpath_pmp_1_cfg_r),.io_dpath_pmp_1_addr(ptw_io_dpath_pmp_1_addr),.io_dpath_pmp_1_mask(ptw_io_dpath_pmp_1_mask),.io_dpath_pmp_2_cfg_l(ptw_io_dpath_pmp_2_cfg_l),.io_dpath_pmp_2_cfg_a(ptw_io_dpath_pmp_2_cfg_a),.io_dpath_pmp_2_cfg_x(ptw_io_dpath_pmp_2_cfg_x),.io_dpath_pmp_2_cfg_w(ptw_io_dpath_pmp_2_cfg_w),.io_dpath_pmp_2_cfg_r(ptw_io_dpath_pmp_2_cfg_r),.io_dpath_pmp_2_addr(ptw_io_dpath_pmp_2_addr),.io_dpath_pmp_2_mask(ptw_io_dpath_pmp_2_mask),.io_dpath_pmp_3_cfg_l(ptw_io_dpath_pmp_3_cfg_l),.io_dpath_pmp_3_cfg_a(ptw_io_dpath_pmp_3_cfg_a),.io_dpath_pmp_3_cfg_x(ptw_io_dpath_pmp_3_cfg_x),.io_dpath_pmp_3_cfg_w(ptw_io_dpath_pmp_3_cfg_w),.io_dpath_pmp_3_cfg_r(ptw_io_dpath_pmp_3_cfg_r),.io_dpath_pmp_3_addr(ptw_io_dpath_pmp_3_addr),.io_dpath_pmp_3_mask(ptw_io_dpath_pmp_3_mask),.io_dpath_pmp_4_cfg_l(ptw_io_dpath_pmp_4_cfg_l),.io_dpath_pmp_4_cfg_a(ptw_io_dpath_pmp_4_cfg_a),.io_dpath_pmp_4_cfg_x(ptw_io_dpath_pmp_4_cfg_x),.io_dpath_pmp_4_cfg_w(ptw_io_dpath_pmp_4_cfg_w),.io_dpath_pmp_4_cfg_r(ptw_io_dpath_pmp_4_cfg_r),.io_dpath_pmp_4_addr(ptw_io_dpath_pmp_4_addr),.io_dpath_pmp_4_mask(ptw_io_dpath_pmp_4_mask),.io_dpath_pmp_5_cfg_l(ptw_io_dpath_pmp_5_cfg_l),.io_dpath_pmp_5_cfg_a(ptw_io_dpath_pmp_5_cfg_a),.io_dpath_pmp_5_cfg_x(ptw_io_dpath_pmp_5_cfg_x),.io_dpath_pmp_5_cfg_w(ptw_io_dpath_pmp_5_cfg_w),.io_dpath_pmp_5_cfg_r(ptw_io_dpath_pmp_5_cfg_r),.io_dpath_pmp_5_addr(ptw_io_dpath_pmp_5_addr),.io_dpath_pmp_5_mask(ptw_io_dpath_pmp_5_mask),.io_dpath_pmp_6_cfg_l(ptw_io_dpath_pmp_6_cfg_l),.io_dpath_pmp_6_cfg_a(ptw_io_dpath_pmp_6_cfg_a),.io_dpath_pmp_6_cfg_x(ptw_io_dpath_pmp_6_cfg_x),.io_dpath_pmp_6_cfg_w(ptw_io_dpath_pmp_6_cfg_w),.io_dpath_pmp_6_cfg_r(ptw_io_dpath_pmp_6_cfg_r),.io_dpath_pmp_6_addr(ptw_io_dpath_pmp_6_addr),.io_dpath_pmp_6_mask(ptw_io_dpath_pmp_6_mask),.io_dpath_pmp_7_cfg_l(ptw_io_dpath_pmp_7_cfg_l),.io_dpath_pmp_7_cfg_a(ptw_io_dpath_pmp_7_cfg_a),.io_dpath_pmp_7_cfg_x(ptw_io_dpath_pmp_7_cfg_x),.io_dpath_pmp_7_cfg_w(ptw_io_dpath_pmp_7_cfg_w),.io_dpath_pmp_7_cfg_r(ptw_io_dpath_pmp_7_cfg_r),.io_dpath_pmp_7_addr(ptw_io_dpath_pmp_7_addr),.io_dpath_pmp_7_mask(ptw_io_dpath_pmp_7_mask),.io_dpath_perf_l2hit(ptw_io_dpath_perf_l2hit),.io_dpath_perf_pte_miss(ptw_io_dpath_perf_pte_miss),.io_dpath_perf_pte_hit(ptw_io_dpath_perf_pte_hit),.io_dpath_customCSRs_csrs_0_value(ptw_io_dpath_customCSRs_csrs_0_value),.io_covSum(ptw_io_covSum),.metaAssert(ptw_metaAssert),.metaReset(ptw_metaReset)); 
  Rocket core(.clock(core_clock),.reset(core_reset),.io_hartid(core_io_hartid),.io_interrupts_debug(core_io_interrupts_debug),.io_interrupts_mtip(core_io_interrupts_mtip),.io_interrupts_msip(core_io_interrupts_msip),.io_interrupts_meip(core_io_interrupts_meip),.io_interrupts_seip(core_io_interrupts_seip),.io_imem_might_request(core_io_imem_might_request),.io_imem_req_valid(core_io_imem_req_valid),.io_imem_req_bits_pc(core_io_imem_req_bits_pc),.io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),.io_imem_sfence_valid(core_io_imem_sfence_valid),.io_imem_sfence_bits_rs1(core_io_imem_sfence_bits_rs1),.io_imem_sfence_bits_rs2(core_io_imem_sfence_bits_rs2),.io_imem_sfence_bits_addr(core_io_imem_sfence_bits_addr),.io_imem_resp_ready(core_io_imem_resp_ready),.io_imem_resp_valid(core_io_imem_resp_valid),.io_imem_resp_bits_btb_taken(core_io_imem_resp_bits_btb_taken),.io_imem_resp_bits_btb_bridx(core_io_imem_resp_bits_btb_bridx),.io_imem_resp_bits_btb_entry(core_io_imem_resp_bits_btb_entry),.io_imem_resp_bits_btb_bht_history(core_io_imem_resp_bits_btb_bht_history),.io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),.io_imem_resp_bits_data(core_io_imem_resp_bits_data),.io_imem_resp_bits_xcpt_pf_inst(core_io_imem_resp_bits_xcpt_pf_inst),.io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),.io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),.io_imem_btb_update_valid(core_io_imem_btb_update_valid),.io_imem_btb_update_bits_prediction_entry(core_io_imem_btb_update_bits_prediction_entry),.io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),.io_imem_btb_update_bits_isValid(core_io_imem_btb_update_bits_isValid),.io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),.io_imem_btb_update_bits_cfiType(core_io_imem_btb_update_bits_cfiType),.io_imem_bht_update_valid(core_io_imem_bht_update_valid),.io_imem_bht_update_bits_prediction_history(core_io_imem_bht_update_bits_prediction_history),.io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),.io_imem_bht_update_bits_branch(core_io_imem_bht_update_bits_branch),.io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),.io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),.io_imem_flush_icache(core_io_imem_flush_icache),.io_dmem_req_ready(core_io_dmem_req_ready),.io_dmem_req_valid(core_io_dmem_req_valid),.io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),.io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),.io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),.io_dmem_req_bits_size(core_io_dmem_req_bits_size),.io_dmem_req_bits_signed(core_io_dmem_req_bits_signed),.io_dmem_s1_kill(core_io_dmem_s1_kill),.io_dmem_s1_data_data(core_io_dmem_s1_data_data),.io_dmem_s2_nack(core_io_dmem_s2_nack),.io_dmem_resp_valid(core_io_dmem_resp_valid),.io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),.io_dmem_resp_bits_size(core_io_dmem_resp_bits_size),.io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),.io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),.io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),.io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),.io_dmem_replay_next(core_io_dmem_replay_next),.io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),.io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),.io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),.io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),.io_dmem_s2_xcpt_ae_ld(core_io_dmem_s2_xcpt_ae_ld),.io_dmem_s2_xcpt_ae_st(core_io_dmem_s2_xcpt_ae_st),.io_dmem_ordered(core_io_dmem_ordered),.io_dmem_perf_release(core_io_dmem_perf_release),.io_dmem_perf_grant(core_io_dmem_perf_grant),.io_ptw_ptbr_mode(core_io_ptw_ptbr_mode),.io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),.io_ptw_sfence_valid(core_io_ptw_sfence_valid),.io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),.io_ptw_status_debug(core_io_ptw_status_debug),.io_ptw_status_dprv(core_io_ptw_status_dprv),.io_ptw_status_prv(core_io_ptw_status_prv),.io_ptw_status_mxr(core_io_ptw_status_mxr),.io_ptw_status_sum(core_io_ptw_status_sum),.io_ptw_pmp_0_cfg_l(core_io_ptw_pmp_0_cfg_l),.io_ptw_pmp_0_cfg_a(core_io_ptw_pmp_0_cfg_a),.io_ptw_pmp_0_cfg_x(core_io_ptw_pmp_0_cfg_x),.io_ptw_pmp_0_cfg_w(core_io_ptw_pmp_0_cfg_w),.io_ptw_pmp_0_cfg_r(core_io_ptw_pmp_0_cfg_r),.io_ptw_pmp_0_addr(core_io_ptw_pmp_0_addr),.io_ptw_pmp_0_mask(core_io_ptw_pmp_0_mask),.io_ptw_pmp_1_cfg_l(core_io_ptw_pmp_1_cfg_l),.io_ptw_pmp_1_cfg_a(core_io_ptw_pmp_1_cfg_a),.io_ptw_pmp_1_cfg_x(core_io_ptw_pmp_1_cfg_x),.io_ptw_pmp_1_cfg_w(core_io_ptw_pmp_1_cfg_w),.io_ptw_pmp_1_cfg_r(core_io_ptw_pmp_1_cfg_r),.io_ptw_pmp_1_addr(core_io_ptw_pmp_1_addr),.io_ptw_pmp_1_mask(core_io_ptw_pmp_1_mask),.io_ptw_pmp_2_cfg_l(core_io_ptw_pmp_2_cfg_l),.io_ptw_pmp_2_cfg_a(core_io_ptw_pmp_2_cfg_a),.io_ptw_pmp_2_cfg_x(core_io_ptw_pmp_2_cfg_x),.io_ptw_pmp_2_cfg_w(core_io_ptw_pmp_2_cfg_w),.io_ptw_pmp_2_cfg_r(core_io_ptw_pmp_2_cfg_r),.io_ptw_pmp_2_addr(core_io_ptw_pmp_2_addr),.io_ptw_pmp_2_mask(core_io_ptw_pmp_2_mask),.io_ptw_pmp_3_cfg_l(core_io_ptw_pmp_3_cfg_l),.io_ptw_pmp_3_cfg_a(core_io_ptw_pmp_3_cfg_a),.io_ptw_pmp_3_cfg_x(core_io_ptw_pmp_3_cfg_x),.io_ptw_pmp_3_cfg_w(core_io_ptw_pmp_3_cfg_w),.io_ptw_pmp_3_cfg_r(core_io_ptw_pmp_3_cfg_r),.io_ptw_pmp_3_addr(core_io_ptw_pmp_3_addr),.io_ptw_pmp_3_mask(core_io_ptw_pmp_3_mask),.io_ptw_pmp_4_cfg_l(core_io_ptw_pmp_4_cfg_l),.io_ptw_pmp_4_cfg_a(core_io_ptw_pmp_4_cfg_a),.io_ptw_pmp_4_cfg_x(core_io_ptw_pmp_4_cfg_x),.io_ptw_pmp_4_cfg_w(core_io_ptw_pmp_4_cfg_w),.io_ptw_pmp_4_cfg_r(core_io_ptw_pmp_4_cfg_r),.io_ptw_pmp_4_addr(core_io_ptw_pmp_4_addr),.io_ptw_pmp_4_mask(core_io_ptw_pmp_4_mask),.io_ptw_pmp_5_cfg_l(core_io_ptw_pmp_5_cfg_l),.io_ptw_pmp_5_cfg_a(core_io_ptw_pmp_5_cfg_a),.io_ptw_pmp_5_cfg_x(core_io_ptw_pmp_5_cfg_x),.io_ptw_pmp_5_cfg_w(core_io_ptw_pmp_5_cfg_w),.io_ptw_pmp_5_cfg_r(core_io_ptw_pmp_5_cfg_r),.io_ptw_pmp_5_addr(core_io_ptw_pmp_5_addr),.io_ptw_pmp_5_mask(core_io_ptw_pmp_5_mask),.io_ptw_pmp_6_cfg_l(core_io_ptw_pmp_6_cfg_l),.io_ptw_pmp_6_cfg_a(core_io_ptw_pmp_6_cfg_a),.io_ptw_pmp_6_cfg_x(core_io_ptw_pmp_6_cfg_x),.io_ptw_pmp_6_cfg_w(core_io_ptw_pmp_6_cfg_w),.io_ptw_pmp_6_cfg_r(core_io_ptw_pmp_6_cfg_r),.io_ptw_pmp_6_addr(core_io_ptw_pmp_6_addr),.io_ptw_pmp_6_mask(core_io_ptw_pmp_6_mask),.io_ptw_pmp_7_cfg_l(core_io_ptw_pmp_7_cfg_l),.io_ptw_pmp_7_cfg_a(core_io_ptw_pmp_7_cfg_a),.io_ptw_pmp_7_cfg_x(core_io_ptw_pmp_7_cfg_x),.io_ptw_pmp_7_cfg_w(core_io_ptw_pmp_7_cfg_w),.io_ptw_pmp_7_cfg_r(core_io_ptw_pmp_7_cfg_r),.io_ptw_pmp_7_addr(core_io_ptw_pmp_7_addr),.io_ptw_pmp_7_mask(core_io_ptw_pmp_7_mask),.io_ptw_customCSRs_csrs_0_value(core_io_ptw_customCSRs_csrs_0_value),.io_fpu_inst(core_io_fpu_inst),.io_fpu_fromint_data(core_io_fpu_fromint_data),.io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),.io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),.io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),.io_fpu_store_data(core_io_fpu_store_data),.io_fpu_toint_data(core_io_fpu_toint_data),.io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),.io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),.io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),.io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),.io_fpu_valid(core_io_fpu_valid),.io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),.io_fpu_nack_mem(core_io_fpu_nack_mem),.io_fpu_illegal_rm(core_io_fpu_illegal_rm),.io_fpu_killx(core_io_fpu_killx),.io_fpu_killm(core_io_fpu_killm),.io_fpu_dec_wen(core_io_fpu_dec_wen),.io_fpu_dec_ren1(core_io_fpu_dec_ren1),.io_fpu_dec_ren2(core_io_fpu_dec_ren2),.io_fpu_dec_ren3(core_io_fpu_dec_ren3),.io_fpu_sboard_set(core_io_fpu_sboard_set),.io_fpu_sboard_clr(core_io_fpu_sboard_clr),.io_fpu_sboard_clra(core_io_fpu_sboard_clra),.io_trace_0_valid(core_io_trace_0_valid),.io_trace_0_iaddr(core_io_trace_0_iaddr),.io_trace_0_insn(core_io_trace_0_insn),.io_trace_0_priv(core_io_trace_0_priv),.io_trace_0_exception(core_io_trace_0_exception),.io_trace_0_interrupt(core_io_trace_0_interrupt),.io_trace_0_cause(core_io_trace_0_cause),.io_trace_0_tval(core_io_trace_0_tval),.io_wfi(core_io_wfi),.io_covSum(core_io_covSum),.metaAssert(core_metaAssert),.metaReset(core_metaReset),.PlusArgTimeout_halt(core_PlusArgTimeout_halt),.csr_halt(core_csr_halt),.ibuf_halt(core_ibuf_halt),.div_halt(core_div_halt)); 
  assign auto_broadcast_out_0_valid=broadcast_3_auto_out_0_valid; 
  assign auto_broadcast_out_0_iaddr=broadcast_3_auto_out_0_iaddr; 
  assign auto_broadcast_out_0_insn=broadcast_3_auto_out_0_insn; 
  assign auto_broadcast_out_0_priv=broadcast_3_auto_out_0_priv; 
  assign auto_broadcast_out_0_exception=broadcast_3_auto_out_0_exception; 
  assign auto_broadcast_out_0_interrupt=broadcast_3_auto_out_0_interrupt; 
  assign auto_broadcast_out_0_cause=broadcast_3_auto_out_0_cause; 
  assign auto_broadcast_out_0_tval=broadcast_3_auto_out_0_tval; 
  assign auto_wfi_out_0=bundleOut_0_0_REG; 
  assign auto_cease_out_0=1'h0; 
  assign auto_halt_out_0=1'h0; 
  assign auto_trace_core_source_out_group_0_iretire=1'h0; 
  assign auto_trace_core_source_out_group_0_iaddr=32'h0; 
  assign auto_trace_core_source_out_group_0_itype=4'h0; 
  assign auto_trace_core_source_out_group_0_ilastsize=1'h0; 
  assign auto_trace_core_source_out_priv=4'h0; 
  assign auto_trace_core_source_out_tval=32'h0; 
  assign auto_trace_core_source_out_cause=32'h0; 
  assign auto_tl_master_xing_out_a_valid=tlMasterXbar_auto_out_a_valid; 
  assign auto_tl_master_xing_out_a_bits_opcode=tlMasterXbar_auto_out_a_bits_opcode; 
  assign auto_tl_master_xing_out_a_bits_param=tlMasterXbar_auto_out_a_bits_param; 
  assign auto_tl_master_xing_out_a_bits_size=tlMasterXbar_auto_out_a_bits_size; 
  assign auto_tl_master_xing_out_a_bits_source=tlMasterXbar_auto_out_a_bits_source; 
  assign auto_tl_master_xing_out_a_bits_address=tlMasterXbar_auto_out_a_bits_address; 
  assign auto_tl_master_xing_out_a_bits_mask=tlMasterXbar_auto_out_a_bits_mask; 
  assign auto_tl_master_xing_out_a_bits_data=tlMasterXbar_auto_out_a_bits_data; 
  assign auto_tl_master_xing_out_a_bits_corrupt=1'h0; 
  assign auto_tl_master_xing_out_b_ready=tlMasterXbar_auto_out_b_ready; 
  assign auto_tl_master_xing_out_c_valid=tlMasterXbar_auto_out_c_valid; 
  assign auto_tl_master_xing_out_c_bits_opcode=tlMasterXbar_auto_out_c_bits_opcode; 
  assign auto_tl_master_xing_out_c_bits_param=tlMasterXbar_auto_out_c_bits_param; 
  assign auto_tl_master_xing_out_c_bits_size=tlMasterXbar_auto_out_c_bits_size; 
  assign auto_tl_master_xing_out_c_bits_source=tlMasterXbar_auto_out_c_bits_source; 
  assign auto_tl_master_xing_out_c_bits_address=tlMasterXbar_auto_out_c_bits_address; 
  assign auto_tl_master_xing_out_c_bits_data=tlMasterXbar_auto_out_c_bits_data; 
  assign auto_tl_master_xing_out_c_bits_corrupt=1'h0; 
  assign auto_tl_master_xing_out_d_ready=tlMasterXbar_auto_out_d_ready; 
  assign auto_tl_master_xing_out_e_valid=tlMasterXbar_auto_out_e_valid; 
  assign auto_tl_master_xing_out_e_bits_sink=tlMasterXbar_auto_out_e_bits_sink; 
  assign tlMasterXbar_clock=clock; 
  assign tlMasterXbar_reset=reset; 
  assign tlMasterXbar_auto_in_1_a_valid=frontend_auto_icache_master_out_a_valid; 
  assign tlMasterXbar_auto_in_1_a_bits_address=frontend_auto_icache_master_out_a_bits_address; 
  assign tlMasterXbar_auto_in_0_a_valid=dcache_auto_out_a_valid; 
  assign tlMasterXbar_auto_in_0_a_bits_opcode=dcache_auto_out_a_bits_opcode; 
  assign tlMasterXbar_auto_in_0_a_bits_param=dcache_auto_out_a_bits_param; 
  assign tlMasterXbar_auto_in_0_a_bits_size=dcache_auto_out_a_bits_size; 
  assign tlMasterXbar_auto_in_0_a_bits_source=dcache_auto_out_a_bits_source; 
  assign tlMasterXbar_auto_in_0_a_bits_address=dcache_auto_out_a_bits_address; 
  assign tlMasterXbar_auto_in_0_a_bits_mask=dcache_auto_out_a_bits_mask; 
  assign tlMasterXbar_auto_in_0_a_bits_data=dcache_auto_out_a_bits_data; 
  assign tlMasterXbar_auto_in_0_b_ready=dcache_auto_out_b_ready; 
  assign tlMasterXbar_auto_in_0_c_valid=dcache_auto_out_c_valid; 
  assign tlMasterXbar_auto_in_0_c_bits_opcode=dcache_auto_out_c_bits_opcode; 
  assign tlMasterXbar_auto_in_0_c_bits_param=dcache_auto_out_c_bits_param; 
  assign tlMasterXbar_auto_in_0_c_bits_size=dcache_auto_out_c_bits_size; 
  assign tlMasterXbar_auto_in_0_c_bits_source=dcache_auto_out_c_bits_source; 
  assign tlMasterXbar_auto_in_0_c_bits_address=dcache_auto_out_c_bits_address; 
  assign tlMasterXbar_auto_in_0_c_bits_data=dcache_auto_out_c_bits_data; 
  assign tlMasterXbar_auto_in_0_d_ready=dcache_auto_out_d_ready; 
  assign tlMasterXbar_auto_in_0_e_valid=dcache_auto_out_e_valid; 
  assign tlMasterXbar_auto_in_0_e_bits_sink=dcache_auto_out_e_bits_sink; 
  assign tlMasterXbar_auto_out_a_ready=auto_tl_master_xing_out_a_ready; 
  assign tlMasterXbar_auto_out_b_valid=auto_tl_master_xing_out_b_valid; 
  assign tlMasterXbar_auto_out_b_bits_opcode=auto_tl_master_xing_out_b_bits_opcode; 
  assign tlMasterXbar_auto_out_b_bits_param=auto_tl_master_xing_out_b_bits_param; 
  assign tlMasterXbar_auto_out_b_bits_size=auto_tl_master_xing_out_b_bits_size; 
  assign tlMasterXbar_auto_out_b_bits_source=auto_tl_master_xing_out_b_bits_source; 
  assign tlMasterXbar_auto_out_b_bits_address=auto_tl_master_xing_out_b_bits_address; 
  assign tlMasterXbar_auto_out_b_bits_mask=auto_tl_master_xing_out_b_bits_mask; 
  assign tlMasterXbar_auto_out_b_bits_corrupt=auto_tl_master_xing_out_b_bits_corrupt; 
  assign tlMasterXbar_auto_out_c_ready=auto_tl_master_xing_out_c_ready; 
  assign tlMasterXbar_auto_out_d_valid=auto_tl_master_xing_out_d_valid; 
  assign tlMasterXbar_auto_out_d_bits_opcode=auto_tl_master_xing_out_d_bits_opcode; 
  assign tlMasterXbar_auto_out_d_bits_param=auto_tl_master_xing_out_d_bits_param; 
  assign tlMasterXbar_auto_out_d_bits_size=auto_tl_master_xing_out_d_bits_size; 
  assign tlMasterXbar_auto_out_d_bits_source=auto_tl_master_xing_out_d_bits_source; 
  assign tlMasterXbar_auto_out_d_bits_sink=auto_tl_master_xing_out_d_bits_sink; 
  assign tlMasterXbar_auto_out_d_bits_denied=auto_tl_master_xing_out_d_bits_denied; 
  assign tlMasterXbar_auto_out_d_bits_data=auto_tl_master_xing_out_d_bits_data; 
  assign tlMasterXbar_auto_out_d_bits_corrupt=auto_tl_master_xing_out_d_bits_corrupt; 
  assign tlMasterXbar_auto_out_e_ready=auto_tl_master_xing_out_e_ready; 
  assign intXbar_auto_int_in_3_0=auto_int_in_xing_in_2_sync_0; 
  assign intXbar_auto_int_in_2_0=auto_int_in_xing_in_1_sync_0; 
  assign intXbar_auto_int_in_1_0=auto_int_in_xing_in_0_sync_0; 
  assign intXbar_auto_int_in_1_1=auto_int_in_xing_in_0_sync_1; 
  assign intXbar_auto_int_in_0_0=auto_intsink_in_sync_0; 
  assign broadcast_auto_in=auto_hartid_in; 
  assign broadcast_1_auto_in=auto_reset_vector_in; 
  assign broadcast_3_auto_in_0_valid=core_io_trace_0_valid; 
  assign broadcast_3_auto_in_0_iaddr=core_io_trace_0_iaddr; 
  assign broadcast_3_auto_in_0_insn=core_io_trace_0_insn; 
  assign broadcast_3_auto_in_0_priv=core_io_trace_0_priv; 
  assign broadcast_3_auto_in_0_exception=core_io_trace_0_exception; 
  assign broadcast_3_auto_in_0_interrupt=core_io_trace_0_interrupt; 
  assign broadcast_3_auto_in_0_cause=core_io_trace_0_cause; 
  assign broadcast_3_auto_in_0_tval=core_io_trace_0_tval; 
  assign dcache_gated_clock=clock; 
  assign dcache_reset=reset; 
  assign dcache_auto_out_a_ready=tlMasterXbar_auto_in_0_a_ready; 
  assign dcache_auto_out_b_valid=tlMasterXbar_auto_in_0_b_valid; 
  assign dcache_auto_out_b_bits_param=tlMasterXbar_auto_in_0_b_bits_param; 
  assign dcache_auto_out_b_bits_size=tlMasterXbar_auto_in_0_b_bits_size; 
  assign dcache_auto_out_b_bits_source=tlMasterXbar_auto_in_0_b_bits_source; 
  assign dcache_auto_out_b_bits_address=tlMasterXbar_auto_in_0_b_bits_address; 
  assign dcache_auto_out_c_ready=tlMasterXbar_auto_in_0_c_ready; 
  assign dcache_auto_out_d_valid=tlMasterXbar_auto_in_0_d_valid; 
  assign dcache_auto_out_d_bits_opcode=tlMasterXbar_auto_in_0_d_bits_opcode; 
  assign dcache_auto_out_d_bits_param=tlMasterXbar_auto_in_0_d_bits_param; 
  assign dcache_auto_out_d_bits_size=tlMasterXbar_auto_in_0_d_bits_size; 
  assign dcache_auto_out_d_bits_source=tlMasterXbar_auto_in_0_d_bits_source; 
  assign dcache_auto_out_d_bits_sink=tlMasterXbar_auto_in_0_d_bits_sink; 
  assign dcache_auto_out_d_bits_denied=tlMasterXbar_auto_in_0_d_bits_denied; 
  assign dcache_auto_out_d_bits_data=tlMasterXbar_auto_in_0_d_bits_data; 
  assign dcache_auto_out_e_ready=tlMasterXbar_auto_in_0_e_ready; 
  assign dcache_io_cpu_req_valid=dcacheArb_io_mem_req_valid; 
  assign dcache_io_cpu_req_bits_addr=dcacheArb_io_mem_req_bits_addr; 
  assign dcache_io_cpu_req_bits_tag=dcacheArb_io_mem_req_bits_tag; 
  assign dcache_io_cpu_req_bits_cmd=dcacheArb_io_mem_req_bits_cmd; 
  assign dcache_io_cpu_req_bits_size=dcacheArb_io_mem_req_bits_size; 
  assign dcache_io_cpu_req_bits_signed=dcacheArb_io_mem_req_bits_signed; 
  assign dcache_io_cpu_req_bits_phys=dcacheArb_io_mem_req_bits_phys; 
  assign dcache_io_cpu_s1_kill=dcacheArb_io_mem_s1_kill; 
  assign dcache_io_cpu_s1_data_data=dcacheArb_io_mem_s1_data_data; 
  assign dcache_io_ptw_req_ready=ptw_io_requestor_0_req_ready; 
  assign dcache_io_ptw_resp_valid=ptw_io_requestor_0_resp_valid; 
  assign dcache_io_ptw_resp_bits_ae=ptw_io_requestor_0_resp_bits_ae; 
  assign dcache_io_ptw_resp_bits_pte_ppn=ptw_io_requestor_0_resp_bits_pte_ppn; 
  assign dcache_io_ptw_resp_bits_pte_d=ptw_io_requestor_0_resp_bits_pte_d; 
  assign dcache_io_ptw_resp_bits_pte_a=ptw_io_requestor_0_resp_bits_pte_a; 
  assign dcache_io_ptw_resp_bits_pte_g=ptw_io_requestor_0_resp_bits_pte_g; 
  assign dcache_io_ptw_resp_bits_pte_u=ptw_io_requestor_0_resp_bits_pte_u; 
  assign dcache_io_ptw_resp_bits_pte_x=ptw_io_requestor_0_resp_bits_pte_x; 
  assign dcache_io_ptw_resp_bits_pte_w=ptw_io_requestor_0_resp_bits_pte_w; 
  assign dcache_io_ptw_resp_bits_pte_r=ptw_io_requestor_0_resp_bits_pte_r; 
  assign dcache_io_ptw_resp_bits_pte_v=ptw_io_requestor_0_resp_bits_pte_v; 
  assign dcache_io_ptw_resp_bits_level=ptw_io_requestor_0_resp_bits_level; 
  assign dcache_io_ptw_resp_bits_homogeneous=ptw_io_requestor_0_resp_bits_homogeneous; 
  assign dcache_io_ptw_ptbr_mode=ptw_io_requestor_0_ptbr_mode; 
  assign dcache_io_ptw_status_debug=ptw_io_requestor_0_status_debug; 
  assign dcache_io_ptw_status_dprv=ptw_io_requestor_0_status_dprv; 
  assign dcache_io_ptw_status_mxr=ptw_io_requestor_0_status_mxr; 
  assign dcache_io_ptw_status_sum=ptw_io_requestor_0_status_sum; 
  assign dcache_io_ptw_pmp_0_cfg_l=ptw_io_requestor_0_pmp_0_cfg_l; 
  assign dcache_io_ptw_pmp_0_cfg_a=ptw_io_requestor_0_pmp_0_cfg_a; 
  assign dcache_io_ptw_pmp_0_cfg_x=ptw_io_requestor_0_pmp_0_cfg_x; 
  assign dcache_io_ptw_pmp_0_cfg_w=ptw_io_requestor_0_pmp_0_cfg_w; 
  assign dcache_io_ptw_pmp_0_cfg_r=ptw_io_requestor_0_pmp_0_cfg_r; 
  assign dcache_io_ptw_pmp_0_addr=ptw_io_requestor_0_pmp_0_addr; 
  assign dcache_io_ptw_pmp_0_mask=ptw_io_requestor_0_pmp_0_mask; 
  assign dcache_io_ptw_pmp_1_cfg_l=ptw_io_requestor_0_pmp_1_cfg_l; 
  assign dcache_io_ptw_pmp_1_cfg_a=ptw_io_requestor_0_pmp_1_cfg_a; 
  assign dcache_io_ptw_pmp_1_cfg_x=ptw_io_requestor_0_pmp_1_cfg_x; 
  assign dcache_io_ptw_pmp_1_cfg_w=ptw_io_requestor_0_pmp_1_cfg_w; 
  assign dcache_io_ptw_pmp_1_cfg_r=ptw_io_requestor_0_pmp_1_cfg_r; 
  assign dcache_io_ptw_pmp_1_addr=ptw_io_requestor_0_pmp_1_addr; 
  assign dcache_io_ptw_pmp_1_mask=ptw_io_requestor_0_pmp_1_mask; 
  assign dcache_io_ptw_pmp_2_cfg_l=ptw_io_requestor_0_pmp_2_cfg_l; 
  assign dcache_io_ptw_pmp_2_cfg_a=ptw_io_requestor_0_pmp_2_cfg_a; 
  assign dcache_io_ptw_pmp_2_cfg_x=ptw_io_requestor_0_pmp_2_cfg_x; 
  assign dcache_io_ptw_pmp_2_cfg_w=ptw_io_requestor_0_pmp_2_cfg_w; 
  assign dcache_io_ptw_pmp_2_cfg_r=ptw_io_requestor_0_pmp_2_cfg_r; 
  assign dcache_io_ptw_pmp_2_addr=ptw_io_requestor_0_pmp_2_addr; 
  assign dcache_io_ptw_pmp_2_mask=ptw_io_requestor_0_pmp_2_mask; 
  assign dcache_io_ptw_pmp_3_cfg_l=ptw_io_requestor_0_pmp_3_cfg_l; 
  assign dcache_io_ptw_pmp_3_cfg_a=ptw_io_requestor_0_pmp_3_cfg_a; 
  assign dcache_io_ptw_pmp_3_cfg_x=ptw_io_requestor_0_pmp_3_cfg_x; 
  assign dcache_io_ptw_pmp_3_cfg_w=ptw_io_requestor_0_pmp_3_cfg_w; 
  assign dcache_io_ptw_pmp_3_cfg_r=ptw_io_requestor_0_pmp_3_cfg_r; 
  assign dcache_io_ptw_pmp_3_addr=ptw_io_requestor_0_pmp_3_addr; 
  assign dcache_io_ptw_pmp_3_mask=ptw_io_requestor_0_pmp_3_mask; 
  assign dcache_io_ptw_pmp_4_cfg_l=ptw_io_requestor_0_pmp_4_cfg_l; 
  assign dcache_io_ptw_pmp_4_cfg_a=ptw_io_requestor_0_pmp_4_cfg_a; 
  assign dcache_io_ptw_pmp_4_cfg_x=ptw_io_requestor_0_pmp_4_cfg_x; 
  assign dcache_io_ptw_pmp_4_cfg_w=ptw_io_requestor_0_pmp_4_cfg_w; 
  assign dcache_io_ptw_pmp_4_cfg_r=ptw_io_requestor_0_pmp_4_cfg_r; 
  assign dcache_io_ptw_pmp_4_addr=ptw_io_requestor_0_pmp_4_addr; 
  assign dcache_io_ptw_pmp_4_mask=ptw_io_requestor_0_pmp_4_mask; 
  assign dcache_io_ptw_pmp_5_cfg_l=ptw_io_requestor_0_pmp_5_cfg_l; 
  assign dcache_io_ptw_pmp_5_cfg_a=ptw_io_requestor_0_pmp_5_cfg_a; 
  assign dcache_io_ptw_pmp_5_cfg_x=ptw_io_requestor_0_pmp_5_cfg_x; 
  assign dcache_io_ptw_pmp_5_cfg_w=ptw_io_requestor_0_pmp_5_cfg_w; 
  assign dcache_io_ptw_pmp_5_cfg_r=ptw_io_requestor_0_pmp_5_cfg_r; 
  assign dcache_io_ptw_pmp_5_addr=ptw_io_requestor_0_pmp_5_addr; 
  assign dcache_io_ptw_pmp_5_mask=ptw_io_requestor_0_pmp_5_mask; 
  assign dcache_io_ptw_pmp_6_cfg_l=ptw_io_requestor_0_pmp_6_cfg_l; 
  assign dcache_io_ptw_pmp_6_cfg_a=ptw_io_requestor_0_pmp_6_cfg_a; 
  assign dcache_io_ptw_pmp_6_cfg_x=ptw_io_requestor_0_pmp_6_cfg_x; 
  assign dcache_io_ptw_pmp_6_cfg_w=ptw_io_requestor_0_pmp_6_cfg_w; 
  assign dcache_io_ptw_pmp_6_cfg_r=ptw_io_requestor_0_pmp_6_cfg_r; 
  assign dcache_io_ptw_pmp_6_addr=ptw_io_requestor_0_pmp_6_addr; 
  assign dcache_io_ptw_pmp_6_mask=ptw_io_requestor_0_pmp_6_mask; 
  assign dcache_io_ptw_pmp_7_cfg_l=ptw_io_requestor_0_pmp_7_cfg_l; 
  assign dcache_io_ptw_pmp_7_cfg_a=ptw_io_requestor_0_pmp_7_cfg_a; 
  assign dcache_io_ptw_pmp_7_cfg_x=ptw_io_requestor_0_pmp_7_cfg_x; 
  assign dcache_io_ptw_pmp_7_cfg_w=ptw_io_requestor_0_pmp_7_cfg_w; 
  assign dcache_io_ptw_pmp_7_cfg_r=ptw_io_requestor_0_pmp_7_cfg_r; 
  assign dcache_io_ptw_pmp_7_addr=ptw_io_requestor_0_pmp_7_addr; 
  assign dcache_io_ptw_pmp_7_mask=ptw_io_requestor_0_pmp_7_mask; 
  assign frontend_gated_clock=clock; 
  assign frontend_reset=reset; 
  assign frontend_auto_icache_master_out_a_ready=tlMasterXbar_auto_in_1_a_ready; 
  assign frontend_auto_icache_master_out_d_valid=tlMasterXbar_auto_in_1_d_valid; 
  assign frontend_auto_icache_master_out_d_bits_opcode=tlMasterXbar_auto_in_1_d_bits_opcode; 
  assign frontend_auto_icache_master_out_d_bits_size=tlMasterXbar_auto_in_1_d_bits_size; 
  assign frontend_auto_icache_master_out_d_bits_data=tlMasterXbar_auto_in_1_d_bits_data; 
  assign frontend_auto_icache_master_out_d_bits_corrupt=tlMasterXbar_auto_in_1_d_bits_corrupt; 
  assign frontend_auto_reset_vector_sink_in=broadcast_1_auto_out_1; 
  assign frontend_io_cpu_might_request=core_io_imem_might_request; 
  assign frontend_io_cpu_req_valid=core_io_imem_req_valid; 
  assign frontend_io_cpu_req_bits_pc=core_io_imem_req_bits_pc; 
  assign frontend_io_cpu_req_bits_speculative=core_io_imem_req_bits_speculative; 
  assign frontend_io_cpu_sfence_valid=core_io_imem_sfence_valid; 
  assign frontend_io_cpu_sfence_bits_rs1=core_io_imem_sfence_bits_rs1; 
  assign frontend_io_cpu_sfence_bits_rs2=core_io_imem_sfence_bits_rs2; 
  assign frontend_io_cpu_sfence_bits_addr=core_io_imem_sfence_bits_addr; 
  assign frontend_io_cpu_resp_ready=core_io_imem_resp_ready; 
  assign frontend_io_cpu_btb_update_valid=core_io_imem_btb_update_valid; 
  assign frontend_io_cpu_btb_update_bits_prediction_entry=core_io_imem_btb_update_bits_prediction_entry; 
  assign frontend_io_cpu_btb_update_bits_pc=core_io_imem_btb_update_bits_pc; 
  assign frontend_io_cpu_btb_update_bits_isValid=core_io_imem_btb_update_bits_isValid; 
  assign frontend_io_cpu_btb_update_bits_br_pc=core_io_imem_btb_update_bits_br_pc; 
  assign frontend_io_cpu_btb_update_bits_cfiType=core_io_imem_btb_update_bits_cfiType; 
  assign frontend_io_cpu_bht_update_valid=core_io_imem_bht_update_valid; 
  assign frontend_io_cpu_bht_update_bits_prediction_history=core_io_imem_bht_update_bits_prediction_history; 
  assign frontend_io_cpu_bht_update_bits_pc=core_io_imem_bht_update_bits_pc; 
  assign frontend_io_cpu_bht_update_bits_branch=core_io_imem_bht_update_bits_branch; 
  assign frontend_io_cpu_bht_update_bits_taken=core_io_imem_bht_update_bits_taken; 
  assign frontend_io_cpu_bht_update_bits_mispredict=core_io_imem_bht_update_bits_mispredict; 
  assign frontend_io_cpu_flush_icache=core_io_imem_flush_icache; 
  assign frontend_io_ptw_req_ready=ptw_io_requestor_1_req_ready; 
  assign frontend_io_ptw_resp_valid=ptw_io_requestor_1_resp_valid; 
  assign frontend_io_ptw_resp_bits_ae=ptw_io_requestor_1_resp_bits_ae; 
  assign frontend_io_ptw_resp_bits_pte_ppn=ptw_io_requestor_1_resp_bits_pte_ppn; 
  assign frontend_io_ptw_resp_bits_pte_d=ptw_io_requestor_1_resp_bits_pte_d; 
  assign frontend_io_ptw_resp_bits_pte_a=ptw_io_requestor_1_resp_bits_pte_a; 
  assign frontend_io_ptw_resp_bits_pte_g=ptw_io_requestor_1_resp_bits_pte_g; 
  assign frontend_io_ptw_resp_bits_pte_u=ptw_io_requestor_1_resp_bits_pte_u; 
  assign frontend_io_ptw_resp_bits_pte_x=ptw_io_requestor_1_resp_bits_pte_x; 
  assign frontend_io_ptw_resp_bits_pte_w=ptw_io_requestor_1_resp_bits_pte_w; 
  assign frontend_io_ptw_resp_bits_pte_r=ptw_io_requestor_1_resp_bits_pte_r; 
  assign frontend_io_ptw_resp_bits_pte_v=ptw_io_requestor_1_resp_bits_pte_v; 
  assign frontend_io_ptw_resp_bits_level=ptw_io_requestor_1_resp_bits_level; 
  assign frontend_io_ptw_resp_bits_homogeneous=ptw_io_requestor_1_resp_bits_homogeneous; 
  assign frontend_io_ptw_ptbr_mode=ptw_io_requestor_1_ptbr_mode; 
  assign frontend_io_ptw_status_debug=ptw_io_requestor_1_status_debug; 
  assign frontend_io_ptw_status_prv=ptw_io_requestor_1_status_prv; 
  assign frontend_io_ptw_pmp_0_cfg_l=ptw_io_requestor_1_pmp_0_cfg_l; 
  assign frontend_io_ptw_pmp_0_cfg_a=ptw_io_requestor_1_pmp_0_cfg_a; 
  assign frontend_io_ptw_pmp_0_cfg_x=ptw_io_requestor_1_pmp_0_cfg_x; 
  assign frontend_io_ptw_pmp_0_cfg_w=ptw_io_requestor_1_pmp_0_cfg_w; 
  assign frontend_io_ptw_pmp_0_cfg_r=ptw_io_requestor_1_pmp_0_cfg_r; 
  assign frontend_io_ptw_pmp_0_addr=ptw_io_requestor_1_pmp_0_addr; 
  assign frontend_io_ptw_pmp_0_mask=ptw_io_requestor_1_pmp_0_mask; 
  assign frontend_io_ptw_pmp_1_cfg_l=ptw_io_requestor_1_pmp_1_cfg_l; 
  assign frontend_io_ptw_pmp_1_cfg_a=ptw_io_requestor_1_pmp_1_cfg_a; 
  assign frontend_io_ptw_pmp_1_cfg_x=ptw_io_requestor_1_pmp_1_cfg_x; 
  assign frontend_io_ptw_pmp_1_cfg_w=ptw_io_requestor_1_pmp_1_cfg_w; 
  assign frontend_io_ptw_pmp_1_cfg_r=ptw_io_requestor_1_pmp_1_cfg_r; 
  assign frontend_io_ptw_pmp_1_addr=ptw_io_requestor_1_pmp_1_addr; 
  assign frontend_io_ptw_pmp_1_mask=ptw_io_requestor_1_pmp_1_mask; 
  assign frontend_io_ptw_pmp_2_cfg_l=ptw_io_requestor_1_pmp_2_cfg_l; 
  assign frontend_io_ptw_pmp_2_cfg_a=ptw_io_requestor_1_pmp_2_cfg_a; 
  assign frontend_io_ptw_pmp_2_cfg_x=ptw_io_requestor_1_pmp_2_cfg_x; 
  assign frontend_io_ptw_pmp_2_cfg_w=ptw_io_requestor_1_pmp_2_cfg_w; 
  assign frontend_io_ptw_pmp_2_cfg_r=ptw_io_requestor_1_pmp_2_cfg_r; 
  assign frontend_io_ptw_pmp_2_addr=ptw_io_requestor_1_pmp_2_addr; 
  assign frontend_io_ptw_pmp_2_mask=ptw_io_requestor_1_pmp_2_mask; 
  assign frontend_io_ptw_pmp_3_cfg_l=ptw_io_requestor_1_pmp_3_cfg_l; 
  assign frontend_io_ptw_pmp_3_cfg_a=ptw_io_requestor_1_pmp_3_cfg_a; 
  assign frontend_io_ptw_pmp_3_cfg_x=ptw_io_requestor_1_pmp_3_cfg_x; 
  assign frontend_io_ptw_pmp_3_cfg_w=ptw_io_requestor_1_pmp_3_cfg_w; 
  assign frontend_io_ptw_pmp_3_cfg_r=ptw_io_requestor_1_pmp_3_cfg_r; 
  assign frontend_io_ptw_pmp_3_addr=ptw_io_requestor_1_pmp_3_addr; 
  assign frontend_io_ptw_pmp_3_mask=ptw_io_requestor_1_pmp_3_mask; 
  assign frontend_io_ptw_pmp_4_cfg_l=ptw_io_requestor_1_pmp_4_cfg_l; 
  assign frontend_io_ptw_pmp_4_cfg_a=ptw_io_requestor_1_pmp_4_cfg_a; 
  assign frontend_io_ptw_pmp_4_cfg_x=ptw_io_requestor_1_pmp_4_cfg_x; 
  assign frontend_io_ptw_pmp_4_cfg_w=ptw_io_requestor_1_pmp_4_cfg_w; 
  assign frontend_io_ptw_pmp_4_cfg_r=ptw_io_requestor_1_pmp_4_cfg_r; 
  assign frontend_io_ptw_pmp_4_addr=ptw_io_requestor_1_pmp_4_addr; 
  assign frontend_io_ptw_pmp_4_mask=ptw_io_requestor_1_pmp_4_mask; 
  assign frontend_io_ptw_pmp_5_cfg_l=ptw_io_requestor_1_pmp_5_cfg_l; 
  assign frontend_io_ptw_pmp_5_cfg_a=ptw_io_requestor_1_pmp_5_cfg_a; 
  assign frontend_io_ptw_pmp_5_cfg_x=ptw_io_requestor_1_pmp_5_cfg_x; 
  assign frontend_io_ptw_pmp_5_cfg_w=ptw_io_requestor_1_pmp_5_cfg_w; 
  assign frontend_io_ptw_pmp_5_cfg_r=ptw_io_requestor_1_pmp_5_cfg_r; 
  assign frontend_io_ptw_pmp_5_addr=ptw_io_requestor_1_pmp_5_addr; 
  assign frontend_io_ptw_pmp_5_mask=ptw_io_requestor_1_pmp_5_mask; 
  assign frontend_io_ptw_pmp_6_cfg_l=ptw_io_requestor_1_pmp_6_cfg_l; 
  assign frontend_io_ptw_pmp_6_cfg_a=ptw_io_requestor_1_pmp_6_cfg_a; 
  assign frontend_io_ptw_pmp_6_cfg_x=ptw_io_requestor_1_pmp_6_cfg_x; 
  assign frontend_io_ptw_pmp_6_cfg_w=ptw_io_requestor_1_pmp_6_cfg_w; 
  assign frontend_io_ptw_pmp_6_cfg_r=ptw_io_requestor_1_pmp_6_cfg_r; 
  assign frontend_io_ptw_pmp_6_addr=ptw_io_requestor_1_pmp_6_addr; 
  assign frontend_io_ptw_pmp_6_mask=ptw_io_requestor_1_pmp_6_mask; 
  assign frontend_io_ptw_pmp_7_cfg_l=ptw_io_requestor_1_pmp_7_cfg_l; 
  assign frontend_io_ptw_pmp_7_cfg_a=ptw_io_requestor_1_pmp_7_cfg_a; 
  assign frontend_io_ptw_pmp_7_cfg_x=ptw_io_requestor_1_pmp_7_cfg_x; 
  assign frontend_io_ptw_pmp_7_cfg_w=ptw_io_requestor_1_pmp_7_cfg_w; 
  assign frontend_io_ptw_pmp_7_cfg_r=ptw_io_requestor_1_pmp_7_cfg_r; 
  assign frontend_io_ptw_pmp_7_addr=ptw_io_requestor_1_pmp_7_addr; 
  assign frontend_io_ptw_pmp_7_mask=ptw_io_requestor_1_pmp_7_mask; 
  assign frontend_io_ptw_customCSRs_csrs_0_value=ptw_io_requestor_1_customCSRs_csrs_0_value; 
  assign fpuOpt_clock=clock; 
  assign fpuOpt_reset=reset; 
  assign fpuOpt_io_inst=core_io_fpu_inst; 
  assign fpuOpt_io_fromint_data=core_io_fpu_fromint_data; 
  assign fpuOpt_io_fcsr_rm=core_io_fpu_fcsr_rm; 
  assign fpuOpt_io_dmem_resp_val=core_io_fpu_dmem_resp_val; 
  assign fpuOpt_io_dmem_resp_type=core_io_fpu_dmem_resp_type; 
  assign fpuOpt_io_dmem_resp_tag=core_io_fpu_dmem_resp_tag; 
  assign fpuOpt_io_dmem_resp_data=core_io_fpu_dmem_resp_data; 
  assign fpuOpt_io_valid=core_io_fpu_valid; 
  assign fpuOpt_io_killx=core_io_fpu_killx; 
  assign fpuOpt_io_killm=core_io_fpu_killm; 
  assign dcacheArb_clock=clock; 
  assign dcacheArb_io_requestor_0_req_valid=ptw_io_mem_req_valid; 
  assign dcacheArb_io_requestor_0_req_bits_addr=ptw_io_mem_req_bits_addr; 
  assign dcacheArb_io_requestor_0_s1_kill=ptw_io_mem_s1_kill; 
  assign dcacheArb_io_requestor_1_req_valid=core_io_dmem_req_valid; 
  assign dcacheArb_io_requestor_1_req_bits_addr=core_io_dmem_req_bits_addr; 
  assign dcacheArb_io_requestor_1_req_bits_tag=core_io_dmem_req_bits_tag; 
  assign dcacheArb_io_requestor_1_req_bits_cmd=core_io_dmem_req_bits_cmd; 
  assign dcacheArb_io_requestor_1_req_bits_size=core_io_dmem_req_bits_size; 
  assign dcacheArb_io_requestor_1_req_bits_signed=core_io_dmem_req_bits_signed; 
  assign dcacheArb_io_requestor_1_s1_kill=core_io_dmem_s1_kill; 
  assign dcacheArb_io_requestor_1_s1_data_data=core_io_dmem_s1_data_data; 
  assign dcacheArb_io_mem_req_ready=dcache_io_cpu_req_ready; 
  assign dcacheArb_io_mem_s2_nack=dcache_io_cpu_s2_nack; 
  assign dcacheArb_io_mem_resp_valid=dcache_io_cpu_resp_valid; 
  assign dcacheArb_io_mem_resp_bits_tag=dcache_io_cpu_resp_bits_tag; 
  assign dcacheArb_io_mem_resp_bits_size=dcache_io_cpu_resp_bits_size; 
  assign dcacheArb_io_mem_resp_bits_data=dcache_io_cpu_resp_bits_data; 
  assign dcacheArb_io_mem_resp_bits_replay=dcache_io_cpu_resp_bits_replay; 
  assign dcacheArb_io_mem_resp_bits_has_data=dcache_io_cpu_resp_bits_has_data; 
  assign dcacheArb_io_mem_resp_bits_data_word_bypass=dcache_io_cpu_resp_bits_data_word_bypass; 
  assign dcacheArb_io_mem_replay_next=dcache_io_cpu_replay_next; 
  assign dcacheArb_io_mem_s2_xcpt_ma_ld=dcache_io_cpu_s2_xcpt_ma_ld; 
  assign dcacheArb_io_mem_s2_xcpt_ma_st=dcache_io_cpu_s2_xcpt_ma_st; 
  assign dcacheArb_io_mem_s2_xcpt_pf_ld=dcache_io_cpu_s2_xcpt_pf_ld; 
  assign dcacheArb_io_mem_s2_xcpt_pf_st=dcache_io_cpu_s2_xcpt_pf_st; 
  assign dcacheArb_io_mem_s2_xcpt_ae_ld=dcache_io_cpu_s2_xcpt_ae_ld; 
  assign dcacheArb_io_mem_s2_xcpt_ae_st=dcache_io_cpu_s2_xcpt_ae_st; 
  assign dcacheArb_io_mem_ordered=dcache_io_cpu_ordered; 
  assign dcacheArb_io_mem_perf_release=dcache_io_cpu_perf_release; 
  assign dcacheArb_io_mem_perf_grant=dcache_io_cpu_perf_grant; 
  assign ptw_clock=clock; 
  assign ptw_reset=reset; 
  assign ptw_io_requestor_0_req_valid=dcache_io_ptw_req_valid; 
  assign ptw_io_requestor_0_req_bits_bits_addr=dcache_io_ptw_req_bits_bits_addr; 
  assign ptw_io_requestor_1_req_valid=frontend_io_ptw_req_valid; 
  assign ptw_io_requestor_1_req_bits_valid=frontend_io_ptw_req_bits_valid; 
  assign ptw_io_requestor_1_req_bits_bits_addr=frontend_io_ptw_req_bits_bits_addr; 
  assign ptw_io_mem_req_ready=dcacheArb_io_requestor_0_req_ready; 
  assign ptw_io_mem_s2_nack=dcacheArb_io_requestor_0_s2_nack; 
  assign ptw_io_mem_resp_valid=dcacheArb_io_requestor_0_resp_valid; 
  assign ptw_io_mem_resp_bits_data=dcacheArb_io_requestor_0_resp_bits_data; 
  assign ptw_io_mem_s2_xcpt_ae_ld=dcacheArb_io_requestor_0_s2_xcpt_ae_ld; 
  assign ptw_io_dpath_ptbr_mode=core_io_ptw_ptbr_mode; 
  assign ptw_io_dpath_ptbr_ppn=core_io_ptw_ptbr_ppn; 
  assign ptw_io_dpath_sfence_valid=core_io_ptw_sfence_valid; 
  assign ptw_io_dpath_sfence_bits_rs1=core_io_ptw_sfence_bits_rs1; 
  assign ptw_io_dpath_status_debug=core_io_ptw_status_debug; 
  assign ptw_io_dpath_status_dprv=core_io_ptw_status_dprv; 
  assign ptw_io_dpath_status_prv=core_io_ptw_status_prv; 
  assign ptw_io_dpath_status_mxr=core_io_ptw_status_mxr; 
  assign ptw_io_dpath_status_sum=core_io_ptw_status_sum; 
  assign ptw_io_dpath_pmp_0_cfg_l=core_io_ptw_pmp_0_cfg_l; 
  assign ptw_io_dpath_pmp_0_cfg_a=core_io_ptw_pmp_0_cfg_a; 
  assign ptw_io_dpath_pmp_0_cfg_x=core_io_ptw_pmp_0_cfg_x; 
  assign ptw_io_dpath_pmp_0_cfg_w=core_io_ptw_pmp_0_cfg_w; 
  assign ptw_io_dpath_pmp_0_cfg_r=core_io_ptw_pmp_0_cfg_r; 
  assign ptw_io_dpath_pmp_0_addr=core_io_ptw_pmp_0_addr; 
  assign ptw_io_dpath_pmp_0_mask=core_io_ptw_pmp_0_mask; 
  assign ptw_io_dpath_pmp_1_cfg_l=core_io_ptw_pmp_1_cfg_l; 
  assign ptw_io_dpath_pmp_1_cfg_a=core_io_ptw_pmp_1_cfg_a; 
  assign ptw_io_dpath_pmp_1_cfg_x=core_io_ptw_pmp_1_cfg_x; 
  assign ptw_io_dpath_pmp_1_cfg_w=core_io_ptw_pmp_1_cfg_w; 
  assign ptw_io_dpath_pmp_1_cfg_r=core_io_ptw_pmp_1_cfg_r; 
  assign ptw_io_dpath_pmp_1_addr=core_io_ptw_pmp_1_addr; 
  assign ptw_io_dpath_pmp_1_mask=core_io_ptw_pmp_1_mask; 
  assign ptw_io_dpath_pmp_2_cfg_l=core_io_ptw_pmp_2_cfg_l; 
  assign ptw_io_dpath_pmp_2_cfg_a=core_io_ptw_pmp_2_cfg_a; 
  assign ptw_io_dpath_pmp_2_cfg_x=core_io_ptw_pmp_2_cfg_x; 
  assign ptw_io_dpath_pmp_2_cfg_w=core_io_ptw_pmp_2_cfg_w; 
  assign ptw_io_dpath_pmp_2_cfg_r=core_io_ptw_pmp_2_cfg_r; 
  assign ptw_io_dpath_pmp_2_addr=core_io_ptw_pmp_2_addr; 
  assign ptw_io_dpath_pmp_2_mask=core_io_ptw_pmp_2_mask; 
  assign ptw_io_dpath_pmp_3_cfg_l=core_io_ptw_pmp_3_cfg_l; 
  assign ptw_io_dpath_pmp_3_cfg_a=core_io_ptw_pmp_3_cfg_a; 
  assign ptw_io_dpath_pmp_3_cfg_x=core_io_ptw_pmp_3_cfg_x; 
  assign ptw_io_dpath_pmp_3_cfg_w=core_io_ptw_pmp_3_cfg_w; 
  assign ptw_io_dpath_pmp_3_cfg_r=core_io_ptw_pmp_3_cfg_r; 
  assign ptw_io_dpath_pmp_3_addr=core_io_ptw_pmp_3_addr; 
  assign ptw_io_dpath_pmp_3_mask=core_io_ptw_pmp_3_mask; 
  assign ptw_io_dpath_pmp_4_cfg_l=core_io_ptw_pmp_4_cfg_l; 
  assign ptw_io_dpath_pmp_4_cfg_a=core_io_ptw_pmp_4_cfg_a; 
  assign ptw_io_dpath_pmp_4_cfg_x=core_io_ptw_pmp_4_cfg_x; 
  assign ptw_io_dpath_pmp_4_cfg_w=core_io_ptw_pmp_4_cfg_w; 
  assign ptw_io_dpath_pmp_4_cfg_r=core_io_ptw_pmp_4_cfg_r; 
  assign ptw_io_dpath_pmp_4_addr=core_io_ptw_pmp_4_addr; 
  assign ptw_io_dpath_pmp_4_mask=core_io_ptw_pmp_4_mask; 
  assign ptw_io_dpath_pmp_5_cfg_l=core_io_ptw_pmp_5_cfg_l; 
  assign ptw_io_dpath_pmp_5_cfg_a=core_io_ptw_pmp_5_cfg_a; 
  assign ptw_io_dpath_pmp_5_cfg_x=core_io_ptw_pmp_5_cfg_x; 
  assign ptw_io_dpath_pmp_5_cfg_w=core_io_ptw_pmp_5_cfg_w; 
  assign ptw_io_dpath_pmp_5_cfg_r=core_io_ptw_pmp_5_cfg_r; 
  assign ptw_io_dpath_pmp_5_addr=core_io_ptw_pmp_5_addr; 
  assign ptw_io_dpath_pmp_5_mask=core_io_ptw_pmp_5_mask; 
  assign ptw_io_dpath_pmp_6_cfg_l=core_io_ptw_pmp_6_cfg_l; 
  assign ptw_io_dpath_pmp_6_cfg_a=core_io_ptw_pmp_6_cfg_a; 
  assign ptw_io_dpath_pmp_6_cfg_x=core_io_ptw_pmp_6_cfg_x; 
  assign ptw_io_dpath_pmp_6_cfg_w=core_io_ptw_pmp_6_cfg_w; 
  assign ptw_io_dpath_pmp_6_cfg_r=core_io_ptw_pmp_6_cfg_r; 
  assign ptw_io_dpath_pmp_6_addr=core_io_ptw_pmp_6_addr; 
  assign ptw_io_dpath_pmp_6_mask=core_io_ptw_pmp_6_mask; 
  assign ptw_io_dpath_pmp_7_cfg_l=core_io_ptw_pmp_7_cfg_l; 
  assign ptw_io_dpath_pmp_7_cfg_a=core_io_ptw_pmp_7_cfg_a; 
  assign ptw_io_dpath_pmp_7_cfg_x=core_io_ptw_pmp_7_cfg_x; 
  assign ptw_io_dpath_pmp_7_cfg_w=core_io_ptw_pmp_7_cfg_w; 
  assign ptw_io_dpath_pmp_7_cfg_r=core_io_ptw_pmp_7_cfg_r; 
  assign ptw_io_dpath_pmp_7_addr=core_io_ptw_pmp_7_addr; 
  assign ptw_io_dpath_pmp_7_mask=core_io_ptw_pmp_7_mask; 
  assign ptw_io_dpath_customCSRs_csrs_0_value=core_io_ptw_customCSRs_csrs_0_value; 
  assign core_clock=clock; 
  assign core_reset=reset; 
  assign core_io_hartid=broadcast_auto_out; 
  assign core_io_interrupts_debug=intXbar_auto_int_out_0; 
  assign core_io_interrupts_mtip=intXbar_auto_int_out_2; 
  assign core_io_interrupts_msip=intXbar_auto_int_out_1; 
  assign core_io_interrupts_meip=intXbar_auto_int_out_3; 
  assign core_io_interrupts_seip=intXbar_auto_int_out_4; 
  assign core_io_imem_resp_valid=frontend_io_cpu_resp_valid; 
  assign core_io_imem_resp_bits_btb_taken=frontend_io_cpu_resp_bits_btb_taken; 
  assign core_io_imem_resp_bits_btb_bridx=frontend_io_cpu_resp_bits_btb_bridx; 
  assign core_io_imem_resp_bits_btb_entry=frontend_io_cpu_resp_bits_btb_entry; 
  assign core_io_imem_resp_bits_btb_bht_history=frontend_io_cpu_resp_bits_btb_bht_history; 
  assign core_io_imem_resp_bits_pc=frontend_io_cpu_resp_bits_pc; 
  assign core_io_imem_resp_bits_data=frontend_io_cpu_resp_bits_data; 
  assign core_io_imem_resp_bits_xcpt_pf_inst=frontend_io_cpu_resp_bits_xcpt_pf_inst; 
  assign core_io_imem_resp_bits_xcpt_ae_inst=frontend_io_cpu_resp_bits_xcpt_ae_inst; 
  assign core_io_imem_resp_bits_replay=frontend_io_cpu_resp_bits_replay; 
  assign core_io_dmem_req_ready=dcacheArb_io_requestor_1_req_ready; 
  assign core_io_dmem_s2_nack=dcacheArb_io_requestor_1_s2_nack; 
  assign core_io_dmem_resp_valid=dcacheArb_io_requestor_1_resp_valid; 
  assign core_io_dmem_resp_bits_tag=dcacheArb_io_requestor_1_resp_bits_tag; 
  assign core_io_dmem_resp_bits_size=dcacheArb_io_requestor_1_resp_bits_size; 
  assign core_io_dmem_resp_bits_data=dcacheArb_io_requestor_1_resp_bits_data; 
  assign core_io_dmem_resp_bits_replay=dcacheArb_io_requestor_1_resp_bits_replay; 
  assign core_io_dmem_resp_bits_has_data=dcacheArb_io_requestor_1_resp_bits_has_data; 
  assign core_io_dmem_resp_bits_data_word_bypass=dcacheArb_io_requestor_1_resp_bits_data_word_bypass; 
  assign core_io_dmem_replay_next=dcacheArb_io_requestor_1_replay_next; 
  assign core_io_dmem_s2_xcpt_ma_ld=dcacheArb_io_requestor_1_s2_xcpt_ma_ld; 
  assign core_io_dmem_s2_xcpt_ma_st=dcacheArb_io_requestor_1_s2_xcpt_ma_st; 
  assign core_io_dmem_s2_xcpt_pf_ld=dcacheArb_io_requestor_1_s2_xcpt_pf_ld; 
  assign core_io_dmem_s2_xcpt_pf_st=dcacheArb_io_requestor_1_s2_xcpt_pf_st; 
  assign core_io_dmem_s2_xcpt_ae_ld=dcacheArb_io_requestor_1_s2_xcpt_ae_ld; 
  assign core_io_dmem_s2_xcpt_ae_st=dcacheArb_io_requestor_1_s2_xcpt_ae_st; 
  assign core_io_dmem_ordered=dcacheArb_io_requestor_1_ordered; 
  assign core_io_dmem_perf_release=dcacheArb_io_requestor_1_perf_release; 
  assign core_io_dmem_perf_grant=dcacheArb_io_requestor_1_perf_grant; 
  assign core_io_fpu_fcsr_flags_valid=fpuOpt_io_fcsr_flags_valid; 
  assign core_io_fpu_fcsr_flags_bits=fpuOpt_io_fcsr_flags_bits; 
  assign core_io_fpu_store_data=fpuOpt_io_store_data; 
  assign core_io_fpu_toint_data=fpuOpt_io_toint_data; 
  assign core_io_fpu_fcsr_rdy=fpuOpt_io_fcsr_rdy; 
  assign core_io_fpu_nack_mem=fpuOpt_io_nack_mem; 
  assign core_io_fpu_illegal_rm=fpuOpt_io_illegal_rm; 
  assign core_io_fpu_dec_wen=fpuOpt_io_dec_wen; 
  assign core_io_fpu_dec_ren1=fpuOpt_io_dec_ren1; 
  assign core_io_fpu_dec_ren2=fpuOpt_io_dec_ren2; 
  assign core_io_fpu_dec_ren3=fpuOpt_io_dec_ren3; 
  assign core_io_fpu_sboard_set=fpuOpt_io_sboard_set; 
  assign core_io_fpu_sboard_clr=fpuOpt_io_sboard_clr; 
  assign core_io_fpu_sboard_clra=fpuOpt_io_sboard_clra; 
  assign RocketTile_covSum=30'h0; 
  assign tlMasterXbar_sum=RocketTile_covSum+tlMasterXbar_io_covSum; 
  assign intXbar_sum=tlMasterXbar_sum+intXbar_io_covSum; 
  assign fpuOpt_sum=intXbar_sum+fpuOpt_io_covSum; 
  assign dcacheArb_sum=fpuOpt_sum+dcacheArb_io_covSum; 
  assign frontend_sum=dcacheArb_sum+frontend_io_covSum; 
  assign dcache_sum=frontend_sum+dcache_io_covSum; 
  assign broadcast_3_sum=dcache_sum+broadcast_3_io_covSum; 
  assign core_sum=broadcast_3_sum+core_io_covSum; 
  assign broadcast_sum=core_sum+broadcast_io_covSum; 
  assign broadcast_1_sum=broadcast_sum+broadcast_1_io_covSum; 
  assign ptw_sum=broadcast_1_sum+ptw_io_covSum; 
  assign io_covSum=ptw_sum; 
  assign broadcast_1_metaAssert_wire=broadcast_1_metaAssert; 
  assign core_metaAssert_wire=core_metaAssert; 
  assign broadcast_metaAssert_wire=broadcast_metaAssert; 
  assign dcache_metaAssert_wire=dcache_metaAssert; 
  assign intXbar_metaAssert_wire=intXbar_metaAssert; 
  assign tlMasterXbar_metaAssert_wire=tlMasterXbar_metaAssert; 
  assign broadcast_3_metaAssert_wire=broadcast_3_metaAssert; 
  assign frontend_metaAssert_wire=frontend_metaAssert; 
  assign dcacheArb_metaAssert_wire=dcacheArb_metaAssert; 
  assign fpuOpt_metaAssert_wire=fpuOpt_metaAssert; 
  assign ptw_metaAssert_wire=ptw_metaAssert; 
  assign RocketTile_or3=tlMasterXbar_metaAssert_wire|broadcast_3_metaAssert_wire; 
  assign RocketTile_or10=dcache_metaAssert_wire|fpuOpt_metaAssert_wire; 
  assign RocketTile_or4=frontend_metaAssert_wire|RocketTile_or10; 
  assign RocketTile_or1=RocketTile_or3|RocketTile_or4; 
  assign RocketTile_or12=intXbar_metaAssert_wire|ptw_metaAssert_wire; 
  assign RocketTile_or5=broadcast_1_metaAssert_wire|RocketTile_or12; 
  assign RocketTile_or14=core_metaAssert_wire|dcacheArb_metaAssert_wire; 
  assign RocketTile_or6=broadcast_metaAssert_wire|RocketTile_or14; 
  assign RocketTile_or2=RocketTile_or5|RocketTile_or6; 
  assign RocketTile_or0=RocketTile_or1|RocketTile_or2; 
  assign metaAssert=RocketTile_metaAssert; 
  assign tlMasterXbar_metaReset=metaReset|tlMasterXbar_halt; 
  assign fpuOpt_metaReset=metaReset|fpuOpt_halt; 
  assign dcacheArb_metaReset=metaReset|dcacheArb_halt; 
  assign frontend_metaReset=metaReset|frontend_halt; 
  assign dcache_metaReset=metaReset|dcache_halt; 
  assign core_metaReset=metaReset|core_halt; 
  assign ptw_metaReset=metaReset|ptw_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              bundleOut_0_0_REG <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 bundleOut_0_0_REG <=1'h0;
               end 
             else 
               begin 
                 bundleOut_0_0_REG <=core_io_wfi;
               end 
         if (metaReset)
            begin 
              RocketTile_metaAssert <=1'h0;
            end 
          else 
            begin 
              RocketTile_metaAssert <=RocketTile_metaAssert|RocketTile_or0;
            end 
       end
  
endmodule
 
module TLXbar_7 (
  input clock,
  input reset,
  output auto_in_1_a_ready,
  input auto_in_1_a_valid,
  input [31:0] auto_in_1_a_bits_address,
  output auto_in_1_d_valid,
  output [2:0] auto_in_1_d_bits_opcode,
  output [3:0] auto_in_1_d_bits_size,
  output [63:0] auto_in_1_d_bits_data,
  output auto_in_1_d_bits_corrupt,
  output auto_in_0_a_ready,
  input auto_in_0_a_valid,
  input [2:0] auto_in_0_a_bits_opcode,
  input [2:0] auto_in_0_a_bits_param,
  input [3:0] auto_in_0_a_bits_size,
  input auto_in_0_a_bits_source,
  input [31:0] auto_in_0_a_bits_address,
  input [7:0] auto_in_0_a_bits_mask,
  input [63:0] auto_in_0_a_bits_data,
  input auto_in_0_b_ready,
  output auto_in_0_b_valid,
  output [1:0] auto_in_0_b_bits_param,
  output [3:0] auto_in_0_b_bits_size,
  output auto_in_0_b_bits_source,
  output [31:0] auto_in_0_b_bits_address,
  output auto_in_0_c_ready,
  input auto_in_0_c_valid,
  input [2:0] auto_in_0_c_bits_opcode,
  input [2:0] auto_in_0_c_bits_param,
  input [3:0] auto_in_0_c_bits_size,
  input auto_in_0_c_bits_source,
  input [31:0] auto_in_0_c_bits_address,
  input [63:0] auto_in_0_c_bits_data,
  input auto_in_0_d_ready,
  output auto_in_0_d_valid,
  output [2:0] auto_in_0_d_bits_opcode,
  output [1:0] auto_in_0_d_bits_param,
  output [3:0] auto_in_0_d_bits_size,
  output auto_in_0_d_bits_source,
  output [1:0] auto_in_0_d_bits_sink,
  output auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output auto_in_0_e_ready,
  input auto_in_0_e_valid,
  input [1:0] auto_in_0_e_bits_sink,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [1:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [2:0] auto_out_b_bits_opcode,
  input [1:0] auto_out_b_bits_param,
  input [3:0] auto_out_b_bits_size,
  input [1:0] auto_out_b_bits_source,
  input [31:0] auto_out_b_bits_address,
  input [7:0] auto_out_b_bits_mask,
  input auto_out_b_bits_corrupt,
  input auto_out_c_ready,
  output auto_out_c_valid,
  output [2:0] auto_out_c_bits_opcode,
  output [2:0] auto_out_c_bits_param,
  output [3:0] auto_out_c_bits_size,
  output [1:0] auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [1:0] auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt,
  input auto_out_e_ready,
  output auto_out_e_valid,
  output [1:0] auto_out_e_bits_sink,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input monitor_halt,
  input monitor_1_halt) ; 
   wire monitor_clock ;  
   wire monitor_reset ;  
   wire monitor_io_in_a_ready ;  
   wire monitor_io_in_a_valid ;  
   wire [2:0] monitor_io_in_a_bits_opcode ;  
   wire [2:0] monitor_io_in_a_bits_param ;  
   wire [3:0] monitor_io_in_a_bits_size ;  
   wire monitor_io_in_a_bits_source ;  
   wire [31:0] monitor_io_in_a_bits_address ;  
   wire [7:0] monitor_io_in_a_bits_mask ;  
   wire monitor_io_in_b_ready ;  
   wire monitor_io_in_b_valid ;  
   wire [2:0] monitor_io_in_b_bits_opcode ;  
   wire [1:0] monitor_io_in_b_bits_param ;  
   wire [3:0] monitor_io_in_b_bits_size ;  
   wire monitor_io_in_b_bits_source ;  
   wire [31:0] monitor_io_in_b_bits_address ;  
   wire [7:0] monitor_io_in_b_bits_mask ;  
   wire monitor_io_in_b_bits_corrupt ;  
   wire monitor_io_in_c_ready ;  
   wire monitor_io_in_c_valid ;  
   wire [2:0] monitor_io_in_c_bits_opcode ;  
   wire [2:0] monitor_io_in_c_bits_param ;  
   wire [3:0] monitor_io_in_c_bits_size ;  
   wire monitor_io_in_c_bits_source ;  
   wire [31:0] monitor_io_in_c_bits_address ;  
   wire monitor_io_in_d_ready ;  
   wire monitor_io_in_d_valid ;  
   wire [2:0] monitor_io_in_d_bits_opcode ;  
   wire [1:0] monitor_io_in_d_bits_param ;  
   wire [3:0] monitor_io_in_d_bits_size ;  
   wire monitor_io_in_d_bits_source ;  
   wire [1:0] monitor_io_in_d_bits_sink ;  
   wire monitor_io_in_d_bits_denied ;  
   wire monitor_io_in_d_bits_corrupt ;  
   wire monitor_io_in_e_ready ;  
   wire monitor_io_in_e_valid ;  
   wire [1:0] monitor_io_in_e_bits_sink ;  
   wire [29:0] monitor_io_covSum ;  
   wire monitor_metaAssert ;  
   wire monitor_metaReset ;  
   wire monitor_1_clock ;  
   wire monitor_1_reset ;  
   wire monitor_1_io_in_a_ready ;  
   wire monitor_1_io_in_a_valid ;  
   wire [31:0] monitor_1_io_in_a_bits_address ;  
   wire monitor_1_io_in_d_valid ;  
   wire [2:0] monitor_1_io_in_d_bits_opcode ;  
   wire [1:0] monitor_1_io_in_d_bits_param ;  
   wire [3:0] monitor_1_io_in_d_bits_size ;  
   wire [1:0] monitor_1_io_in_d_bits_sink ;  
   wire monitor_1_io_in_d_bits_denied ;  
   wire monitor_1_io_in_d_bits_corrupt ;  
   wire [29:0] monitor_1_io_covSum ;  
   wire monitor_1_metaAssert ;  
   wire monitor_1_metaReset ;  
   wire requestBOI_0_0 ;  
   wire requestDOI_0_0 ;  
   wire requestDOI_0_1 ;  
   wire [26:0] _beatsAI_decode_T_1 ;  
   wire [8:0] beatsAI_decode ;  
   wire beatsAI_opdata ;  
   wire _portsDIO_out_0_d_ready_T ;  
   reg [8:0] beatsLeft ;  
   reg [31:0] _RAND_0 ;  
   wire idle ;  
   wire latch ;  
   wire [1:0] readys_filter_lo ;  
   wire _readys_T_1 ;  
   wire _readys_T_3 ;  
   reg [1:0] readys_mask ;  
   reg [31:0] _RAND_1 ;  
   wire [1:0] readys_filter_hi ;  
   wire [3:0] readys_filter ;  
   wire [3:0] _GEN_1 ;  
   wire [3:0] _readys_unready_T_1 ;  
   wire [3:0] _readys_unready_T_4 ;  
   wire [3:0] _GEN_2 ;  
   wire [3:0] readys_unready ;  
   wire [1:0] _readys_readys_T_2 ;  
   wire [1:0] readys_readys ;  
   wire _readys_T_5 ;  
   wire _readys_T_6 ;  
   wire [1:0] _readys_mask_T ;  
   wire [2:0] _readys_mask_T_1 ;  
   wire [1:0] _readys_mask_T_3 ;  
   wire readys_0 ;  
   wire readys_1 ;  
   wire earlyWinner_0 ;  
   wire earlyWinner_1 ;  
   wire _prefixOR_T ;  
   wire _T_6 ;  
   wire _T_9 ;  
   wire _T_11 ;  
   wire _T_14 ;  
   wire _T_16 ;  
   wire _T_21 ;  
   wire _T_23 ;  
   reg state_0 ;  
   reg [31:0] _RAND_2 ;  
   wire muxStateEarly_0 ;  
   reg state_1 ;  
   reg [31:0] _RAND_3 ;  
   wire muxStateEarly_1 ;  
   wire _out_0_a_earlyValid_T_1 ;  
   wire _out_0_a_earlyValid_T_2 ;  
   wire _out_0_a_earlyValid_T_3 ;  
   wire out_2_0_a_earlyValid ;  
   wire _beatsLeft_T_2 ;  
   wire [8:0] _GEN_3 ;  
   wire [8:0] _beatsLeft_T_4 ;  
   wire allowed_0 ;  
   wire allowed_1 ;  
   wire [7:0] _T_31 ;  
   wire [7:0] _T_32 ;  
   wire [31:0] _T_34 ;  
   wire [31:0] _T_35 ;  
   wire [1:0] in_0_a_bits_source ;  
   wire [1:0] _T_37 ;  
   wire [1:0] _T_38 ;  
   wire [3:0] _T_40 ;  
   wire [3:0] _T_41 ;  
   wire [2:0] _T_46 ;  
   wire [2:0] _T_47 ;  
   reg [2:0] TLXbar_7_state ;  
   reg [31:0] _RAND_4 ;  
   reg TLXbar_7_cov[0:7] ;  
   reg [31:0] _RAND_5 ;  
   wire TLXbar_7_cov_read_data ;  
   wire [2:0] TLXbar_7_cov_read_addr ;  
   wire TLXbar_7_cov_write_data ;  
   wire [2:0] TLXbar_7_cov_write_addr ;  
   wire TLXbar_7_cov_write_mask ;  
   wire TLXbar_7_cov_write_en ;  
   reg [29:0] TLXbar_7_covSum ;  
   reg [31:0] _RAND_6 ;  
   wire [1:0] readys_mask_shl ;  
   wire [2:0] readys_mask_pad ;  
   wire [2:0] state_0_shl ;  
   wire [2:0] state_0_pad ;  
   wire [2:0] state_1_shl ;  
   wire [2:0] state_1_pad ;  
   wire [2:0] TLXbar_7_xor2 ;  
   wire [2:0] TLXbar_7_xor0 ;  
   wire [29:0] monitor_sum ;  
   wire [29:0] monitor_1_sum ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire stopEn2 ;  
   wire stopEn3 ;  
   wire monitor_metaAssert_wire ;  
   wire monitor_1_metaAssert_wire ;  
   wire TLXbar_7_or4 ;  
   wire TLXbar_7_or1 ;  
   wire TLXbar_7_or6 ;  
   wire TLXbar_7_or2 ;  
   wire TLXbar_7_or0 ;  
   reg TLXbar_7_metaAssert ;  
   reg [31:0] _RAND_7 ;  
  TLMonitor_23 monitor(.clock(monitor_clock),.reset(monitor_reset),.io_in_a_ready(monitor_io_in_a_ready),.io_in_a_valid(monitor_io_in_a_valid),.io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),.io_in_a_bits_param(monitor_io_in_a_bits_param),.io_in_a_bits_size(monitor_io_in_a_bits_size),.io_in_a_bits_source(monitor_io_in_a_bits_source),.io_in_a_bits_address(monitor_io_in_a_bits_address),.io_in_a_bits_mask(monitor_io_in_a_bits_mask),.io_in_b_ready(monitor_io_in_b_ready),.io_in_b_valid(monitor_io_in_b_valid),.io_in_b_bits_opcode(monitor_io_in_b_bits_opcode),.io_in_b_bits_param(monitor_io_in_b_bits_param),.io_in_b_bits_size(monitor_io_in_b_bits_size),.io_in_b_bits_source(monitor_io_in_b_bits_source),.io_in_b_bits_address(monitor_io_in_b_bits_address),.io_in_b_bits_mask(monitor_io_in_b_bits_mask),.io_in_b_bits_corrupt(monitor_io_in_b_bits_corrupt),.io_in_c_ready(monitor_io_in_c_ready),.io_in_c_valid(monitor_io_in_c_valid),.io_in_c_bits_opcode(monitor_io_in_c_bits_opcode),.io_in_c_bits_param(monitor_io_in_c_bits_param),.io_in_c_bits_size(monitor_io_in_c_bits_size),.io_in_c_bits_source(monitor_io_in_c_bits_source),.io_in_c_bits_address(monitor_io_in_c_bits_address),.io_in_d_ready(monitor_io_in_d_ready),.io_in_d_valid(monitor_io_in_d_valid),.io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),.io_in_d_bits_param(monitor_io_in_d_bits_param),.io_in_d_bits_size(monitor_io_in_d_bits_size),.io_in_d_bits_source(monitor_io_in_d_bits_source),.io_in_d_bits_sink(monitor_io_in_d_bits_sink),.io_in_d_bits_denied(monitor_io_in_d_bits_denied),.io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt),.io_in_e_ready(monitor_io_in_e_ready),.io_in_e_valid(monitor_io_in_e_valid),.io_in_e_bits_sink(monitor_io_in_e_bits_sink),.io_covSum(monitor_io_covSum),.metaAssert(monitor_metaAssert),.metaReset(monitor_metaReset)); 
  TLMonitor_24 monitor_1(.clock(monitor_1_clock),.reset(monitor_1_reset),.io_in_a_ready(monitor_1_io_in_a_ready),.io_in_a_valid(monitor_1_io_in_a_valid),.io_in_a_bits_address(monitor_1_io_in_a_bits_address),.io_in_d_valid(monitor_1_io_in_d_valid),.io_in_d_bits_opcode(monitor_1_io_in_d_bits_opcode),.io_in_d_bits_param(monitor_1_io_in_d_bits_param),.io_in_d_bits_size(monitor_1_io_in_d_bits_size),.io_in_d_bits_sink(monitor_1_io_in_d_bits_sink),.io_in_d_bits_denied(monitor_1_io_in_d_bits_denied),.io_in_d_bits_corrupt(monitor_1_io_in_d_bits_corrupt),.io_covSum(monitor_1_io_covSum),.metaAssert(monitor_1_metaAssert),.metaReset(monitor_1_metaReset)); 
  assign requestBOI_0_0=~auto_out_b_bits_source[1]; 
  assign requestDOI_0_0=~auto_out_d_bits_source[1]; 
  assign requestDOI_0_1=auto_out_d_bits_source==2'h2; 
  assign _beatsAI_decode_T_1=27'hfff<<auto_in_0_a_bits_size; 
  assign beatsAI_decode=~_beatsAI_decode_T_1[11:3]; 
  assign beatsAI_opdata=~auto_in_0_a_bits_opcode[2]; 
  assign _portsDIO_out_0_d_ready_T=requestDOI_0_0&auto_in_0_d_ready; 
  assign idle=beatsLeft==9'h0; 
  assign latch=idle&auto_out_a_ready; 
  assign readys_filter_lo={auto_in_1_a_valid,auto_in_0_a_valid}; 
  assign _readys_T_1=readys_filter_lo==readys_filter_lo; 
  assign _readys_T_3=_readys_T_1|reset; 
  assign readys_filter_hi=readys_filter_lo&~readys_mask; 
  assign readys_filter={readys_filter_hi,auto_in_1_a_valid,auto_in_0_a_valid}; 
  assign _GEN_1={1'b0,readys_filter[3:1]}; 
  assign _readys_unready_T_1=readys_filter|_GEN_1; 
  assign _readys_unready_T_4={readys_mask,2'h0}; 
  assign _GEN_2={1'b0,_readys_unready_T_1[3:1]}; 
  assign readys_unready=_GEN_2|_readys_unready_T_4; 
  assign _readys_readys_T_2=readys_unready[3:2]&readys_unready[1:0]; 
  assign readys_readys=~_readys_readys_T_2; 
  assign _readys_T_5=|readys_filter_lo; 
  assign _readys_T_6=latch&_readys_T_5; 
  assign _readys_mask_T=readys_readys&readys_filter_lo; 
  assign _readys_mask_T_1={_readys_mask_T,1'h0}; 
  assign _readys_mask_T_3=_readys_mask_T|_readys_mask_T_1[1:0]; 
  assign readys_0=readys_readys[0]; 
  assign readys_1=readys_readys[1]; 
  assign earlyWinner_0=readys_0&auto_in_0_a_valid; 
  assign earlyWinner_1=readys_1&auto_in_1_a_valid; 
  assign _prefixOR_T=earlyWinner_0|earlyWinner_1; 
  assign _T_6=~earlyWinner_0|~earlyWinner_1; 
  assign _T_9=_T_6|reset; 
  assign _T_11=auto_in_0_a_valid|auto_in_1_a_valid; 
  assign _T_14=~_T_11|_prefixOR_T; 
  assign _T_16=_T_14|reset; 
  assign _T_21=~_T_11|_T_11; 
  assign _T_23=_T_21|reset; 
  assign muxStateEarly_0=idle ? earlyWinner_0:state_0; 
  assign muxStateEarly_1=idle ? earlyWinner_1:state_1; 
  assign _out_0_a_earlyValid_T_1=state_0&auto_in_0_a_valid; 
  assign _out_0_a_earlyValid_T_2=state_1&auto_in_1_a_valid; 
  assign _out_0_a_earlyValid_T_3=_out_0_a_earlyValid_T_1|_out_0_a_earlyValid_T_2; 
  assign out_2_0_a_earlyValid=idle ? _T_11:_out_0_a_earlyValid_T_3; 
  assign _beatsLeft_T_2=auto_out_a_ready&out_2_0_a_earlyValid; 
  assign _GEN_3={8'b0,_beatsLeft_T_2}; 
  assign _beatsLeft_T_4=beatsLeft-_GEN_3; 
  assign allowed_0=idle ? readys_0:state_0; 
  assign allowed_1=idle ? readys_1:state_1; 
  assign _T_31=muxStateEarly_0 ? auto_in_0_a_bits_mask:8'h0; 
  assign _T_32=muxStateEarly_1 ? 8'hff:8'h0; 
  assign _T_34=muxStateEarly_0 ? auto_in_0_a_bits_address:32'h0; 
  assign _T_35=muxStateEarly_1 ? auto_in_1_a_bits_address:32'h0; 
  assign in_0_a_bits_source={1'b0,auto_in_0_a_bits_source}; 
  assign _T_37=muxStateEarly_0 ? in_0_a_bits_source:2'h0; 
  assign _T_38=muxStateEarly_1 ? 2'h2:2'h0; 
  assign _T_40=muxStateEarly_0 ? auto_in_0_a_bits_size:4'h0; 
  assign _T_41=muxStateEarly_1 ? 4'h6:4'h0; 
  assign _T_46=muxStateEarly_0 ? auto_in_0_a_bits_opcode:3'h0; 
  assign _T_47=muxStateEarly_1 ? 3'h4:3'h0; 
  assign auto_in_1_a_ready=auto_out_a_ready&allowed_1; 
  assign auto_in_1_d_valid=auto_out_d_valid&requestDOI_0_1; 
  assign auto_in_1_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_1_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_1_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_1_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign auto_in_0_a_ready=auto_out_a_ready&allowed_0; 
  assign auto_in_0_b_valid=auto_out_b_valid&requestBOI_0_0; 
  assign auto_in_0_b_bits_param=auto_out_b_bits_param; 
  assign auto_in_0_b_bits_size=auto_out_b_bits_size; 
  assign auto_in_0_b_bits_source=auto_out_b_bits_source[0]; 
  assign auto_in_0_b_bits_address=auto_out_b_bits_address; 
  assign auto_in_0_c_ready=auto_out_c_ready; 
  assign auto_in_0_d_valid=auto_out_d_valid&requestDOI_0_0; 
  assign auto_in_0_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_0_d_bits_param=auto_out_d_bits_param; 
  assign auto_in_0_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_0_d_bits_source=auto_out_d_bits_source[0]; 
  assign auto_in_0_d_bits_sink=auto_out_d_bits_sink; 
  assign auto_in_0_d_bits_denied=auto_out_d_bits_denied; 
  assign auto_in_0_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_0_e_ready=auto_out_e_ready; 
  assign auto_out_a_valid=idle ? _T_11:_out_0_a_earlyValid_T_3; 
  assign auto_out_a_bits_opcode=_T_46|_T_47; 
  assign auto_out_a_bits_param=muxStateEarly_0 ? auto_in_0_a_bits_param:3'h0; 
  assign auto_out_a_bits_size=_T_40|_T_41; 
  assign auto_out_a_bits_source=_T_37|_T_38; 
  assign auto_out_a_bits_address=_T_34|_T_35; 
  assign auto_out_a_bits_mask=_T_31|_T_32; 
  assign auto_out_a_bits_data=muxStateEarly_0 ? auto_in_0_a_bits_data:64'h0; 
  assign auto_out_b_ready=requestBOI_0_0&auto_in_0_b_ready; 
  assign auto_out_c_valid=auto_in_0_c_valid; 
  assign auto_out_c_bits_opcode=auto_in_0_c_bits_opcode; 
  assign auto_out_c_bits_param=auto_in_0_c_bits_param; 
  assign auto_out_c_bits_size=auto_in_0_c_bits_size; 
  assign auto_out_c_bits_source={1'b0,auto_in_0_c_bits_source}; 
  assign auto_out_c_bits_address=auto_in_0_c_bits_address; 
  assign auto_out_c_bits_data=auto_in_0_c_bits_data; 
  assign auto_out_d_ready=_portsDIO_out_0_d_ready_T|requestDOI_0_1; 
  assign auto_out_e_valid=auto_in_0_e_valid; 
  assign auto_out_e_bits_sink=auto_in_0_e_bits_sink; 
  assign monitor_clock=clock; 
  assign monitor_reset=reset; 
  assign monitor_io_in_a_ready=auto_out_a_ready&allowed_0; 
  assign monitor_io_in_a_valid=auto_in_0_a_valid; 
  assign monitor_io_in_a_bits_opcode=auto_in_0_a_bits_opcode; 
  assign monitor_io_in_a_bits_param=auto_in_0_a_bits_param; 
  assign monitor_io_in_a_bits_size=auto_in_0_a_bits_size; 
  assign monitor_io_in_a_bits_source=auto_in_0_a_bits_source; 
  assign monitor_io_in_a_bits_address=auto_in_0_a_bits_address; 
  assign monitor_io_in_a_bits_mask=auto_in_0_a_bits_mask; 
  assign monitor_io_in_b_ready=auto_in_0_b_ready; 
  assign monitor_io_in_b_valid=auto_out_b_valid&requestBOI_0_0; 
  assign monitor_io_in_b_bits_opcode=auto_out_b_bits_opcode; 
  assign monitor_io_in_b_bits_param=auto_out_b_bits_param; 
  assign monitor_io_in_b_bits_size=auto_out_b_bits_size; 
  assign monitor_io_in_b_bits_source=auto_out_b_bits_source[0]; 
  assign monitor_io_in_b_bits_address=auto_out_b_bits_address; 
  assign monitor_io_in_b_bits_mask=auto_out_b_bits_mask; 
  assign monitor_io_in_b_bits_corrupt=auto_out_b_bits_corrupt; 
  assign monitor_io_in_c_ready=auto_out_c_ready; 
  assign monitor_io_in_c_valid=auto_in_0_c_valid; 
  assign monitor_io_in_c_bits_opcode=auto_in_0_c_bits_opcode; 
  assign monitor_io_in_c_bits_param=auto_in_0_c_bits_param; 
  assign monitor_io_in_c_bits_size=auto_in_0_c_bits_size; 
  assign monitor_io_in_c_bits_source=auto_in_0_c_bits_source; 
  assign monitor_io_in_c_bits_address=auto_in_0_c_bits_address; 
  assign monitor_io_in_d_ready=auto_in_0_d_ready; 
  assign monitor_io_in_d_valid=auto_out_d_valid&requestDOI_0_0; 
  assign monitor_io_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign monitor_io_in_d_bits_param=auto_out_d_bits_param; 
  assign monitor_io_in_d_bits_size=auto_out_d_bits_size; 
  assign monitor_io_in_d_bits_source=auto_out_d_bits_source[0]; 
  assign monitor_io_in_d_bits_sink=auto_out_d_bits_sink; 
  assign monitor_io_in_d_bits_denied=auto_out_d_bits_denied; 
  assign monitor_io_in_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign monitor_io_in_e_ready=auto_out_e_ready; 
  assign monitor_io_in_e_valid=auto_in_0_e_valid; 
  assign monitor_io_in_e_bits_sink=auto_in_0_e_bits_sink; 
  assign monitor_1_clock=clock; 
  assign monitor_1_reset=reset; 
  assign monitor_1_io_in_a_ready=auto_out_a_ready&allowed_1; 
  assign monitor_1_io_in_a_valid=auto_in_1_a_valid; 
  assign monitor_1_io_in_a_bits_address=auto_in_1_a_bits_address; 
  assign monitor_1_io_in_d_valid=auto_out_d_valid&requestDOI_0_1; 
  assign monitor_1_io_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign monitor_1_io_in_d_bits_param=auto_out_d_bits_param; 
  assign monitor_1_io_in_d_bits_size=auto_out_d_bits_size; 
  assign monitor_1_io_in_d_bits_sink=auto_out_d_bits_sink; 
  assign monitor_1_io_in_d_bits_denied=auto_out_d_bits_denied; 
  assign monitor_1_io_in_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign TLXbar_7_cov_read_addr=TLXbar_7_state; 
  assign TLXbar_7_cov_read_data=TLXbar_7_cov[TLXbar_7_cov_read_addr]; 
  assign TLXbar_7_cov_write_data=1'h1; 
  assign TLXbar_7_cov_write_addr=TLXbar_7_state; 
  assign TLXbar_7_cov_write_mask=1'h1; 
  assign TLXbar_7_cov_write_en=1'h1; 
  assign readys_mask_shl=readys_mask; 
  assign readys_mask_pad={1'h0,readys_mask_shl}; 
  assign state_0_shl={state_0,2'h0}; 
  assign state_0_pad=state_0_shl; 
  assign state_1_shl={state_1,2'h0}; 
  assign state_1_pad=state_1_shl; 
  assign TLXbar_7_xor2=state_0_pad^state_1_pad; 
  assign TLXbar_7_xor0=readys_mask_pad^TLXbar_7_xor2; 
  assign monitor_sum=TLXbar_7_covSum+monitor_io_covSum; 
  assign monitor_1_sum=monitor_sum+monitor_1_io_covSum; 
  assign io_covSum=monitor_1_sum; 
  assign stopEn0=~_readys_T_3; 
  assign stopEn1=~_T_9; 
  assign stopEn2=~_T_16; 
  assign stopEn3=~_T_23; 
  assign monitor_metaAssert_wire=monitor_metaAssert; 
  assign monitor_1_metaAssert_wire=monitor_1_metaAssert; 
  assign TLXbar_7_or4=stopEn1|stopEn2; 
  assign TLXbar_7_or1=stopEn0|TLXbar_7_or4; 
  assign TLXbar_7_or6=monitor_metaAssert_wire|monitor_1_metaAssert_wire; 
  assign TLXbar_7_or2=stopEn3|TLXbar_7_or6; 
  assign TLXbar_7_or0=TLXbar_7_or1|TLXbar_7_or2; 
  assign metaAssert=TLXbar_7_metaAssert; 
  assign monitor_metaReset=metaReset|monitor_halt; 
  assign monitor_1_metaReset=metaReset|monitor_1_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              beatsLeft <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 beatsLeft <=9'h0;
               end 
             else 
               if (latch)
                  begin 
                    if (earlyWinner_0)
                       begin 
                         if (beatsAI_opdata)
                            begin 
                              beatsLeft <=beatsAI_decode;
                            end 
                          else 
                            begin 
                              beatsLeft <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         beatsLeft <=9'h0;
                       end 
                  end 
                else 
                  begin 
                    beatsLeft <=_beatsLeft_T_4;
                  end 
         if (metaReset)
            begin 
              readys_mask <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 readys_mask <=2'h3;
               end 
             else 
               if (_readys_T_6)
                  begin 
                    readys_mask <=_readys_mask_T_3;
                  end 
         if (metaReset)
            begin 
              state_0 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_0 <=1'h0;
               end 
             else 
               if (idle)
                  begin 
                    state_0 <=earlyWinner_0;
                  end 
         if (metaReset)
            begin 
              state_1 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_1 <=1'h0;
               end 
             else 
               if (idle)
                  begin 
                    state_1 <=earlyWinner_1;
                  end 
         if (~_readys_T_3)
            begin $display("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");
            end 
         if (~_readys_T_3)
            begin $display("fatal");
            end 
         if (~_T_9)
            begin $display("Assertion failed\n    at Arbiter.scala:105 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
            end 
         if (~_T_9)
            begin $display("fatal");
            end 
         if (~_T_16)
            begin $display("Assertion failed\n    at Arbiter.scala:107 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n");
            end 
         if (~_T_16)
            begin $display("fatal");
            end 
         if (~_T_23)
            begin $display("Assertion failed\n    at Arbiter.scala:108 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n");
            end 
         if (~_T_23)
            begin $display("fatal");
            end 
         TLXbar_7_state <=TLXbar_7_xor0;
         if (!(TLXbar_7_cov_read_data))
            begin 
              TLXbar_7_covSum <=TLXbar_7_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              TLXbar_7_metaAssert <=1'h0;
            end 
          else 
            begin 
              TLXbar_7_metaAssert <=TLXbar_7_metaAssert|TLXbar_7_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (TLXbar_7_cov_write_en&TLXbar_7_cov_write_mask)
            begin 
              TLXbar_7_cov [TLXbar_7_cov_write_addr]<=TLXbar_7_cov_write_data;
            end 
       end
  
endmodule
 
module IntXbar_1 (
  input auto_int_in_3_0,
  input auto_int_in_2_0,
  input auto_int_in_1_0,
  input auto_int_in_1_1,
  input auto_int_in_0_0,
  output auto_int_out_0,
  output auto_int_out_1,
  output auto_int_out_2,
  output auto_int_out_3,
  output auto_int_out_4,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [29:0] IntXbar_1_covSum ;  
  assign auto_int_out_0=auto_int_in_0_0; 
  assign auto_int_out_1=auto_int_in_1_0; 
  assign auto_int_out_2=auto_int_in_1_1; 
  assign auto_int_out_3=auto_int_in_2_0; 
  assign auto_int_out_4=auto_int_in_3_0; 
  assign IntXbar_1_covSum=30'h0; 
  assign io_covSum=IntXbar_1_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module BundleBridgeNexus_6 (
  input auto_in,
  output auto_out,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [29:0] BundleBridgeNexus_6_covSum ;  
  assign auto_out=auto_in; 
  assign BundleBridgeNexus_6_covSum=30'h0; 
  assign io_covSum=BundleBridgeNexus_6_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module BundleBridgeNexus_7 (
  input [31:0] auto_in,
  output [31:0] auto_out_1,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [29:0] BundleBridgeNexus_7_covSum ;  
  assign auto_out_1=auto_in; 
  assign BundleBridgeNexus_7_covSum=30'h0; 
  assign io_covSum=BundleBridgeNexus_7_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module BundleBridgeNexus_10 (
  input auto_in_0_valid,
  input [39:0] auto_in_0_iaddr,
  input [31:0] auto_in_0_insn,
  input [2:0] auto_in_0_priv,
  input auto_in_0_exception,
  input auto_in_0_interrupt,
  input [63:0] auto_in_0_cause,
  input [39:0] auto_in_0_tval,
  output auto_out_0_valid,
  output [39:0] auto_out_0_iaddr,
  output [31:0] auto_out_0_insn,
  output [2:0] auto_out_0_priv,
  output auto_out_0_exception,
  output auto_out_0_interrupt,
  output [63:0] auto_out_0_cause,
  output [39:0] auto_out_0_tval,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [29:0] BundleBridgeNexus_10_covSum ;  
  assign auto_out_0_valid=auto_in_0_valid; 
  assign auto_out_0_iaddr=auto_in_0_iaddr; 
  assign auto_out_0_insn=auto_in_0_insn; 
  assign auto_out_0_priv=auto_in_0_priv; 
  assign auto_out_0_exception=auto_in_0_exception; 
  assign auto_out_0_interrupt=auto_in_0_interrupt; 
  assign auto_out_0_cause=auto_in_0_cause; 
  assign auto_out_0_tval=auto_in_0_tval; 
  assign BundleBridgeNexus_10_covSum=30'h0; 
  assign io_covSum=BundleBridgeNexus_10_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module DCache (
  input gated_clock,
  input reset,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [1:0] auto_out_b_bits_param,
  input [3:0] auto_out_b_bits_size,
  input auto_out_b_bits_source,
  input [31:0] auto_out_b_bits_address,
  input auto_out_c_ready,
  output auto_out_c_valid,
  output [2:0] auto_out_c_bits_opcode,
  output [2:0] auto_out_c_bits_param,
  output [3:0] auto_out_c_bits_size,
  output auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_e_ready,
  output auto_out_e_valid,
  output [1:0] auto_out_e_bits_sink,
  output io_cpu_req_ready,
  input io_cpu_req_valid,
  input [39:0] io_cpu_req_bits_addr,
  input [6:0] io_cpu_req_bits_tag,
  input [4:0] io_cpu_req_bits_cmd,
  input [1:0] io_cpu_req_bits_size,
  input io_cpu_req_bits_signed,
  input io_cpu_req_bits_phys,
  input io_cpu_s1_kill,
  input [63:0] io_cpu_s1_data_data,
  output io_cpu_s2_nack,
  output io_cpu_resp_valid,
  output [6:0] io_cpu_resp_bits_tag,
  output [1:0] io_cpu_resp_bits_size,
  output [63:0] io_cpu_resp_bits_data,
  output io_cpu_resp_bits_replay,
  output io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output io_cpu_replay_next,
  output io_cpu_s2_xcpt_ma_ld,
  output io_cpu_s2_xcpt_ma_st,
  output io_cpu_s2_xcpt_pf_ld,
  output io_cpu_s2_xcpt_pf_st,
  output io_cpu_s2_xcpt_ae_ld,
  output io_cpu_s2_xcpt_ae_st,
  output io_cpu_ordered,
  output io_cpu_perf_release,
  output io_cpu_perf_grant,
  input io_ptw_req_ready,
  output io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input io_ptw_resp_valid,
  input io_ptw_resp_bits_ae,
  input [53:0] io_ptw_resp_bits_pte_ppn,
  input io_ptw_resp_bits_pte_d,
  input io_ptw_resp_bits_pte_a,
  input io_ptw_resp_bits_pte_g,
  input io_ptw_resp_bits_pte_u,
  input io_ptw_resp_bits_pte_x,
  input io_ptw_resp_bits_pte_w,
  input io_ptw_resp_bits_pte_r,
  input io_ptw_resp_bits_pte_v,
  input [1:0] io_ptw_resp_bits_level,
  input io_ptw_resp_bits_homogeneous,
  input [3:0] io_ptw_ptbr_mode,
  input io_ptw_status_debug,
  input [1:0] io_ptw_status_dprv,
  input io_ptw_status_mxr,
  input io_ptw_status_sum,
  input io_ptw_pmp_0_cfg_l,
  input [1:0] io_ptw_pmp_0_cfg_a,
  input io_ptw_pmp_0_cfg_x,
  input io_ptw_pmp_0_cfg_w,
  input io_ptw_pmp_0_cfg_r,
  input [29:0] io_ptw_pmp_0_addr,
  input [31:0] io_ptw_pmp_0_mask,
  input io_ptw_pmp_1_cfg_l,
  input [1:0] io_ptw_pmp_1_cfg_a,
  input io_ptw_pmp_1_cfg_x,
  input io_ptw_pmp_1_cfg_w,
  input io_ptw_pmp_1_cfg_r,
  input [29:0] io_ptw_pmp_1_addr,
  input [31:0] io_ptw_pmp_1_mask,
  input io_ptw_pmp_2_cfg_l,
  input [1:0] io_ptw_pmp_2_cfg_a,
  input io_ptw_pmp_2_cfg_x,
  input io_ptw_pmp_2_cfg_w,
  input io_ptw_pmp_2_cfg_r,
  input [29:0] io_ptw_pmp_2_addr,
  input [31:0] io_ptw_pmp_2_mask,
  input io_ptw_pmp_3_cfg_l,
  input [1:0] io_ptw_pmp_3_cfg_a,
  input io_ptw_pmp_3_cfg_x,
  input io_ptw_pmp_3_cfg_w,
  input io_ptw_pmp_3_cfg_r,
  input [29:0] io_ptw_pmp_3_addr,
  input [31:0] io_ptw_pmp_3_mask,
  input io_ptw_pmp_4_cfg_l,
  input [1:0] io_ptw_pmp_4_cfg_a,
  input io_ptw_pmp_4_cfg_x,
  input io_ptw_pmp_4_cfg_w,
  input io_ptw_pmp_4_cfg_r,
  input [29:0] io_ptw_pmp_4_addr,
  input [31:0] io_ptw_pmp_4_mask,
  input io_ptw_pmp_5_cfg_l,
  input [1:0] io_ptw_pmp_5_cfg_a,
  input io_ptw_pmp_5_cfg_x,
  input io_ptw_pmp_5_cfg_w,
  input io_ptw_pmp_5_cfg_r,
  input [29:0] io_ptw_pmp_5_addr,
  input [31:0] io_ptw_pmp_5_mask,
  input io_ptw_pmp_6_cfg_l,
  input [1:0] io_ptw_pmp_6_cfg_a,
  input io_ptw_pmp_6_cfg_x,
  input io_ptw_pmp_6_cfg_w,
  input io_ptw_pmp_6_cfg_r,
  input [29:0] io_ptw_pmp_6_addr,
  input [31:0] io_ptw_pmp_6_mask,
  input io_ptw_pmp_7_cfg_l,
  input [1:0] io_ptw_pmp_7_cfg_a,
  input io_ptw_pmp_7_cfg_x,
  input io_ptw_pmp_7_cfg_w,
  input io_ptw_pmp_7_cfg_r,
  input [29:0] io_ptw_pmp_7_addr,
  input [31:0] io_ptw_pmp_7_mask,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input data_halt,
  input tlb_halt,
  input pma_checker_halt,
  input lfsr_prng_halt) ; 
   wire tlb_clock ;  
   wire tlb_reset ;  
   wire tlb_io_req_ready ;  
   wire tlb_io_req_valid ;  
   wire [39:0] tlb_io_req_bits_vaddr ;  
   wire tlb_io_req_bits_passthrough ;  
   wire [1:0] tlb_io_req_bits_size ;  
   wire [4:0] tlb_io_req_bits_cmd ;  
   wire tlb_io_resp_miss ;  
   wire [31:0] tlb_io_resp_paddr ;  
   wire tlb_io_resp_pf_ld ;  
   wire tlb_io_resp_pf_st ;  
   wire tlb_io_resp_ae_ld ;  
   wire tlb_io_resp_ae_st ;  
   wire tlb_io_resp_ma_ld ;  
   wire tlb_io_resp_ma_st ;  
   wire tlb_io_resp_cacheable ;  
   wire tlb_io_sfence_valid ;  
   wire tlb_io_sfence_bits_rs1 ;  
   wire tlb_io_sfence_bits_rs2 ;  
   wire [38:0] tlb_io_sfence_bits_addr ;  
   wire tlb_io_ptw_req_ready ;  
   wire tlb_io_ptw_req_valid ;  
   wire [26:0] tlb_io_ptw_req_bits_bits_addr ;  
   wire tlb_io_ptw_resp_valid ;  
   wire tlb_io_ptw_resp_bits_ae ;  
   wire [53:0] tlb_io_ptw_resp_bits_pte_ppn ;  
   wire tlb_io_ptw_resp_bits_pte_d ;  
   wire tlb_io_ptw_resp_bits_pte_a ;  
   wire tlb_io_ptw_resp_bits_pte_g ;  
   wire tlb_io_ptw_resp_bits_pte_u ;  
   wire tlb_io_ptw_resp_bits_pte_x ;  
   wire tlb_io_ptw_resp_bits_pte_w ;  
   wire tlb_io_ptw_resp_bits_pte_r ;  
   wire tlb_io_ptw_resp_bits_pte_v ;  
   wire [1:0] tlb_io_ptw_resp_bits_level ;  
   wire tlb_io_ptw_resp_bits_homogeneous ;  
   wire [3:0] tlb_io_ptw_ptbr_mode ;  
   wire tlb_io_ptw_status_debug ;  
   wire [1:0] tlb_io_ptw_status_dprv ;  
   wire tlb_io_ptw_status_mxr ;  
   wire tlb_io_ptw_status_sum ;  
   wire tlb_io_ptw_pmp_0_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_0_cfg_a ;  
   wire tlb_io_ptw_pmp_0_cfg_x ;  
   wire tlb_io_ptw_pmp_0_cfg_w ;  
   wire tlb_io_ptw_pmp_0_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_0_addr ;  
   wire [31:0] tlb_io_ptw_pmp_0_mask ;  
   wire tlb_io_ptw_pmp_1_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_1_cfg_a ;  
   wire tlb_io_ptw_pmp_1_cfg_x ;  
   wire tlb_io_ptw_pmp_1_cfg_w ;  
   wire tlb_io_ptw_pmp_1_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_1_addr ;  
   wire [31:0] tlb_io_ptw_pmp_1_mask ;  
   wire tlb_io_ptw_pmp_2_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_2_cfg_a ;  
   wire tlb_io_ptw_pmp_2_cfg_x ;  
   wire tlb_io_ptw_pmp_2_cfg_w ;  
   wire tlb_io_ptw_pmp_2_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_2_addr ;  
   wire [31:0] tlb_io_ptw_pmp_2_mask ;  
   wire tlb_io_ptw_pmp_3_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_3_cfg_a ;  
   wire tlb_io_ptw_pmp_3_cfg_x ;  
   wire tlb_io_ptw_pmp_3_cfg_w ;  
   wire tlb_io_ptw_pmp_3_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_3_addr ;  
   wire [31:0] tlb_io_ptw_pmp_3_mask ;  
   wire tlb_io_ptw_pmp_4_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_4_cfg_a ;  
   wire tlb_io_ptw_pmp_4_cfg_x ;  
   wire tlb_io_ptw_pmp_4_cfg_w ;  
   wire tlb_io_ptw_pmp_4_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_4_addr ;  
   wire [31:0] tlb_io_ptw_pmp_4_mask ;  
   wire tlb_io_ptw_pmp_5_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_5_cfg_a ;  
   wire tlb_io_ptw_pmp_5_cfg_x ;  
   wire tlb_io_ptw_pmp_5_cfg_w ;  
   wire tlb_io_ptw_pmp_5_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_5_addr ;  
   wire [31:0] tlb_io_ptw_pmp_5_mask ;  
   wire tlb_io_ptw_pmp_6_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_6_cfg_a ;  
   wire tlb_io_ptw_pmp_6_cfg_x ;  
   wire tlb_io_ptw_pmp_6_cfg_w ;  
   wire tlb_io_ptw_pmp_6_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_6_addr ;  
   wire [31:0] tlb_io_ptw_pmp_6_mask ;  
   wire tlb_io_ptw_pmp_7_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_7_cfg_a ;  
   wire tlb_io_ptw_pmp_7_cfg_x ;  
   wire tlb_io_ptw_pmp_7_cfg_w ;  
   wire tlb_io_ptw_pmp_7_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_7_addr ;  
   wire [31:0] tlb_io_ptw_pmp_7_mask ;  
   wire [29:0] tlb_io_covSum ;  
   wire tlb_metaAssert ;  
   wire tlb_metaReset ;  
   wire pma_checker_clock ;  
   wire pma_checker_reset ;  
   wire pma_checker_io_req_ready ;  
   wire pma_checker_io_req_valid ;  
   wire [39:0] pma_checker_io_req_bits_vaddr ;  
   wire pma_checker_io_req_bits_passthrough ;  
   wire [1:0] pma_checker_io_req_bits_size ;  
   wire [4:0] pma_checker_io_req_bits_cmd ;  
   wire pma_checker_io_resp_miss ;  
   wire [31:0] pma_checker_io_resp_paddr ;  
   wire pma_checker_io_resp_pf_ld ;  
   wire pma_checker_io_resp_pf_st ;  
   wire pma_checker_io_resp_ae_ld ;  
   wire pma_checker_io_resp_ae_st ;  
   wire pma_checker_io_resp_ma_ld ;  
   wire pma_checker_io_resp_ma_st ;  
   wire pma_checker_io_resp_cacheable ;  
   wire pma_checker_io_sfence_valid ;  
   wire pma_checker_io_sfence_bits_rs1 ;  
   wire pma_checker_io_sfence_bits_rs2 ;  
   wire [38:0] pma_checker_io_sfence_bits_addr ;  
   wire pma_checker_io_ptw_req_ready ;  
   wire pma_checker_io_ptw_req_valid ;  
   wire [26:0] pma_checker_io_ptw_req_bits_bits_addr ;  
   wire pma_checker_io_ptw_resp_valid ;  
   wire pma_checker_io_ptw_resp_bits_ae ;  
   wire [53:0] pma_checker_io_ptw_resp_bits_pte_ppn ;  
   wire pma_checker_io_ptw_resp_bits_pte_d ;  
   wire pma_checker_io_ptw_resp_bits_pte_a ;  
   wire pma_checker_io_ptw_resp_bits_pte_g ;  
   wire pma_checker_io_ptw_resp_bits_pte_u ;  
   wire pma_checker_io_ptw_resp_bits_pte_x ;  
   wire pma_checker_io_ptw_resp_bits_pte_w ;  
   wire pma_checker_io_ptw_resp_bits_pte_r ;  
   wire pma_checker_io_ptw_resp_bits_pte_v ;  
   wire [1:0] pma_checker_io_ptw_resp_bits_level ;  
   wire pma_checker_io_ptw_resp_bits_homogeneous ;  
   wire [3:0] pma_checker_io_ptw_ptbr_mode ;  
   wire pma_checker_io_ptw_status_debug ;  
   wire [1:0] pma_checker_io_ptw_status_dprv ;  
   wire pma_checker_io_ptw_status_mxr ;  
   wire pma_checker_io_ptw_status_sum ;  
   wire pma_checker_io_ptw_pmp_0_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_0_cfg_a ;  
   wire pma_checker_io_ptw_pmp_0_cfg_x ;  
   wire pma_checker_io_ptw_pmp_0_cfg_w ;  
   wire pma_checker_io_ptw_pmp_0_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_0_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_0_mask ;  
   wire pma_checker_io_ptw_pmp_1_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_1_cfg_a ;  
   wire pma_checker_io_ptw_pmp_1_cfg_x ;  
   wire pma_checker_io_ptw_pmp_1_cfg_w ;  
   wire pma_checker_io_ptw_pmp_1_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_1_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_1_mask ;  
   wire pma_checker_io_ptw_pmp_2_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_2_cfg_a ;  
   wire pma_checker_io_ptw_pmp_2_cfg_x ;  
   wire pma_checker_io_ptw_pmp_2_cfg_w ;  
   wire pma_checker_io_ptw_pmp_2_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_2_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_2_mask ;  
   wire pma_checker_io_ptw_pmp_3_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_3_cfg_a ;  
   wire pma_checker_io_ptw_pmp_3_cfg_x ;  
   wire pma_checker_io_ptw_pmp_3_cfg_w ;  
   wire pma_checker_io_ptw_pmp_3_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_3_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_3_mask ;  
   wire pma_checker_io_ptw_pmp_4_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_4_cfg_a ;  
   wire pma_checker_io_ptw_pmp_4_cfg_x ;  
   wire pma_checker_io_ptw_pmp_4_cfg_w ;  
   wire pma_checker_io_ptw_pmp_4_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_4_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_4_mask ;  
   wire pma_checker_io_ptw_pmp_5_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_5_cfg_a ;  
   wire pma_checker_io_ptw_pmp_5_cfg_x ;  
   wire pma_checker_io_ptw_pmp_5_cfg_w ;  
   wire pma_checker_io_ptw_pmp_5_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_5_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_5_mask ;  
   wire pma_checker_io_ptw_pmp_6_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_6_cfg_a ;  
   wire pma_checker_io_ptw_pmp_6_cfg_x ;  
   wire pma_checker_io_ptw_pmp_6_cfg_w ;  
   wire pma_checker_io_ptw_pmp_6_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_6_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_6_mask ;  
   wire pma_checker_io_ptw_pmp_7_cfg_l ;  
   wire [1:0] pma_checker_io_ptw_pmp_7_cfg_a ;  
   wire pma_checker_io_ptw_pmp_7_cfg_x ;  
   wire pma_checker_io_ptw_pmp_7_cfg_w ;  
   wire pma_checker_io_ptw_pmp_7_cfg_r ;  
   wire [29:0] pma_checker_io_ptw_pmp_7_addr ;  
   wire [31:0] pma_checker_io_ptw_pmp_7_mask ;  
   wire [29:0] pma_checker_io_covSum ;  
   wire pma_checker_metaAssert ;  
   wire pma_checker_metaReset ;  
   wire lfsr_prng_clock ;  
   wire lfsr_prng_reset ;  
   wire lfsr_prng_io_increment ;  
   wire lfsr_prng_io_out_0 ;  
   wire lfsr_prng_io_out_1 ;  
   wire lfsr_prng_io_out_2 ;  
   wire lfsr_prng_io_out_3 ;  
   wire lfsr_prng_io_out_4 ;  
   wire lfsr_prng_io_out_5 ;  
   wire lfsr_prng_io_out_6 ;  
   wire lfsr_prng_io_out_7 ;  
   wire lfsr_prng_io_out_8 ;  
   wire lfsr_prng_io_out_9 ;  
   wire lfsr_prng_io_out_10 ;  
   wire lfsr_prng_io_out_11 ;  
   wire lfsr_prng_io_out_12 ;  
   wire lfsr_prng_io_out_13 ;  
   wire lfsr_prng_io_out_14 ;  
   wire lfsr_prng_io_out_15 ;  
   wire [29:0] lfsr_prng_io_covSum ;  
   wire lfsr_prng_metaAssert ;  
   wire lfsr_prng_metaReset ;  
   wire metaArb_io_in_0_valid ;  
   wire [39:0] metaArb_io_in_0_bits_addr ;  
   wire [5:0] metaArb_io_in_0_bits_idx ;  
   wire metaArb_io_in_1_valid ;  
   wire [39:0] metaArb_io_in_1_bits_addr ;  
   wire [5:0] metaArb_io_in_1_bits_idx ;  
   wire [21:0] metaArb_io_in_1_bits_data ;  
   wire metaArb_io_in_2_valid ;  
   wire [39:0] metaArb_io_in_2_bits_addr ;  
   wire [5:0] metaArb_io_in_2_bits_idx ;  
   wire [3:0] metaArb_io_in_2_bits_way_en ;  
   wire [21:0] metaArb_io_in_2_bits_data ;  
   wire metaArb_io_in_3_valid ;  
   wire [39:0] metaArb_io_in_3_bits_addr ;  
   wire [5:0] metaArb_io_in_3_bits_idx ;  
   wire [3:0] metaArb_io_in_3_bits_way_en ;  
   wire [21:0] metaArb_io_in_3_bits_data ;  
   wire metaArb_io_in_4_ready ;  
   wire metaArb_io_in_4_valid ;  
   wire [39:0] metaArb_io_in_4_bits_addr ;  
   wire [5:0] metaArb_io_in_4_bits_idx ;  
   wire [3:0] metaArb_io_in_4_bits_way_en ;  
   wire [21:0] metaArb_io_in_4_bits_data ;  
   wire metaArb_io_in_5_ready ;  
   wire metaArb_io_in_5_valid ;  
   wire [39:0] metaArb_io_in_5_bits_addr ;  
   wire [5:0] metaArb_io_in_5_bits_idx ;  
   wire metaArb_io_in_6_ready ;  
   wire metaArb_io_in_6_valid ;  
   wire [39:0] metaArb_io_in_6_bits_addr ;  
   wire [5:0] metaArb_io_in_6_bits_idx ;  
   wire [3:0] metaArb_io_in_6_bits_way_en ;  
   wire [21:0] metaArb_io_in_6_bits_data ;  
   wire metaArb_io_in_7_ready ;  
   wire metaArb_io_in_7_valid ;  
   wire [39:0] metaArb_io_in_7_bits_addr ;  
   wire [5:0] metaArb_io_in_7_bits_idx ;  
   wire [3:0] metaArb_io_in_7_bits_way_en ;  
   wire [21:0] metaArb_io_in_7_bits_data ;  
   wire metaArb_io_out_valid ;  
   wire metaArb_io_out_bits_write ;  
   wire [39:0] metaArb_io_out_bits_addr ;  
   wire [5:0] metaArb_io_out_bits_idx ;  
   wire [3:0] metaArb_io_out_bits_way_en ;  
   wire [21:0] metaArb_io_out_bits_data ;  
   wire [29:0] metaArb_io_covSum ;  
   wire metaArb_metaAssert ;  
   reg [21:0] tag_array_0[0:63] ;  
   reg [31:0] _RAND_0 ;  
   wire [21:0] tag_array_0_s1_meta_data ;  
   wire [5:0] tag_array_0_s1_meta_addr ;  
   wire [21:0] tag_array_0_MPORT_data ;  
   wire [5:0] tag_array_0_MPORT_addr ;  
   wire tag_array_0_MPORT_mask ;  
   wire tag_array_0_MPORT_en ;  
   reg tag_array_0_s1_meta_en_pipe_0 ;  
   reg [31:0] _RAND_1 ;  
   reg [5:0] tag_array_0_s1_meta_addr_pipe_0 ;  
   reg [31:0] _RAND_2 ;  
   reg [21:0] tag_array_1[0:63] ;  
   reg [31:0] _RAND_3 ;  
   wire [21:0] tag_array_1_s1_meta_data ;  
   wire [5:0] tag_array_1_s1_meta_addr ;  
   wire [21:0] tag_array_1_MPORT_data ;  
   wire [5:0] tag_array_1_MPORT_addr ;  
   wire tag_array_1_MPORT_mask ;  
   wire tag_array_1_MPORT_en ;  
   reg tag_array_1_s1_meta_en_pipe_0 ;  
   reg [31:0] _RAND_4 ;  
   reg [5:0] tag_array_1_s1_meta_addr_pipe_0 ;  
   reg [31:0] _RAND_5 ;  
   reg [21:0] tag_array_2[0:63] ;  
   reg [31:0] _RAND_6 ;  
   wire [21:0] tag_array_2_s1_meta_data ;  
   wire [5:0] tag_array_2_s1_meta_addr ;  
   wire [21:0] tag_array_2_MPORT_data ;  
   wire [5:0] tag_array_2_MPORT_addr ;  
   wire tag_array_2_MPORT_mask ;  
   wire tag_array_2_MPORT_en ;  
   reg tag_array_2_s1_meta_en_pipe_0 ;  
   reg [31:0] _RAND_7 ;  
   reg [5:0] tag_array_2_s1_meta_addr_pipe_0 ;  
   reg [31:0] _RAND_8 ;  
   reg [21:0] tag_array_3[0:63] ;  
   reg [31:0] _RAND_9 ;  
   wire [21:0] tag_array_3_s1_meta_data ;  
   wire [5:0] tag_array_3_s1_meta_addr ;  
   wire [21:0] tag_array_3_MPORT_data ;  
   wire [5:0] tag_array_3_MPORT_addr ;  
   wire tag_array_3_MPORT_mask ;  
   wire tag_array_3_MPORT_en ;  
   reg tag_array_3_s1_meta_en_pipe_0 ;  
   reg [31:0] _RAND_10 ;  
   reg [5:0] tag_array_3_s1_meta_addr_pipe_0 ;  
   reg [31:0] _RAND_11 ;  
   wire data_clock ;  
   wire data_io_req_valid ;  
   wire [11:0] data_io_req_bits_addr ;  
   wire data_io_req_bits_write ;  
   wire [63:0] data_io_req_bits_wdata ;  
   wire [7:0] data_io_req_bits_eccMask ;  
   wire [3:0] data_io_req_bits_way_en ;  
   wire [63:0] data_io_resp_0 ;  
   wire [63:0] data_io_resp_1 ;  
   wire [63:0] data_io_resp_2 ;  
   wire [63:0] data_io_resp_3 ;  
   wire [29:0] data_io_covSum ;  
   wire data_metaAssert ;  
   wire data_metaReset ;  
   wire dataArb_io_in_0_valid ;  
   wire [11:0] dataArb_io_in_0_bits_addr ;  
   wire dataArb_io_in_0_bits_write ;  
   wire [63:0] dataArb_io_in_0_bits_wdata ;  
   wire [7:0] dataArb_io_in_0_bits_eccMask ;  
   wire [3:0] dataArb_io_in_0_bits_way_en ;  
   wire dataArb_io_in_1_ready ;  
   wire dataArb_io_in_1_valid ;  
   wire [11:0] dataArb_io_in_1_bits_addr ;  
   wire dataArb_io_in_1_bits_write ;  
   wire [63:0] dataArb_io_in_1_bits_wdata ;  
   wire [3:0] dataArb_io_in_1_bits_way_en ;  
   wire dataArb_io_in_2_ready ;  
   wire dataArb_io_in_2_valid ;  
   wire [11:0] dataArb_io_in_2_bits_addr ;  
   wire [63:0] dataArb_io_in_2_bits_wdata ;  
   wire dataArb_io_in_3_ready ;  
   wire dataArb_io_in_3_valid ;  
   wire [11:0] dataArb_io_in_3_bits_addr ;  
   wire [63:0] dataArb_io_in_3_bits_wdata ;  
   wire dataArb_io_in_3_bits_wordMask ;  
   wire dataArb_io_out_valid ;  
   wire [11:0] dataArb_io_out_bits_addr ;  
   wire dataArb_io_out_bits_write ;  
   wire [63:0] dataArb_io_out_bits_wdata ;  
   wire [7:0] dataArb_io_out_bits_eccMask ;  
   wire [3:0] dataArb_io_out_bits_way_en ;  
   wire [29:0] dataArb_io_covSum ;  
   wire dataArb_metaAssert ;  
   wire [7:0] amoalu_io_mask ;  
   wire [4:0] amoalu_io_cmd ;  
   wire [63:0] amoalu_io_lhs ;  
   wire [63:0] amoalu_io_rhs ;  
   wire [63:0] amoalu_io_out ;  
   wire [29:0] amoalu_io_covSum ;  
   wire amoalu_metaAssert ;  
   wire [7:0] lfsr_lo ;  
   wire [15:0] lfsr ;  
   wire s1_valid_x9 ;  
   reg s1_valid ;  
   reg [31:0] _RAND_12 ;  
   reg [2:0] blockProbeAfterGrantCount ;  
   reg [31:0] _RAND_13 ;  
   wire _block_probe_for_core_progress_T ;  
   reg [6:0] lrscCount ;  
   reg [31:0] _RAND_14 ;  
   wire lrscValid ;  
   wire block_probe_for_core_progress ;  
   reg s1_probe ;  
   reg [31:0] _RAND_15 ;  
   reg s2_probe ;  
   reg [31:0] _RAND_16 ;  
   wire _releaseInFlight_T ;  
   reg [3:0] release_state ;  
   reg [31:0] _RAND_17 ;  
   wire _releaseInFlight_T_1 ;  
   wire releaseInFlight ;  
   reg release_ack_wait ;  
   reg [31:0] _RAND_18 ;  
   reg [31:0] release_ack_addr ;  
   reg [31:0] _RAND_19 ;  
   wire [31:0] _block_probe_for_pending_release_ack_T ;  
   wire _block_probe_for_pending_release_ack_T_2 ;  
   wire block_probe_for_pending_release_ack ;  
   wire _block_probe_for_ordering_T ;  
   reg grantInProgress ;  
   reg [31:0] _RAND_20 ;  
   wire block_probe_for_ordering ;  
   wire _bundleOut_0_b_ready_T ;  
   wire _bundleOut_0_b_ready_T_1 ;  
   reg s2_valid ;  
   reg [31:0] _RAND_21 ;  
   wire _bundleOut_0_b_ready_T_2 ;  
   wire tl_out__b_ready ;  
   wire s1_probe_x12 ;  
   reg [1:0] probe_bits_param ;  
   reg [31:0] _RAND_22 ;  
   reg [3:0] probe_bits_size ;  
   reg [31:0] _RAND_23 ;  
   reg probe_bits_source ;  
   reg [31:0] _RAND_24 ;  
   reg [31:0] probe_bits_address ;  
   reg [31:0] _RAND_25 ;  
   wire s1_valid_masked ;  
   wire s2_meta_error ;  
   reg [1:0] s2_probe_state_state ;  
   reg [31:0] _RAND_26 ;  
   wire [3:0] _T_118 ;  
   wire _T_175 ;  
   wire _T_171 ;  
   wire _T_167 ;  
   wire _T_163 ;  
   wire _T_159 ;  
   wire _T_155 ;  
   wire _T_151 ;  
   wire _T_147 ;  
   wire _T_143 ;  
   wire _T_139 ;  
   wire _T_135 ;  
   wire _T_131 ;  
   wire _T_148 ;  
   wire _T_152 ;  
   wire _T_156 ;  
   wire _T_160 ;  
   wire _T_164 ;  
   wire _T_168 ;  
   wire _T_172 ;  
   wire s2_prb_ack_data ;  
   wire _T_303 ;  
   reg [8:0] counter_1 ;  
   reg [31:0] _RAND_27 ;  
   wire _last_T_2 ;  
   wire _T_308 ;  
   wire _T_309 ;  
   wire _T_311 ;  
   wire _T_310 ;  
   wire _T_312 ;  
   wire [2:0] _GEN_323 ;  
   wire _T_307 ;  
   wire _T_306 ;  
   wire [2:0] _GEN_315 ;  
   wire [2:0] tl_out__c_bits_opcode ;  
   wire beats1_opdata_1 ;  
   wire [3:0] tl_out__c_bits_size ;  
   wire [26:0] _beats1_decode_T_5 ;  
   wire [8:0] beats1_decode_1 ;  
   wire [8:0] beats1_1 ;  
   wire _last_T_3 ;  
   wire c_last ;  
   wire _T_305 ;  
   reg s2_release_data_valid ;  
   reg [31:0] _RAND_28 ;  
   wire c_first ;  
   wire _bundleOut_0_c_valid_T_3 ;  
   wire _bundleOut_0_c_valid_T_5 ;  
   wire _GEN_264 ;  
   wire _GEN_274 ;  
   wire _GEN_285 ;  
   wire _GEN_302 ;  
   wire tl_out__c_valid ;  
   wire _T_297 ;  
   wire releaseDone ;  
   wire _GEN_262 ;  
   wire _GEN_272 ;  
   wire probeNack ;  
   reg [4:0] s1_req_cmd ;  
   reg [31:0] _RAND_29 ;  
   wire _s1_read_T ;  
   wire _s1_read_T_1 ;  
   wire _s1_read_T_2 ;  
   wire _s1_read_T_3 ;  
   wire _s1_read_T_4 ;  
   wire _s1_read_T_5 ;  
   wire _s1_read_T_6 ;  
   wire _s1_read_T_9 ;  
   wire _s1_read_T_7 ;  
   wire _s1_read_T_10 ;  
   wire _s1_read_T_8 ;  
   wire _s1_read_T_11 ;  
   wire _s1_read_T_12 ;  
   wire _s1_read_T_13 ;  
   wire _s1_read_T_17 ;  
   wire _s1_read_T_14 ;  
   wire _s1_read_T_18 ;  
   wire _s1_read_T_15 ;  
   wire _s1_read_T_19 ;  
   wire _s1_read_T_16 ;  
   wire _s1_read_T_20 ;  
   wire _s1_read_T_21 ;  
   wire s1_read ;  
   reg [4:0] s2_req_cmd ;  
   reg [31:0] _RAND_30 ;  
   wire _s2_write_T ;  
   wire _s2_write_T_1 ;  
   wire _s2_write_T_2 ;  
   wire _s2_write_T_3 ;  
   wire _s2_write_T_4 ;  
   wire _s2_write_T_5 ;  
   wire _s2_write_T_6 ;  
   wire _s2_write_T_9 ;  
   wire _s2_write_T_7 ;  
   wire _s2_write_T_10 ;  
   wire _s2_write_T_8 ;  
   wire _s2_write_T_11 ;  
   wire _s2_write_T_12 ;  
   wire _s2_write_T_13 ;  
   wire _s2_write_T_17 ;  
   wire _s2_write_T_14 ;  
   wire _s2_write_T_18 ;  
   wire _s2_write_T_15 ;  
   wire _s2_write_T_19 ;  
   wire _s2_write_T_16 ;  
   wire _s2_write_T_20 ;  
   wire _s2_write_T_21 ;  
   wire s2_write ;  
   wire _pstore1_valid_likely_T ;  
   reg pstore1_held ;  
   reg [31:0] _RAND_31 ;  
   wire pstore1_valid_likely ;  
   reg [39:0] pstore1_addr ;  
   reg [63:0] _RAND_32 ;  
   reg [39:0] s1_req_addr ;  
   reg [63:0] _RAND_33 ;  
   wire [27:0] s1_vaddr_hi ;  
   wire [11:0] s1_vaddr_lo ;  
   wire [39:0] s1_vaddr ;  
   wire _s1_hazard_T_2 ;  
   wire _s1_write_T ;  
   wire _s1_write_T_1 ;  
   wire _s1_write_T_2 ;  
   wire _s1_write_T_4 ;  
   wire s1_write ;  
   reg [7:0] pstore1_mask ;  
   reg [31:0] _RAND_34 ;  
   wire s1_hazard_hi_hi_hi ;  
   wire s1_hazard_hi_hi_lo ;  
   wire s1_hazard_hi_lo_hi ;  
   wire s1_hazard_hi_lo_lo ;  
   wire s1_hazard_lo_hi_hi ;  
   wire s1_hazard_lo_hi_lo ;  
   wire s1_hazard_lo_lo_hi ;  
   wire s1_hazard_lo_lo_lo ;  
   wire [7:0] _s1_hazard_T_11 ;  
   wire s1_hazard_hi_hi_hi_1 ;  
   wire s1_hazard_hi_hi_lo_1 ;  
   wire s1_hazard_hi_lo_hi_1 ;  
   wire s1_hazard_hi_lo_lo_1 ;  
   wire s1_hazard_lo_hi_hi_1 ;  
   wire s1_hazard_lo_hi_lo_1 ;  
   wire s1_hazard_lo_lo_hi_1 ;  
   wire s1_hazard_lo_lo_lo_1 ;  
   wire [7:0] _s1_hazard_T_12 ;  
   reg [1:0] s1_req_size ;  
   reg [31:0] _RAND_35 ;  
   wire _s1_mask_xwr_upper_T_2 ;  
   wire s1_mask_xwr_hi ;  
   wire s1_mask_xwr_lo ;  
   wire [1:0] _s1_mask_xwr_T ;  
   wire [1:0] _s1_mask_xwr_upper_T_5 ;  
   wire _s1_mask_xwr_upper_T_6 ;  
   wire [1:0] _s1_mask_xwr_upper_T_7 ;  
   wire [1:0] s1_mask_xwr_hi_1 ;  
   wire [1:0] s1_mask_xwr_lo_1 ;  
   wire [3:0] _s1_mask_xwr_T_1 ;  
   wire [3:0] _s1_mask_xwr_upper_T_9 ;  
   wire _s1_mask_xwr_upper_T_10 ;  
   wire [3:0] _s1_mask_xwr_upper_T_11 ;  
   wire [3:0] s1_mask_xwr_hi_2 ;  
   wire [3:0] s1_mask_xwr_lo_2 ;  
   wire [7:0] s1_mask_xwr ;  
   wire s1_hazard_hi_hi_hi_2 ;  
   wire s1_hazard_hi_hi_lo_2 ;  
   wire s1_hazard_hi_lo_hi_2 ;  
   wire s1_hazard_hi_lo_lo_2 ;  
   wire s1_hazard_lo_hi_hi_2 ;  
   wire s1_hazard_lo_hi_lo_2 ;  
   wire s1_hazard_lo_lo_hi_2 ;  
   wire s1_hazard_lo_lo_lo_2 ;  
   wire [7:0] _s1_hazard_T_21 ;  
   wire s1_hazard_hi_hi_hi_3 ;  
   wire s1_hazard_hi_hi_lo_3 ;  
   wire s1_hazard_hi_lo_hi_3 ;  
   wire s1_hazard_hi_lo_lo_3 ;  
   wire s1_hazard_lo_hi_hi_3 ;  
   wire s1_hazard_lo_hi_lo_3 ;  
   wire s1_hazard_lo_lo_hi_3 ;  
   wire s1_hazard_lo_lo_lo_3 ;  
   wire [7:0] _s1_hazard_T_22 ;  
   wire [7:0] _s1_hazard_T_23 ;  
   wire _s1_hazard_T_24 ;  
   wire [7:0] _s1_hazard_T_25 ;  
   wire _s1_hazard_T_26 ;  
   wire _s1_hazard_T_27 ;  
   wire _s1_hazard_T_28 ;  
   wire _s1_hazard_T_29 ;  
   reg pstore2_valid ;  
   reg [31:0] _RAND_36 ;  
   reg [39:0] pstore2_addr ;  
   reg [63:0] _RAND_37 ;  
   wire _s1_hazard_T_32 ;  
   reg [7:0] mask ;  
   reg [31:0] _RAND_38 ;  
   wire s1_hazard_hi_hi_hi_4 ;  
   wire s1_hazard_hi_hi_lo_4 ;  
   wire s1_hazard_hi_lo_hi_4 ;  
   wire s1_hazard_hi_lo_lo_4 ;  
   wire s1_hazard_lo_hi_hi_4 ;  
   wire s1_hazard_lo_hi_lo_4 ;  
   wire s1_hazard_lo_lo_hi_4 ;  
   wire s1_hazard_lo_lo_lo_4 ;  
   wire [7:0] _s1_hazard_T_41 ;  
   wire s1_hazard_hi_hi_hi_5 ;  
   wire s1_hazard_hi_hi_lo_5 ;  
   wire s1_hazard_hi_lo_hi_5 ;  
   wire s1_hazard_hi_lo_lo_5 ;  
   wire s1_hazard_lo_hi_hi_5 ;  
   wire s1_hazard_lo_hi_lo_5 ;  
   wire s1_hazard_lo_lo_hi_5 ;  
   wire s1_hazard_lo_lo_lo_5 ;  
   wire [7:0] _s1_hazard_T_42 ;  
   wire [7:0] _s1_hazard_T_53 ;  
   wire _s1_hazard_T_54 ;  
   wire [7:0] _s1_hazard_T_55 ;  
   wire _s1_hazard_T_56 ;  
   wire _s1_hazard_T_57 ;  
   wire _s1_hazard_T_58 ;  
   wire _s1_hazard_T_59 ;  
   wire s1_hazard ;  
   wire s1_raw_hazard ;  
   wire _T_262 ;  
   wire [5:0] _s2_valid_no_xcpt_T ;  
   wire _s2_valid_no_xcpt_T_1 ;  
   wire s2_valid_no_xcpt ;  
   reg s2_not_nacked_in_s1 ;  
   reg [31:0] _RAND_39 ;  
   wire s2_valid_masked ;  
   wire _s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1 ;  
   wire _c_cat_T_45 ;  
   wire _c_cat_T_46 ;  
   wire _c_cat_T_47 ;  
   wire c_cat_lo ;  
   reg [1:0] s2_hit_state_state ;  
   reg [31:0] _RAND_40 ;  
   wire [3:0] _T_71 ;  
   wire _T_117 ;  
   wire _T_114 ;  
   wire _T_111 ;  
   wire _T_108 ;  
   wire _T_105 ;  
   wire _T_102 ;  
   wire _T_99 ;  
   wire _T_96 ;  
   wire _T_93 ;  
   wire _T_90 ;  
   wire _T_87 ;  
   wire _T_84 ;  
   wire _T_103 ;  
   wire _T_106 ;  
   wire _T_109 ;  
   wire _T_112 ;  
   wire _T_115 ;  
   wire s2_hit ;  
   wire s2_valid_hit_maybe_flush_pre_data_ecc_and_waw ;  
   wire _s2_read_T ;  
   wire _s2_read_T_2 ;  
   wire _s2_read_T_4 ;  
   wire s2_read ;  
   wire s2_readwrite ;  
   wire s2_valid_hit_pre_data_ecc_and_waw ;  
   wire [1:0] _T_86 ;  
   wire [1:0] _T_89 ;  
   wire [1:0] _T_92 ;  
   wire [1:0] _T_95 ;  
   wire [1:0] _T_98 ;  
   wire [1:0] _T_101 ;  
   wire [1:0] _T_104 ;  
   wire [1:0] _T_107 ;  
   wire [1:0] _T_110 ;  
   wire [1:0] _T_113 ;  
   wire [1:0] _T_116 ;  
   wire [1:0] s2_grow_param ;  
   wire _s2_update_meta_T ;  
   wire s2_update_meta ;  
   wire _T_241 ;  
   wire _T_242 ;  
   wire s1_readwrite ;  
   wire _s1_flush_line_T ;  
   wire s1_flush_line ;  
   wire _s1_cmd_uses_tlb_T ;  
   wire _s1_cmd_uses_tlb_T_1 ;  
   wire s1_cmd_uses_tlb ;  
   wire _T_13 ;  
   wire _T_14 ;  
   wire _GEN_117 ;  
   wire _GEN_141 ;  
   wire _GEN_283 ;  
   wire s1_nack ;  
   wire s1_valid_not_nacked ;  
   wire s0_clk_en ;  
   wire [33:0] s0_req_addr_hi ;  
   wire [5:0] s0_req_addr_lo ;  
   wire [39:0] s0_req_addr ;  
   wire s0_req_phys ;  
   reg [6:0] s1_req_tag ;  
   reg [31:0] _RAND_41 ;  
   reg s1_req_signed ;  
   reg [31:0] _RAND_42 ;  
   reg [39:0] s1_tlb_req_vaddr ;  
   reg [63:0] _RAND_43 ;  
   reg s1_tlb_req_passthrough ;  
   reg [31:0] _RAND_44 ;  
   reg [1:0] s1_tlb_req_size ;  
   reg [31:0] _RAND_45 ;  
   reg [4:0] s1_tlb_req_cmd ;  
   reg [31:0] _RAND_46 ;  
   wire s1_sfence ;  
   reg s1_flush_valid ;  
   reg [31:0] _RAND_47 ;  
   reg cached_grant_wait ;  
   reg [31:0] _RAND_48 ;  
   reg resetting ;  
   reg [31:0] _RAND_49 ;  
   reg [7:0] flushCounter ;  
   reg [31:0] _RAND_50 ;  
   reg [3:0] refill_way ;  
   reg [31:0] _RAND_51 ;  
   wire inWriteback ;  
   wire _io_cpu_req_ready_T ;  
   wire _io_cpu_req_ready_T_2 ;  
   wire _io_cpu_req_ready_T_4 ;  
   reg uncachedInFlight_0 ;  
   reg [31:0] _RAND_52 ;  
   reg [39:0] uncachedReqs_0_addr ;  
   reg [63:0] _RAND_53 ;  
   reg [6:0] uncachedReqs_0_tag ;  
   reg [31:0] _RAND_54 ;  
   reg [1:0] uncachedReqs_0_size ;  
   reg [31:0] _RAND_55 ;  
   reg uncachedReqs_0_signed ;  
   reg [31:0] _RAND_56 ;  
   wire _s0_read_T ;  
   wire _s0_read_T_1 ;  
   wire _s0_read_T_2 ;  
   wire _s0_read_T_3 ;  
   wire _s0_read_T_4 ;  
   wire _s0_read_T_5 ;  
   wire _s0_read_T_6 ;  
   wire _s0_read_T_7 ;  
   wire _s0_read_T_8 ;  
   wire _s0_read_T_9 ;  
   wire _s0_read_T_10 ;  
   wire _s0_read_T_11 ;  
   wire _s0_read_T_12 ;  
   wire _s0_read_T_13 ;  
   wire _s0_read_T_14 ;  
   wire _s0_read_T_15 ;  
   wire _s0_read_T_16 ;  
   wire _s0_read_T_17 ;  
   wire _s0_read_T_18 ;  
   wire _s0_read_T_19 ;  
   wire _s0_read_T_20 ;  
   wire _s0_read_T_21 ;  
   wire s0_read ;  
   wire _dataArb_io_in_3_valid_res_T ;  
   wire _dataArb_io_in_3_valid_res_T_1 ;  
   wire _dataArb_io_in_3_valid_res_T_2 ;  
   wire res ;  
   wire _dataArb_io_in_3_valid_T_24 ;  
   wire _dataArb_io_in_3_valid_T_25 ;  
   wire _dataArb_io_in_3_valid_T_27 ;  
   wire _dataArb_io_in_3_valid_T_45 ;  
   wire _dataArb_io_in_3_valid_T_49 ;  
   wire _dataArb_io_in_3_valid_T_50 ;  
   wire _dataArb_io_in_3_valid_T_52 ;  
   wire _dataArb_io_in_3_valid_T_54 ;  
   wire _dataArb_io_in_3_valid_T_56 ;  
   wire [27:0] dataArb_io_in_3_bits_addr_hi ;  
   wire [11:0] dataArb_io_in_3_bits_addr_lo ;  
   wire [39:0] _dataArb_io_in_3_bits_addr_T ;  
   wire _T_4 ;  
   wire _GEN_28 ;  
   wire _s1_did_read_T_51 ;  
   wire _s1_did_read_T_52 ;  
   reg s1_did_read ;  
   reg [31:0] _RAND_57 ;  
   reg s1_read_mask ;  
   reg [31:0] _RAND_58 ;  
   wire _GEN_31 ;  
   wire _T_8 ;  
   wire _T_10 ;  
   wire _GEN_32 ;  
   wire [19:0] s1_paddr_hi ;  
   wire [31:0] s1_paddr ;  
   wire [21:0] _WIRE_2 ;  
   wire [19:0] s1_meta_uncorrected_0_tag ;  
   wire [1:0] s1_meta_uncorrected_0_coh_state ;  
   wire [21:0] _WIRE_3 ;  
   wire [19:0] s1_meta_uncorrected_1_tag ;  
   wire [1:0] s1_meta_uncorrected_1_coh_state ;  
   wire [21:0] _WIRE_4 ;  
   wire [19:0] s1_meta_uncorrected_2_tag ;  
   wire [1:0] s1_meta_uncorrected_2_coh_state ;  
   wire [21:0] _WIRE_5 ;  
   wire [19:0] s1_meta_uncorrected_3_tag ;  
   wire [1:0] s1_meta_uncorrected_3_coh_state ;  
   wire [19:0] s1_tag ;  
   wire _T_32 ;  
   wire _T_33 ;  
   wire lo_lo ;  
   wire _T_34 ;  
   wire _T_35 ;  
   wire lo_hi ;  
   wire _T_36 ;  
   wire _T_37 ;  
   wire hi_lo ;  
   wire _T_38 ;  
   wire _T_39 ;  
   wire hi_hi ;  
   wire [3:0] s1_meta_hit_way ;  
   wire _T_42 ;  
   wire [1:0] _T_43 ;  
   wire _T_46 ;  
   wire [1:0] _T_47 ;  
   wire _T_50 ;  
   wire [1:0] _T_51 ;  
   wire _T_54 ;  
   wire [1:0] _T_55 ;  
   wire [1:0] _T_56 ;  
   wire [1:0] _T_57 ;  
   wire [1:0] s1_meta_hit_state_state ;  
   wire s2_hit_valid ;  
   reg [3:0] s2_hit_way ;  
   reg [31:0] _RAND_59 ;  
   reg [1:0] s2_victim_way_r ;  
   reg [31:0] _RAND_60 ;  
   wire [3:0] s2_victim_way ;  
   wire [3:0] s2_victim_or_hit_way ;  
   reg [3:0] s2_probe_way ;  
   reg [31:0] _RAND_61 ;  
   wire [3:0] releaseWay ;  
   wire [3:0] s1_data_way_x35 ;  
   wire [7:0] tl_d_data_encoded_lo_lo_lo ;  
   wire [7:0] tl_d_data_encoded_lo_lo_hi ;  
   wire [7:0] tl_d_data_encoded_lo_hi_lo ;  
   wire [7:0] tl_d_data_encoded_lo_hi_hi ;  
   wire [7:0] tl_d_data_encoded_hi_lo_lo ;  
   wire [7:0] tl_d_data_encoded_hi_lo_hi ;  
   wire [7:0] tl_d_data_encoded_hi_hi_lo ;  
   wire [7:0] tl_d_data_encoded_hi_hi_hi ;  
   wire [31:0] tl_d_data_encoded_lo ;  
   wire [31:0] tl_d_data_encoded_hi ;  
   wire [63:0] _tl_d_data_encoded_T ;  
   wire _T_61 ;  
   wire _T_65 ;  
   wire _T_66 ;  
   wire _T_68 ;  
   wire s2_valid_x37 ;  
   reg [39:0] s2_req_addr ;  
   reg [63:0] _RAND_62 ;  
   reg [6:0] s2_req_tag ;  
   reg [31:0] _RAND_63 ;  
   reg [1:0] s2_req_size ;  
   reg [31:0] _RAND_64 ;  
   reg s2_req_signed ;  
   reg [31:0] _RAND_65 ;  
   wire _s2_cmd_flush_all_T ;  
   wire s2_cmd_flush_line ;  
   reg s2_tlb_xcpt_pf_ld ;  
   reg [31:0] _RAND_66 ;  
   reg s2_tlb_xcpt_pf_st ;  
   reg [31:0] _RAND_67 ;  
   reg s2_tlb_xcpt_ae_ld ;  
   reg [31:0] _RAND_68 ;  
   reg s2_tlb_xcpt_ae_st ;  
   reg [31:0] _RAND_69 ;  
   reg s2_tlb_xcpt_ma_ld ;  
   reg [31:0] _RAND_70 ;  
   reg s2_tlb_xcpt_ma_st ;  
   reg [31:0] _RAND_71 ;  
   reg s2_pma_cacheable ;  
   reg [31:0] _RAND_72 ;  
   wire _T_70 ;  
   wire _s2_pma_T_cacheable ;  
   reg [39:0] s2_vaddr_r ;  
   reg [63:0] _RAND_73 ;  
   wire [27:0] s2_vaddr_hi ;  
   wire [11:0] s2_vaddr_lo ;  
   wire [39:0] s2_vaddr ;  
   reg s2_flush_valid_pre_tag_ecc ;  
   reg [31:0] _RAND_74 ;  
   wire s1_meta_clk_en ;  
   reg [21:0] s2_meta_corrected_r ;  
   reg [31:0] _RAND_75 ;  
   wire [19:0] s2_meta_corrected_0_tag ;  
   wire [1:0] s2_meta_corrected_0_coh_state ;  
   reg [21:0] s2_meta_corrected_r_1 ;  
   reg [31:0] _RAND_76 ;  
   wire [19:0] s2_meta_corrected_1_tag ;  
   wire [1:0] s2_meta_corrected_1_coh_state ;  
   reg [21:0] s2_meta_corrected_r_2 ;  
   reg [31:0] _RAND_77 ;  
   wire [19:0] s2_meta_corrected_2_tag ;  
   wire [1:0] s2_meta_corrected_2_coh_state ;  
   reg [21:0] s2_meta_corrected_r_3 ;  
   reg [31:0] _RAND_78 ;  
   wire [19:0] s2_meta_corrected_3_tag ;  
   wire [1:0] s2_meta_corrected_3_coh_state ;  
   wire s2_flush_valid ;  
   wire _s2_data_en_T ;  
   wire en ;  
   wire _s2_data_word_en_T ;  
   wire word_en ;  
   wire [63:0] s1_all_data_ways_0 ;  
   wire [63:0] s1_all_data_ways_1 ;  
   wire [63:0] s1_all_data_ways_2 ;  
   wire [63:0] s1_all_data_ways_3 ;  
   wire s1_word_en ;  
   wire grantIsUncachedData ;  
   reg blockUncachedGrant ;  
   reg [31:0] _RAND_79 ;  
   wire _T_293 ;  
   wire _T_294 ;  
   wire grantIsRefill ;  
   wire _T_292 ;  
   wire _grantIsCached_T ;  
   wire grantIsCached ;  
   reg [8:0] counter ;  
   reg [31:0] _RAND_80 ;  
   wire d_first ;  
   wire _bundleOut_0_d_ready_T_1 ;  
   wire canAcceptCachedGrant ;  
   wire _bundleOut_0_d_ready_T_2 ;  
   wire _bundleOut_0_d_ready_T_3 ;  
   wire _GEN_233 ;  
   wire tl_out__d_ready ;  
   wire _T_271 ;  
   wire _T_267 ;  
   wire _T_269 ;  
   wire _T_268 ;  
   wire grantIsUncached ;  
   wire [4:0] _GEN_189 ;  
   wire [4:0] _GEN_198 ;  
   wire [4:0] _GEN_211 ;  
   wire [4:0] s1_data_way ;  
   wire [4:0] _s2_data_T_1 ;  
   wire [63:0] _s2_data_T_7 ;  
   wire [63:0] _s2_data_T_8 ;  
   wire [63:0] _s2_data_T_9 ;  
   wire [63:0] _s2_data_T_10 ;  
   wire [63:0] _s2_data_T_11 ;  
   wire [63:0] _s2_data_T_12 ;  
   wire [63:0] _s2_data_T_13 ;  
   wire [63:0] _s2_data_T_14 ;  
   wire [63:0] _s2_data_T_15 ;  
   reg [63:0] s2_data ;  
   reg [63:0] _RAND_81 ;  
   wire [7:0] s2_data_uncorrected_lo_lo_lo ;  
   wire [7:0] s2_data_uncorrected_lo_lo_hi ;  
   wire [7:0] s2_data_uncorrected_lo_hi_lo ;  
   wire [7:0] s2_data_uncorrected_lo_hi_hi ;  
   wire [7:0] s2_data_uncorrected_hi_lo_lo ;  
   wire [7:0] s2_data_uncorrected_hi_lo_hi ;  
   wire [7:0] s2_data_uncorrected_hi_hi_lo ;  
   wire [7:0] s2_data_uncorrected_hi_hi_hi ;  
   wire [31:0] s2_data_corrected_lo ;  
   wire [31:0] s2_data_corrected_hi ;  
   wire [63:0] s2_data_corrected ;  
   wire s2_valid_flush_line ;  
   wire _s2_valid_miss_T ;  
   wire _s2_valid_miss_T_2 ;  
   wire s2_valid_miss ;  
   wire s2_uncached ;  
   wire _s2_valid_cached_miss_T_1 ;  
   wire _s2_valid_cached_miss_T_2 ;  
   wire s2_valid_cached_miss ;  
   wire _s2_want_victimize_T ;  
   wire s2_want_victimize ;  
   wire _s2_valid_uncached_pending_T ;  
   wire _s2_valid_uncached_pending_T_1 ;  
   wire s2_valid_uncached_pending ;  
   wire [1:0] s1_victim_way ;  
   wire [19:0] _s2_victim_tag_T_6 ;  
   wire [19:0] _s2_victim_tag_T_7 ;  
   wire [19:0] _s2_victim_tag_T_8 ;  
   wire [19:0] _s2_victim_tag_T_9 ;  
   wire [19:0] _s2_victim_tag_T_10 ;  
   wire [19:0] _s2_victim_tag_T_11 ;  
   wire [19:0] _s2_victim_tag_T_12 ;  
   wire [1:0] _s2_victim_tag_T_13 ;  
   wire [1:0] _s2_victim_tag_T_14 ;  
   wire [1:0] _s2_victim_tag_T_15 ;  
   wire [1:0] _s2_victim_tag_T_16 ;  
   wire [1:0] _s2_victim_tag_T_17 ;  
   wire [1:0] _s2_victim_tag_T_18 ;  
   wire [1:0] _s2_victim_tag_T_19 ;  
   wire [19:0] s2_victim_tag ;  
   wire [1:0] s2_victim_state_state ;  
   wire [2:0] _T_133 ;  
   wire [2:0] _T_137 ;  
   wire [2:0] _T_141 ;  
   wire [2:0] _T_145 ;  
   wire [2:0] _T_149 ;  
   wire [2:0] _T_153 ;  
   wire [1:0] _T_154 ;  
   wire [2:0] _T_157 ;  
   wire [1:0] _T_158 ;  
   wire [2:0] _T_161 ;  
   wire [1:0] _T_162 ;  
   wire [2:0] _T_165 ;  
   wire [1:0] _T_166 ;  
   wire [2:0] _T_169 ;  
   wire [1:0] _T_170 ;  
   wire [2:0] _T_173 ;  
   wire [1:0] _T_174 ;  
   wire [2:0] s2_report_param ;  
   wire [1:0] probeNewCoh_state ;  
   wire [3:0] _T_182 ;  
   wire _T_195 ;  
   wire [2:0] _T_197 ;  
   wire _T_199 ;  
   wire [2:0] _T_201 ;  
   wire _T_203 ;  
   wire [2:0] _T_205 ;  
   wire _T_207 ;  
   wire [2:0] _T_209 ;  
   wire _T_211 ;  
   wire _T_212 ;  
   wire [2:0] _T_213 ;  
   wire _T_215 ;  
   wire _T_216 ;  
   wire [2:0] _T_217 ;  
   wire [1:0] _T_218 ;  
   wire _T_219 ;  
   wire _T_220 ;  
   wire [2:0] _T_221 ;  
   wire [1:0] _T_222 ;  
   wire _T_223 ;  
   wire _T_224 ;  
   wire [2:0] _T_225 ;  
   wire [1:0] _T_226 ;  
   wire _T_227 ;  
   wire _T_228 ;  
   wire [2:0] _T_229 ;  
   wire [1:0] _T_230 ;  
   wire _T_231 ;  
   wire _T_232 ;  
   wire [2:0] _T_233 ;  
   wire [1:0] _T_234 ;  
   wire _T_235 ;  
   wire _T_236 ;  
   wire [2:0] _T_237 ;  
   wire [1:0] _T_238 ;  
   wire _T_239 ;  
   wire s2_victim_dirty ;  
   wire [2:0] s2_shrink_param ;  
   wire [1:0] voluntaryNewCoh_state ;  
   wire s2_dont_nack_uncached ;  
   wire _s2_dont_nack_misc_T_10 ;  
   wire s2_dont_nack_misc ;  
   wire _io_cpu_s2_nack_T_1 ;  
   wire _io_cpu_s2_nack_T_3 ;  
   wire _metaArb_io_in_1_valid_T ;  
   wire _metaArb_io_in_1_valid_T_1 ;  
   wire [11:0] metaArb_io_in_1_bits_addr_lo ;  
   wire [1:0] new_meta_coh_state ;  
   wire [11:0] metaArb_io_in_2_bits_addr_lo ;  
   wire [19:0] metaArb_io_in_2_bits_data_meta_tag ;  
   wire _lrscBackingOff_T ;  
   wire lrscBackingOff ;  
   reg [33:0] lrscAddr ;  
   reg [63:0] _RAND_82 ;  
   wire lrscAddrMatch ;  
   wire _s2_sc_fail_T ;  
   wire s2_sc_fail ;  
   wire _T_243 ;  
   wire _T_245 ;  
   wire _T_246 ;  
   wire [6:0] _lrscCount_T_2 ;  
   wire _T_250 ;  
   wire _pstore1_cmd_T ;  
   reg [4:0] pstore1_cmd ;  
   reg [31:0] _RAND_83 ;  
   reg [63:0] pstore1_data ;  
   reg [63:0] _RAND_84 ;  
   reg [3:0] pstore1_way ;  
   reg [31:0] _RAND_85 ;  
   wire _pstore1_rmw_T_49 ;  
   wire _pstore1_rmw_T_50 ;  
   reg pstore1_rmw_r ;  
   reg [31:0] _RAND_86 ;  
   wire _pstore1_merge_T ;  
   wire _pstore1_merge_T_2 ;  
   wire pstore_drain_opportunistic ;  
   reg pstore_drain_on_miss_REG ;  
   reg [31:0] _RAND_87 ;  
   wire pstore_drain_on_miss ;  
   wire pstore1_valid ;  
   wire _pstore_drain_structural_T ;  
   wire _pstore_drain_structural_T_1 ;  
   wire _pstore_drain_structural_T_2 ;  
   wire pstore_drain_structural ;  
   wire _T_254 ;  
   wire _T_255 ;  
   wire _T_256 ;  
   wire _T_258 ;  
   wire _pstore_drain_T_7 ;  
   wire _pstore_drain_T_8 ;  
   wire _pstore_drain_T_9 ;  
   wire _pstore_drain_T_10 ;  
   wire pstore_drain ;  
   wire _pstore1_held_T_8 ;  
   wire _pstore1_held_T_10 ;  
   wire _advance_pstore1_T_1 ;  
   wire advance_pstore1 ;  
   wire _pstore2_valid_T_1 ;  
   wire _pstore2_valid_T_2 ;  
   reg [3:0] pstore2_way ;  
   reg [31:0] _RAND_88 ;  
   wire [63:0] pstore1_storegen_data ;  
   reg [7:0] pstore2_storegen_data_lo_lo_lo ;  
   reg [31:0] _RAND_89 ;  
   reg [7:0] pstore2_storegen_data_lo_lo_hi ;  
   reg [31:0] _RAND_90 ;  
   reg [7:0] pstore2_storegen_data_lo_hi_lo ;  
   reg [31:0] _RAND_91 ;  
   reg [7:0] pstore2_storegen_data_lo_hi_hi ;  
   reg [31:0] _RAND_92 ;  
   reg [7:0] pstore2_storegen_data_hi_lo_lo ;  
   reg [31:0] _RAND_93 ;  
   reg [7:0] pstore2_storegen_data_hi_lo_hi ;  
   reg [31:0] _RAND_94 ;  
   reg [7:0] pstore2_storegen_data_hi_hi_lo ;  
   reg [31:0] _RAND_95 ;  
   reg [7:0] pstore2_storegen_data_hi_hi_hi ;  
   reg [31:0] _RAND_96 ;  
   wire [63:0] pstore2_storegen_data ;  
   wire [39:0] _dataArb_io_in_0_bits_addr_T ;  
   wire [63:0] _dataArb_io_in_0_bits_wdata_T ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_lo_lo_lo ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_lo_lo_hi ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_lo_hi_lo ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_lo_hi_hi ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_hi_lo_lo ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_hi_lo_hi ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_hi_hi_lo ;  
   wire [7:0] dataArb_io_in_0_bits_wdata_hi_hi_hi ;  
   wire [31:0] dataArb_io_in_0_bits_wdata_lo ;  
   wire [31:0] dataArb_io_in_0_bits_wdata_hi ;  
   wire [7:0] _dataArb_io_in_0_bits_eccMask_T ;  
   wire dataArb_io_in_0_bits_eccMask_lo_lo_lo ;  
   wire dataArb_io_in_0_bits_eccMask_lo_lo_hi ;  
   wire dataArb_io_in_0_bits_eccMask_lo_hi_lo ;  
   wire dataArb_io_in_0_bits_eccMask_lo_hi_hi ;  
   wire dataArb_io_in_0_bits_eccMask_hi_lo_lo ;  
   wire dataArb_io_in_0_bits_eccMask_hi_lo_hi ;  
   wire dataArb_io_in_0_bits_eccMask_hi_hi_lo ;  
   wire dataArb_io_in_0_bits_eccMask_hi_hi_hi ;  
   wire [3:0] dataArb_io_in_0_bits_eccMask_lo ;  
   wire [3:0] dataArb_io_in_0_bits_eccMask_hi ;  
   wire [1:0] _a_source_T_1 ;  
   wire a_source ;  
   wire [39:0] acquire_address ;  
   wire [22:0] a_mask ;  
   wire [2:0] _get_a_mask_sizeOH_T ;  
   wire [1:0] get_a_mask_sizeOH_shiftAmount ;  
   wire [3:0] _get_a_mask_sizeOH_T_1 ;  
   wire [2:0] get_a_mask_sizeOH ;  
   wire _get_a_mask_T ;  
   wire get_a_mask_size ;  
   wire get_a_mask_bit ;  
   wire get_a_mask_nbit ;  
   wire _get_a_mask_acc_T ;  
   wire get_a_mask_acc ;  
   wire _get_a_mask_acc_T_1 ;  
   wire get_a_mask_acc_1 ;  
   wire get_a_mask_size_1 ;  
   wire get_a_mask_bit_1 ;  
   wire get_a_mask_nbit_1 ;  
   wire get_a_mask_eq_2 ;  
   wire _get_a_mask_acc_T_2 ;  
   wire get_a_mask_acc_2 ;  
   wire get_a_mask_eq_3 ;  
   wire _get_a_mask_acc_T_3 ;  
   wire get_a_mask_acc_3 ;  
   wire get_a_mask_eq_4 ;  
   wire _get_a_mask_acc_T_4 ;  
   wire get_a_mask_acc_4 ;  
   wire get_a_mask_eq_5 ;  
   wire _get_a_mask_acc_T_5 ;  
   wire get_a_mask_acc_5 ;  
   wire get_a_mask_size_2 ;  
   wire get_a_mask_bit_2 ;  
   wire get_a_mask_nbit_2 ;  
   wire get_a_mask_eq_6 ;  
   wire _get_a_mask_acc_T_6 ;  
   wire get_a_mask_lo_lo_lo ;  
   wire get_a_mask_eq_7 ;  
   wire _get_a_mask_acc_T_7 ;  
   wire get_a_mask_lo_lo_hi ;  
   wire get_a_mask_eq_8 ;  
   wire _get_a_mask_acc_T_8 ;  
   wire get_a_mask_lo_hi_lo ;  
   wire get_a_mask_eq_9 ;  
   wire _get_a_mask_acc_T_9 ;  
   wire get_a_mask_lo_hi_hi ;  
   wire get_a_mask_eq_10 ;  
   wire _get_a_mask_acc_T_10 ;  
   wire get_a_mask_hi_lo_lo ;  
   wire get_a_mask_eq_11 ;  
   wire _get_a_mask_acc_T_11 ;  
   wire get_a_mask_hi_lo_hi ;  
   wire get_a_mask_eq_12 ;  
   wire _get_a_mask_acc_T_12 ;  
   wire get_a_mask_hi_hi_lo ;  
   wire get_a_mask_eq_13 ;  
   wire _get_a_mask_acc_T_13 ;  
   wire get_a_mask_hi_hi_hi ;  
   wire [7:0] get_mask ;  
   wire _atomics_T ;  
   wire [2:0] _atomics_T_1_opcode ;  
   wire [3:0] atomics_a_size ;  
   wire [3:0] _atomics_T_1_size ;  
   wire _atomics_T_1_source ;  
   wire [31:0] atomics_a_address ;  
   wire [31:0] _atomics_T_1_address ;  
   wire [7:0] _atomics_T_1_mask ;  
   wire [63:0] _atomics_T_1_data ;  
   wire _atomics_T_2 ;  
   wire [2:0] _atomics_T_3_opcode ;  
   wire [2:0] _atomics_T_3_param ;  
   wire [3:0] _atomics_T_3_size ;  
   wire _atomics_T_3_source ;  
   wire [31:0] _atomics_T_3_address ;  
   wire [7:0] _atomics_T_3_mask ;  
   wire [63:0] _atomics_T_3_data ;  
   wire _atomics_T_4 ;  
   wire [2:0] _atomics_T_5_opcode ;  
   wire [2:0] _atomics_T_5_param ;  
   wire [3:0] _atomics_T_5_size ;  
   wire _atomics_T_5_source ;  
   wire [31:0] _atomics_T_5_address ;  
   wire [7:0] _atomics_T_5_mask ;  
   wire [63:0] _atomics_T_5_data ;  
   wire _atomics_T_6 ;  
   wire [2:0] _atomics_T_7_opcode ;  
   wire [2:0] _atomics_T_7_param ;  
   wire [3:0] _atomics_T_7_size ;  
   wire _atomics_T_7_source ;  
   wire [31:0] _atomics_T_7_address ;  
   wire [7:0] _atomics_T_7_mask ;  
   wire [63:0] _atomics_T_7_data ;  
   wire _atomics_T_8 ;  
   wire [2:0] _atomics_T_9_opcode ;  
   wire [2:0] _atomics_T_9_param ;  
   wire [3:0] _atomics_T_9_size ;  
   wire _atomics_T_9_source ;  
   wire [31:0] _atomics_T_9_address ;  
   wire [7:0] _atomics_T_9_mask ;  
   wire [63:0] _atomics_T_9_data ;  
   wire _atomics_T_10 ;  
   wire [2:0] _atomics_T_11_opcode ;  
   wire [2:0] _atomics_T_11_param ;  
   wire [3:0] _atomics_T_11_size ;  
   wire _atomics_T_11_source ;  
   wire [31:0] _atomics_T_11_address ;  
   wire [7:0] _atomics_T_11_mask ;  
   wire [63:0] _atomics_T_11_data ;  
   wire _atomics_T_12 ;  
   wire [2:0] _atomics_T_13_opcode ;  
   wire [2:0] _atomics_T_13_param ;  
   wire [3:0] _atomics_T_13_size ;  
   wire _atomics_T_13_source ;  
   wire [31:0] _atomics_T_13_address ;  
   wire [7:0] _atomics_T_13_mask ;  
   wire [63:0] _atomics_T_13_data ;  
   wire _atomics_T_14 ;  
   wire [2:0] _atomics_T_15_opcode ;  
   wire [2:0] _atomics_T_15_param ;  
   wire [3:0] _atomics_T_15_size ;  
   wire _atomics_T_15_source ;  
   wire [31:0] _atomics_T_15_address ;  
   wire [7:0] _atomics_T_15_mask ;  
   wire [63:0] _atomics_T_15_data ;  
   wire _atomics_T_16 ;  
   wire [2:0] atomics_opcode ;  
   wire [2:0] atomics_param ;  
   wire [3:0] atomics_size ;  
   wire atomics_source ;  
   wire [31:0] atomics_address ;  
   wire [7:0] atomics_mask ;  
   wire [63:0] atomics_data ;  
   wire [39:0] _GEN_356 ;  
   wire [39:0] _tl_out_a_valid_T_1 ;  
   wire _tl_out_a_valid_T_3 ;  
   wire _tl_out_a_valid_T_4 ;  
   wire _tl_out_a_valid_T_6 ;  
   wire _tl_out_a_valid_T_12 ;  
   wire tl_out_a_valid ;  
   wire [2:0] _tl_out_a_bits_T_6_opcode ;  
   wire [2:0] _tl_out_a_bits_T_6_param ;  
   wire [3:0] _tl_out_a_bits_T_6_size ;  
   wire _tl_out_a_bits_T_6_source ;  
   wire [31:0] _tl_out_a_bits_T_6_address ;  
   wire [7:0] _tl_out_a_bits_T_6_mask ;  
   wire [63:0] _tl_out_a_bits_T_6_data ;  
   wire [2:0] _tl_out_a_bits_T_7_opcode ;  
   wire [2:0] _tl_out_a_bits_T_7_param ;  
   wire [3:0] _tl_out_a_bits_T_7_size ;  
   wire _tl_out_a_bits_T_7_source ;  
   wire [31:0] _tl_out_a_bits_T_7_address ;  
   wire [7:0] putpartial_mask ;  
   wire [7:0] _tl_out_a_bits_T_7_mask ;  
   wire [63:0] _tl_out_a_bits_T_7_data ;  
   wire [2:0] _tl_out_a_bits_T_8_opcode ;  
   wire [2:0] _tl_out_a_bits_T_8_param ;  
   wire [3:0] _tl_out_a_bits_T_8_size ;  
   wire _tl_out_a_bits_T_8_source ;  
   wire [31:0] _tl_out_a_bits_T_8_address ;  
   wire [7:0] _tl_out_a_bits_T_8_mask ;  
   wire [63:0] _tl_out_a_bits_T_8_data ;  
   wire [2:0] tl_out_a_bits_a_param ;  
   wire [31:0] tl_out_a_bits_a_address ;  
   wire [1:0] _a_sel_T ;  
   wire a_sel ;  
   wire _T_263 ;  
   wire _GEN_142 ;  
   wire [26:0] _beats1_decode_T_1 ;  
   wire [8:0] beats1_decode ;  
   wire beats1_opdata ;  
   wire [8:0] beats1 ;  
   wire [8:0] counter1 ;  
   wire _last_T ;  
   wire _last_T_1 ;  
   wire d_last ;  
   wire d_done ;  
   wire [8:0] count ;  
   wire [11:0] d_address_inc ;  
   wire grantIsVoluntary ;  
   wire [2:0] _blockProbeAfterGrantCount_T_1 ;  
   wire [1:0] _uncachedRespIdxOH_T ;  
   wire uncachedRespIdxOH ;  
   wire _T_273 ;  
   wire _T_276 ;  
   wire _T_278 ;  
   wire [31:0] dontCareBits ;  
   wire [31:0] _GEN_357 ;  
   wire [31:0] _s2_req_addr_T_1 ;  
   wire _T_281 ;  
   wire _GEN_196 ;  
   wire _GEN_205 ;  
   wire _GEN_209 ;  
   wire _GEN_218 ;  
   wire _GEN_231 ;  
   wire _bundleOut_0_e_valid_T ;  
   wire _bundleOut_0_e_valid_T_1 ;  
   wire _bundleOut_0_e_valid_T_2 ;  
   wire tl_out__e_valid ;  
   wire _T_283 ;  
   wire _T_285 ;  
   wire _T_286 ;  
   wire _T_287 ;  
   wire _T_289 ;  
   wire _dataArb_io_in_1_valid_T ;  
   wire _dataArb_io_in_1_valid_T_1 ;  
   wire [39:0] _dataArb_io_in_1_bits_addr_T_1 ;  
   wire [39:0] _GEN_358 ;  
   wire [39:0] _dataArb_io_in_1_bits_addr_T_2 ;  
   wire _metaArb_io_in_3_valid_T ;  
   wire [3:0] _metaArb_io_in_3_bits_data_T_1 ;  
   wire _metaArb_io_in_3_bits_data_T_6 ;  
   wire [1:0] _metaArb_io_in_3_bits_data_T_7 ;  
   wire _metaArb_io_in_3_bits_data_T_8 ;  
   wire [1:0] _metaArb_io_in_3_bits_data_T_9 ;  
   wire _metaArb_io_in_3_bits_data_T_10 ;  
   wire [1:0] _metaArb_io_in_3_bits_data_T_11 ;  
   wire _metaArb_io_in_3_bits_data_T_12 ;  
   wire [1:0] metaArb_io_in_3_bits_data_meta_state ;  
   wire _GEN_234 ;  
   wire _GEN_235 ;  
   wire _GEN_236 ;  
   wire _metaArb_io_in_6_valid_T_1 ;  
   wire _metaArb_io_in_6_valid_T_2 ;  
   wire [7:0] metaArb_io_in_6_bits_addr_hi ;  
   wire [39:0] _metaArb_io_in_6_bits_addr_T ;  
   wire [8:0] counter1_1 ;  
   wire [8:0] c_count ;  
   reg s1_release_data_valid ;  
   reg [31:0] _RAND_97 ;  
   wire releaseRejected ;  
   wire [9:0] _releaseDataBeat_T ;  
   wire [1:0] _releaseDataBeat_T_1 ;  
   wire [1:0] _GEN_359 ;  
   wire [1:0] _releaseDataBeat_T_3 ;  
   wire [1:0] _releaseDataBeat_T_4 ;  
   wire [9:0] _GEN_360 ;  
   wire [9:0] releaseDataBeat ;  
   wire _T_298 ;  
   wire _T_299 ;  
   wire _T_301 ;  
   wire discard_line ;  
   wire _release_state_T_1 ;  
   wire [3:0] _release_state_T_13 ;  
   wire [5:0] probe_bits_lo ;  
   wire [25:0] _probe_bits_T_1 ;  
   wire [31:0] res_2_address ;  
   wire [3:0] _GEN_244 ;  
   wire [3:0] _release_state_T_14 ;  
   wire [3:0] _release_state_T_15 ;  
   wire [2:0] _GEN_255 ;  
   wire [3:0] _GEN_261 ;  
   wire [3:0] _GEN_263 ;  
   wire [2:0] _GEN_266 ;  
   wire [3:0] _GEN_273 ;  
   wire [2:0] _GEN_276 ;  
   wire [3:0] _GEN_284 ;  
   wire [2:0] _GEN_287 ;  
   wire _T_304 ;  
   wire [39:0] _metaArb_io_in_6_bits_addr_T_1 ;  
   wire [3:0] _GEN_294 ;  
   wire _GEN_295 ;  
   wire [3:0] _GEN_299 ;  
   wire [3:0] _GEN_301 ;  
   wire [3:0] _GEN_303 ;  
   wire [2:0] _GEN_307 ;  
   wire [2:0] _GEN_316 ;  
   wire _T_315 ;  
   wire _GEN_331 ;  
   wire [1:0] newCoh_state ;  
   wire _dataArb_io_in_2_valid_T ;  
   wire [11:0] _dataArb_io_in_2_bits_addr_T_1 ;  
   wire [5:0] _dataArb_io_in_2_bits_addr_T_3 ;  
   wire [11:0] _GEN_363 ;  
   wire _metaArb_io_in_4_valid_T_1 ;  
   wire [11:0] metaArb_io_in_4_bits_addr_lo ;  
   wire [19:0] metaArb_io_in_4_bits_data_meta_tag ;  
   wire _T_316 ;  
   wire _io_cpu_ordered_T_4 ;  
   wire _io_cpu_ordered_T_5 ;  
   wire _io_cpu_ordered_T_7 ;  
   wire _s1_xcpt_valid_T_1 ;  
   reg io_cpu_s2_xcpt_REG ;  
   reg [31:0] _RAND_98 ;  
   reg doUncachedResp ;  
   reg [31:0] _RAND_99 ;  
   wire _T_321 ;  
   wire [31:0] io_cpu_resp_bits_data_shifted ;  
   wire _io_cpu_resp_bits_data_T ;  
   wire _io_cpu_resp_bits_data_T_3 ;  
   wire [31:0] _io_cpu_resp_bits_data_T_5 ;  
   wire [31:0] io_cpu_resp_bits_data_hi ;  
   wire [63:0] _io_cpu_resp_bits_data_T_7 ;  
   wire [15:0] io_cpu_resp_bits_data_shifted_1 ;  
   wire _io_cpu_resp_bits_data_T_8 ;  
   wire _io_cpu_resp_bits_data_T_11 ;  
   wire [47:0] _io_cpu_resp_bits_data_T_13 ;  
   wire [47:0] io_cpu_resp_bits_data_hi_1 ;  
   wire [63:0] _io_cpu_resp_bits_data_T_15 ;  
   wire [7:0] io_cpu_resp_bits_data_shifted_2 ;  
   wire [7:0] io_cpu_resp_bits_data_lo_2 ;  
   wire _io_cpu_resp_bits_data_T_16 ;  
   wire _io_cpu_resp_bits_data_T_17 ;  
   wire _io_cpu_resp_bits_data_T_19 ;  
   wire [55:0] _io_cpu_resp_bits_data_T_21 ;  
   wire [55:0] io_cpu_resp_bits_data_hi_2 ;  
   wire [63:0] _io_cpu_resp_bits_data_T_23 ;  
   wire [63:0] _GEN_364 ;  
   reg REG ;  
   reg [31:0] _RAND_100 ;  
   wire _GEN_349 ;  
   wire [8:0] flushCounterNext ;  
   wire flushDone ;  
   wire _s1_flush_valid_T ;  
   wire _s1_flush_valid_T_2 ;  
   wire _s1_flush_valid_T_4 ;  
   wire _s1_flush_valid_T_6 ;  
   wire [11:0] metaArb_io_in_5_bits_addr_lo ;  
   wire [8:0] _GEN_351 ;  
   reg [8:0] io_cpu_perf_release_counter ;  
   reg [31:0] _RAND_101 ;  
   wire [8:0] io_cpu_perf_release_counter1 ;  
   wire io_cpu_perf_release_first ;  
   wire _io_cpu_perf_release_last_T ;  
   wire io_cpu_perf_release_last ;  
   wire _GEN_367 ;  
   wire _GEN_370 ;  
   wire _GEN_371 ;  
   wire _GEN_372 ;  
   wire _GEN_380 ;  
   wire _GEN_381 ;  
   reg [19:0] DCache_state ;  
   reg [31:0] _RAND_102 ;  
   reg DCache_cov[0:1048575] ;  
   reg [31:0] _RAND_103 ;  
   wire DCache_cov_read_data ;  
   wire [19:0] DCache_cov_read_addr ;  
   wire DCache_cov_write_data ;  
   wire [19:0] DCache_cov_write_addr ;  
   wire DCache_cov_write_mask ;  
   wire DCache_cov_write_en ;  
   reg [29:0] DCache_covSum ;  
   reg [31:0] _RAND_104 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire mux_cond_4 ;  
   wire mux_cond_5 ;  
   wire [4:0] s2_req_size_shl ;  
   wire [19:0] s2_req_size_pad ;  
   wire [9:0] pstore1_held_shl ;  
   wire [19:0] pstore1_held_pad ;  
   wire [5:0] s2_req_signed_shl ;  
   wire [19:0] s2_req_signed_pad ;  
   wire [10:0] pstore2_valid_shl ;  
   wire [19:0] pstore2_valid_pad ;  
   wire [17:0] s1_flush_valid_shl ;  
   wire [19:0] s1_flush_valid_pad ;  
   wire [8:0] uncachedInFlight_0_shl ;  
   wire [19:0] uncachedInFlight_0_pad ;  
   wire [18:0] blockUncachedGrant_shl ;  
   wire [19:0] blockUncachedGrant_pad ;  
   wire [13:0] probe_bits_param_shl ;  
   wire [19:0] probe_bits_param_pad ;  
   wire [16:0] s2_flush_valid_pre_tag_ecc_shl ;  
   wire [19:0] s2_flush_valid_pre_tag_ecc_pad ;  
   wire [10:0] s1_read_mask_shl ;  
   wire [19:0] s1_read_mask_pad ;  
   wire [13:0] s2_victim_way_r_shl ;  
   wire [19:0] s2_victim_way_r_pad ;  
   wire [13:0] s1_probe_shl ;  
   wire [19:0] s1_probe_pad ;  
   wire [2:0] release_ack_wait_shl ;  
   wire [19:0] release_ack_wait_pad ;  
   wire [12:0] s2_hit_state_state_shl ;  
   wire [19:0] s2_hit_state_state_pad ;  
   wire [15:0] cached_grant_wait_shl ;  
   wire [19:0] cached_grant_wait_pad ;  
   wire [19:0] s1_valid_shl ;  
   wire [19:0] s1_valid_pad ;  
   wire [18:0] s2_pma_cacheable_shl ;  
   wire [19:0] s2_pma_cacheable_pad ;  
   wire [17:0] s1_did_read_shl ;  
   wire [19:0] s1_did_read_pad ;  
   wire [19:0] s2_probe_shl ;  
   wire [19:0] s2_probe_pad ;  
   wire [6:0] s2_hit_way_shl ;  
   wire [19:0] s2_hit_way_pad ;  
   wire [9:0] s2_not_nacked_in_s1_shl ;  
   wire [19:0] s2_not_nacked_in_s1_pad ;  
   wire [18:0] s2_probe_state_state_shl ;  
   wire [19:0] s2_probe_state_state_pad ;  
   wire [4:0] s1_req_size_shl ;  
   wire [19:0] s1_req_size_pad ;  
   wire [14:0] pstore1_rmw_r_shl ;  
   wire [19:0] pstore1_rmw_r_pad ;  
   wire [7:0] s2_release_data_valid_shl ;  
   wire [19:0] s2_release_data_valid_pad ;  
   wire [8:0] s2_valid_shl ;  
   wire [19:0] s2_valid_pad ;  
   wire [19:0] pstore_drain_on_miss_REG_shl ;  
   wire [19:0] pstore_drain_on_miss_REG_pad ;  
   wire [15:0] resetting_shl ;  
   wire [19:0] resetting_pad ;  
   wire [19:0] grantInProgress_shl ;  
   wire [19:0] grantInProgress_pad ;  
   wire [12:0] s2_probe_way_shl ;  
   wire [19:0] s2_probe_way_pad ;  
   wire [11:0] mux_cond_0_shl ;  
   wire [19:0] mux_cond_0_pad ;  
   wire [1:0] mux_cond_1_shl ;  
   wire [19:0] mux_cond_1_pad ;  
   wire [15:0] mux_cond_2_shl ;  
   wire [19:0] mux_cond_2_pad ;  
   wire [6:0] mux_cond_3_shl ;  
   wire [19:0] mux_cond_3_pad ;  
   wire [7:0] mux_cond_4_shl ;  
   wire [19:0] mux_cond_4_pad ;  
   wire [7:0] mux_cond_5_shl ;  
   wire [19:0] mux_cond_5_pad ;  
   wire [19:0] DCache_xor15 ;  
   wire [19:0] DCache_xor16 ;  
   wire [19:0] DCache_xor7 ;  
   wire [19:0] DCache_xor17 ;  
   wire [19:0] DCache_xor38 ;  
   wire [19:0] DCache_xor18 ;  
   wire [19:0] DCache_xor8 ;  
   wire [19:0] DCache_xor3 ;  
   wire [19:0] DCache_xor19 ;  
   wire [19:0] DCache_xor20 ;  
   wire [19:0] DCache_xor9 ;  
   wire [19:0] DCache_xor21 ;  
   wire [19:0] DCache_xor46 ;  
   wire [19:0] DCache_xor22 ;  
   wire [19:0] DCache_xor10 ;  
   wire [19:0] DCache_xor4 ;  
   wire [19:0] DCache_xor1 ;  
   wire [19:0] DCache_xor23 ;  
   wire [19:0] DCache_xor24 ;  
   wire [19:0] DCache_xor11 ;  
   wire [19:0] DCache_xor25 ;  
   wire [19:0] DCache_xor54 ;  
   wire [19:0] DCache_xor26 ;  
   wire [19:0] DCache_xor12 ;  
   wire [19:0] DCache_xor5 ;  
   wire [19:0] DCache_xor27 ;  
   wire [19:0] DCache_xor28 ;  
   wire [19:0] DCache_xor13 ;  
   wire [19:0] DCache_xor29 ;  
   wire [19:0] DCache_xor62 ;  
   wire [19:0] DCache_xor30 ;  
   wire [19:0] DCache_xor14 ;  
   wire [19:0] DCache_xor6 ;  
   wire [19:0] DCache_xor2 ;  
   wire [19:0] DCache_xor0 ;  
   wire [29:0] data_sum ;  
   wire [29:0] tlb_sum ;  
   wire [29:0] pma_checker_sum ;  
   wire [29:0] metaArb_sum ;  
   wire [29:0] lfsr_prng_sum ;  
   wire [29:0] amoalu_sum ;  
   wire [29:0] dataArb_sum ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire stopEn2 ;  
   wire stopEn3 ;  
   wire stopEn4 ;  
   wire stopEn5 ;  
   wire stopEn6 ;  
   wire stopEn7 ;  
   wire stopEn8 ;  
   wire stopEn9 ;  
   wire dataArb_metaAssert_wire ;  
   wire metaArb_metaAssert_wire ;  
   wire lfsr_prng_metaAssert_wire ;  
   wire tlb_metaAssert_wire ;  
   wire pma_checker_metaAssert_wire ;  
   wire data_metaAssert_wire ;  
   wire amoalu_metaAssert_wire ;  
   wire DCache_or7 ;  
   wire DCache_or8 ;  
   wire DCache_or3 ;  
   wire DCache_or9 ;  
   wire DCache_or10 ;  
   wire DCache_or4 ;  
   wire DCache_or1 ;  
   wire DCache_or11 ;  
   wire DCache_or12 ;  
   wire DCache_or5 ;  
   wire DCache_or13 ;  
   wire DCache_or30 ;  
   wire DCache_or14 ;  
   wire DCache_or6 ;  
   wire DCache_or2 ;  
   wire DCache_or0 ;  
  TLB tlb(.clock(tlb_clock),.reset(tlb_reset),.io_req_ready(tlb_io_req_ready),.io_req_valid(tlb_io_req_valid),.io_req_bits_vaddr(tlb_io_req_bits_vaddr),.io_req_bits_passthrough(tlb_io_req_bits_passthrough),.io_req_bits_size(tlb_io_req_bits_size),.io_req_bits_cmd(tlb_io_req_bits_cmd),.io_resp_miss(tlb_io_resp_miss),.io_resp_paddr(tlb_io_resp_paddr),.io_resp_pf_ld(tlb_io_resp_pf_ld),.io_resp_pf_st(tlb_io_resp_pf_st),.io_resp_ae_ld(tlb_io_resp_ae_ld),.io_resp_ae_st(tlb_io_resp_ae_st),.io_resp_ma_ld(tlb_io_resp_ma_ld),.io_resp_ma_st(tlb_io_resp_ma_st),.io_resp_cacheable(tlb_io_resp_cacheable),.io_sfence_valid(tlb_io_sfence_valid),.io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),.io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),.io_sfence_bits_addr(tlb_io_sfence_bits_addr),.io_ptw_req_ready(tlb_io_ptw_req_ready),.io_ptw_req_valid(tlb_io_ptw_req_valid),.io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),.io_ptw_resp_valid(tlb_io_ptw_resp_valid),.io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),.io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),.io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),.io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),.io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),.io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),.io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),.io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),.io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),.io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),.io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),.io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),.io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),.io_ptw_status_debug(tlb_io_ptw_status_debug),.io_ptw_status_dprv(tlb_io_ptw_status_dprv),.io_ptw_status_mxr(tlb_io_ptw_status_mxr),.io_ptw_status_sum(tlb_io_ptw_status_sum),.io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),.io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),.io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),.io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),.io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),.io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),.io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),.io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),.io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),.io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),.io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),.io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),.io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),.io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),.io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),.io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),.io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),.io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),.io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),.io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),.io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),.io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),.io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),.io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),.io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),.io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),.io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),.io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),.io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),.io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),.io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),.io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),.io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),.io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),.io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),.io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),.io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),.io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),.io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),.io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),.io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),.io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),.io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),.io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),.io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),.io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),.io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),.io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),.io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),.io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),.io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),.io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),.io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),.io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),.io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),.io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),.io_covSum(tlb_io_covSum),.metaAssert(tlb_metaAssert),.metaReset(tlb_metaReset)); 
  TLB pma_checker(.clock(pma_checker_clock),.reset(pma_checker_reset),.io_req_ready(pma_checker_io_req_ready),.io_req_valid(pma_checker_io_req_valid),.io_req_bits_vaddr(pma_checker_io_req_bits_vaddr),.io_req_bits_passthrough(pma_checker_io_req_bits_passthrough),.io_req_bits_size(pma_checker_io_req_bits_size),.io_req_bits_cmd(pma_checker_io_req_bits_cmd),.io_resp_miss(pma_checker_io_resp_miss),.io_resp_paddr(pma_checker_io_resp_paddr),.io_resp_pf_ld(pma_checker_io_resp_pf_ld),.io_resp_pf_st(pma_checker_io_resp_pf_st),.io_resp_ae_ld(pma_checker_io_resp_ae_ld),.io_resp_ae_st(pma_checker_io_resp_ae_st),.io_resp_ma_ld(pma_checker_io_resp_ma_ld),.io_resp_ma_st(pma_checker_io_resp_ma_st),.io_resp_cacheable(pma_checker_io_resp_cacheable),.io_sfence_valid(pma_checker_io_sfence_valid),.io_sfence_bits_rs1(pma_checker_io_sfence_bits_rs1),.io_sfence_bits_rs2(pma_checker_io_sfence_bits_rs2),.io_sfence_bits_addr(pma_checker_io_sfence_bits_addr),.io_ptw_req_ready(pma_checker_io_ptw_req_ready),.io_ptw_req_valid(pma_checker_io_ptw_req_valid),.io_ptw_req_bits_bits_addr(pma_checker_io_ptw_req_bits_bits_addr),.io_ptw_resp_valid(pma_checker_io_ptw_resp_valid),.io_ptw_resp_bits_ae(pma_checker_io_ptw_resp_bits_ae),.io_ptw_resp_bits_pte_ppn(pma_checker_io_ptw_resp_bits_pte_ppn),.io_ptw_resp_bits_pte_d(pma_checker_io_ptw_resp_bits_pte_d),.io_ptw_resp_bits_pte_a(pma_checker_io_ptw_resp_bits_pte_a),.io_ptw_resp_bits_pte_g(pma_checker_io_ptw_resp_bits_pte_g),.io_ptw_resp_bits_pte_u(pma_checker_io_ptw_resp_bits_pte_u),.io_ptw_resp_bits_pte_x(pma_checker_io_ptw_resp_bits_pte_x),.io_ptw_resp_bits_pte_w(pma_checker_io_ptw_resp_bits_pte_w),.io_ptw_resp_bits_pte_r(pma_checker_io_ptw_resp_bits_pte_r),.io_ptw_resp_bits_pte_v(pma_checker_io_ptw_resp_bits_pte_v),.io_ptw_resp_bits_level(pma_checker_io_ptw_resp_bits_level),.io_ptw_resp_bits_homogeneous(pma_checker_io_ptw_resp_bits_homogeneous),.io_ptw_ptbr_mode(pma_checker_io_ptw_ptbr_mode),.io_ptw_status_debug(pma_checker_io_ptw_status_debug),.io_ptw_status_dprv(pma_checker_io_ptw_status_dprv),.io_ptw_status_mxr(pma_checker_io_ptw_status_mxr),.io_ptw_status_sum(pma_checker_io_ptw_status_sum),.io_ptw_pmp_0_cfg_l(pma_checker_io_ptw_pmp_0_cfg_l),.io_ptw_pmp_0_cfg_a(pma_checker_io_ptw_pmp_0_cfg_a),.io_ptw_pmp_0_cfg_x(pma_checker_io_ptw_pmp_0_cfg_x),.io_ptw_pmp_0_cfg_w(pma_checker_io_ptw_pmp_0_cfg_w),.io_ptw_pmp_0_cfg_r(pma_checker_io_ptw_pmp_0_cfg_r),.io_ptw_pmp_0_addr(pma_checker_io_ptw_pmp_0_addr),.io_ptw_pmp_0_mask(pma_checker_io_ptw_pmp_0_mask),.io_ptw_pmp_1_cfg_l(pma_checker_io_ptw_pmp_1_cfg_l),.io_ptw_pmp_1_cfg_a(pma_checker_io_ptw_pmp_1_cfg_a),.io_ptw_pmp_1_cfg_x(pma_checker_io_ptw_pmp_1_cfg_x),.io_ptw_pmp_1_cfg_w(pma_checker_io_ptw_pmp_1_cfg_w),.io_ptw_pmp_1_cfg_r(pma_checker_io_ptw_pmp_1_cfg_r),.io_ptw_pmp_1_addr(pma_checker_io_ptw_pmp_1_addr),.io_ptw_pmp_1_mask(pma_checker_io_ptw_pmp_1_mask),.io_ptw_pmp_2_cfg_l(pma_checker_io_ptw_pmp_2_cfg_l),.io_ptw_pmp_2_cfg_a(pma_checker_io_ptw_pmp_2_cfg_a),.io_ptw_pmp_2_cfg_x(pma_checker_io_ptw_pmp_2_cfg_x),.io_ptw_pmp_2_cfg_w(pma_checker_io_ptw_pmp_2_cfg_w),.io_ptw_pmp_2_cfg_r(pma_checker_io_ptw_pmp_2_cfg_r),.io_ptw_pmp_2_addr(pma_checker_io_ptw_pmp_2_addr),.io_ptw_pmp_2_mask(pma_checker_io_ptw_pmp_2_mask),.io_ptw_pmp_3_cfg_l(pma_checker_io_ptw_pmp_3_cfg_l),.io_ptw_pmp_3_cfg_a(pma_checker_io_ptw_pmp_3_cfg_a),.io_ptw_pmp_3_cfg_x(pma_checker_io_ptw_pmp_3_cfg_x),.io_ptw_pmp_3_cfg_w(pma_checker_io_ptw_pmp_3_cfg_w),.io_ptw_pmp_3_cfg_r(pma_checker_io_ptw_pmp_3_cfg_r),.io_ptw_pmp_3_addr(pma_checker_io_ptw_pmp_3_addr),.io_ptw_pmp_3_mask(pma_checker_io_ptw_pmp_3_mask),.io_ptw_pmp_4_cfg_l(pma_checker_io_ptw_pmp_4_cfg_l),.io_ptw_pmp_4_cfg_a(pma_checker_io_ptw_pmp_4_cfg_a),.io_ptw_pmp_4_cfg_x(pma_checker_io_ptw_pmp_4_cfg_x),.io_ptw_pmp_4_cfg_w(pma_checker_io_ptw_pmp_4_cfg_w),.io_ptw_pmp_4_cfg_r(pma_checker_io_ptw_pmp_4_cfg_r),.io_ptw_pmp_4_addr(pma_checker_io_ptw_pmp_4_addr),.io_ptw_pmp_4_mask(pma_checker_io_ptw_pmp_4_mask),.io_ptw_pmp_5_cfg_l(pma_checker_io_ptw_pmp_5_cfg_l),.io_ptw_pmp_5_cfg_a(pma_checker_io_ptw_pmp_5_cfg_a),.io_ptw_pmp_5_cfg_x(pma_checker_io_ptw_pmp_5_cfg_x),.io_ptw_pmp_5_cfg_w(pma_checker_io_ptw_pmp_5_cfg_w),.io_ptw_pmp_5_cfg_r(pma_checker_io_ptw_pmp_5_cfg_r),.io_ptw_pmp_5_addr(pma_checker_io_ptw_pmp_5_addr),.io_ptw_pmp_5_mask(pma_checker_io_ptw_pmp_5_mask),.io_ptw_pmp_6_cfg_l(pma_checker_io_ptw_pmp_6_cfg_l),.io_ptw_pmp_6_cfg_a(pma_checker_io_ptw_pmp_6_cfg_a),.io_ptw_pmp_6_cfg_x(pma_checker_io_ptw_pmp_6_cfg_x),.io_ptw_pmp_6_cfg_w(pma_checker_io_ptw_pmp_6_cfg_w),.io_ptw_pmp_6_cfg_r(pma_checker_io_ptw_pmp_6_cfg_r),.io_ptw_pmp_6_addr(pma_checker_io_ptw_pmp_6_addr),.io_ptw_pmp_6_mask(pma_checker_io_ptw_pmp_6_mask),.io_ptw_pmp_7_cfg_l(pma_checker_io_ptw_pmp_7_cfg_l),.io_ptw_pmp_7_cfg_a(pma_checker_io_ptw_pmp_7_cfg_a),.io_ptw_pmp_7_cfg_x(pma_checker_io_ptw_pmp_7_cfg_x),.io_ptw_pmp_7_cfg_w(pma_checker_io_ptw_pmp_7_cfg_w),.io_ptw_pmp_7_cfg_r(pma_checker_io_ptw_pmp_7_cfg_r),.io_ptw_pmp_7_addr(pma_checker_io_ptw_pmp_7_addr),.io_ptw_pmp_7_mask(pma_checker_io_ptw_pmp_7_mask),.io_covSum(pma_checker_io_covSum),.metaAssert(pma_checker_metaAssert),.metaReset(pma_checker_metaReset)); 
  MaxPeriodFibonacciLFSR lfsr_prng(.clock(lfsr_prng_clock),.reset(lfsr_prng_reset),.io_increment(lfsr_prng_io_increment),.io_out_0(lfsr_prng_io_out_0),.io_out_1(lfsr_prng_io_out_1),.io_out_2(lfsr_prng_io_out_2),.io_out_3(lfsr_prng_io_out_3),.io_out_4(lfsr_prng_io_out_4),.io_out_5(lfsr_prng_io_out_5),.io_out_6(lfsr_prng_io_out_6),.io_out_7(lfsr_prng_io_out_7),.io_out_8(lfsr_prng_io_out_8),.io_out_9(lfsr_prng_io_out_9),.io_out_10(lfsr_prng_io_out_10),.io_out_11(lfsr_prng_io_out_11),.io_out_12(lfsr_prng_io_out_12),.io_out_13(lfsr_prng_io_out_13),.io_out_14(lfsr_prng_io_out_14),.io_out_15(lfsr_prng_io_out_15),.io_covSum(lfsr_prng_io_covSum),.metaAssert(lfsr_prng_metaAssert),.metaReset(lfsr_prng_metaReset)); 
  DCacheModuleImpl_Anon_1 metaArb(.io_in_0_valid(metaArb_io_in_0_valid),.io_in_0_bits_addr(metaArb_io_in_0_bits_addr),.io_in_0_bits_idx(metaArb_io_in_0_bits_idx),.io_in_1_valid(metaArb_io_in_1_valid),.io_in_1_bits_addr(metaArb_io_in_1_bits_addr),.io_in_1_bits_idx(metaArb_io_in_1_bits_idx),.io_in_1_bits_data(metaArb_io_in_1_bits_data),.io_in_2_valid(metaArb_io_in_2_valid),.io_in_2_bits_addr(metaArb_io_in_2_bits_addr),.io_in_2_bits_idx(metaArb_io_in_2_bits_idx),.io_in_2_bits_way_en(metaArb_io_in_2_bits_way_en),.io_in_2_bits_data(metaArb_io_in_2_bits_data),.io_in_3_valid(metaArb_io_in_3_valid),.io_in_3_bits_addr(metaArb_io_in_3_bits_addr),.io_in_3_bits_idx(metaArb_io_in_3_bits_idx),.io_in_3_bits_way_en(metaArb_io_in_3_bits_way_en),.io_in_3_bits_data(metaArb_io_in_3_bits_data),.io_in_4_ready(metaArb_io_in_4_ready),.io_in_4_valid(metaArb_io_in_4_valid),.io_in_4_bits_addr(metaArb_io_in_4_bits_addr),.io_in_4_bits_idx(metaArb_io_in_4_bits_idx),.io_in_4_bits_way_en(metaArb_io_in_4_bits_way_en),.io_in_4_bits_data(metaArb_io_in_4_bits_data),.io_in_5_ready(metaArb_io_in_5_ready),.io_in_5_valid(metaArb_io_in_5_valid),.io_in_5_bits_addr(metaArb_io_in_5_bits_addr),.io_in_5_bits_idx(metaArb_io_in_5_bits_idx),.io_in_6_ready(metaArb_io_in_6_ready),.io_in_6_valid(metaArb_io_in_6_valid),.io_in_6_bits_addr(metaArb_io_in_6_bits_addr),.io_in_6_bits_idx(metaArb_io_in_6_bits_idx),.io_in_6_bits_way_en(metaArb_io_in_6_bits_way_en),.io_in_6_bits_data(metaArb_io_in_6_bits_data),.io_in_7_ready(metaArb_io_in_7_ready),.io_in_7_valid(metaArb_io_in_7_valid),.io_in_7_bits_addr(metaArb_io_in_7_bits_addr),.io_in_7_bits_idx(metaArb_io_in_7_bits_idx),.io_in_7_bits_way_en(metaArb_io_in_7_bits_way_en),.io_in_7_bits_data(metaArb_io_in_7_bits_data),.io_out_valid(metaArb_io_out_valid),.io_out_bits_write(metaArb_io_out_bits_write),.io_out_bits_addr(metaArb_io_out_bits_addr),.io_out_bits_idx(metaArb_io_out_bits_idx),.io_out_bits_way_en(metaArb_io_out_bits_way_en),.io_out_bits_data(metaArb_io_out_bits_data),.io_covSum(metaArb_io_covSum),.metaAssert(metaArb_metaAssert)); 
  DCacheDataArray data(.clock(data_clock),.io_req_valid(data_io_req_valid),.io_req_bits_addr(data_io_req_bits_addr),.io_req_bits_write(data_io_req_bits_write),.io_req_bits_wdata(data_io_req_bits_wdata),.io_req_bits_eccMask(data_io_req_bits_eccMask),.io_req_bits_way_en(data_io_req_bits_way_en),.io_resp_0(data_io_resp_0),.io_resp_1(data_io_resp_1),.io_resp_2(data_io_resp_2),.io_resp_3(data_io_resp_3),.io_covSum(data_io_covSum),.metaAssert(data_metaAssert),.metaReset(data_metaReset)); 
  DCacheModuleImpl_Anon_2 dataArb(.io_in_0_valid(dataArb_io_in_0_valid),.io_in_0_bits_addr(dataArb_io_in_0_bits_addr),.io_in_0_bits_write(dataArb_io_in_0_bits_write),.io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),.io_in_0_bits_eccMask(dataArb_io_in_0_bits_eccMask),.io_in_0_bits_way_en(dataArb_io_in_0_bits_way_en),.io_in_1_ready(dataArb_io_in_1_ready),.io_in_1_valid(dataArb_io_in_1_valid),.io_in_1_bits_addr(dataArb_io_in_1_bits_addr),.io_in_1_bits_write(dataArb_io_in_1_bits_write),.io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),.io_in_1_bits_way_en(dataArb_io_in_1_bits_way_en),.io_in_2_ready(dataArb_io_in_2_ready),.io_in_2_valid(dataArb_io_in_2_valid),.io_in_2_bits_addr(dataArb_io_in_2_bits_addr),.io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),.io_in_3_ready(dataArb_io_in_3_ready),.io_in_3_valid(dataArb_io_in_3_valid),.io_in_3_bits_addr(dataArb_io_in_3_bits_addr),.io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),.io_in_3_bits_wordMask(dataArb_io_in_3_bits_wordMask),.io_out_valid(dataArb_io_out_valid),.io_out_bits_addr(dataArb_io_out_bits_addr),.io_out_bits_write(dataArb_io_out_bits_write),.io_out_bits_wdata(dataArb_io_out_bits_wdata),.io_out_bits_eccMask(dataArb_io_out_bits_eccMask),.io_out_bits_way_en(dataArb_io_out_bits_way_en),.io_covSum(dataArb_io_covSum),.metaAssert(dataArb_metaAssert)); 
  AMOALU amoalu(.io_mask(amoalu_io_mask),.io_cmd(amoalu_io_cmd),.io_lhs(amoalu_io_lhs),.io_rhs(amoalu_io_rhs),.io_out(amoalu_io_out),.io_covSum(amoalu_io_covSum),.metaAssert(amoalu_metaAssert)); 
  assign tag_array_0_s1_meta_addr=tag_array_0_s1_meta_addr_pipe_0; 
  assign tag_array_0_s1_meta_data=tag_array_0[tag_array_0_s1_meta_addr]; 
  assign tag_array_0_MPORT_data=metaArb_io_out_bits_data; 
  assign tag_array_0_MPORT_addr=metaArb_io_out_bits_idx; 
  assign tag_array_0_MPORT_mask=metaArb_io_out_bits_way_en[0]; 
  assign tag_array_0_MPORT_en=metaArb_io_out_valid&metaArb_io_out_bits_write; 
  assign tag_array_1_s1_meta_addr=tag_array_1_s1_meta_addr_pipe_0; 
  assign tag_array_1_s1_meta_data=tag_array_1[tag_array_1_s1_meta_addr]; 
  assign tag_array_1_MPORT_data=metaArb_io_out_bits_data; 
  assign tag_array_1_MPORT_addr=metaArb_io_out_bits_idx; 
  assign tag_array_1_MPORT_mask=metaArb_io_out_bits_way_en[1]; 
  assign tag_array_1_MPORT_en=metaArb_io_out_valid&metaArb_io_out_bits_write; 
  assign tag_array_2_s1_meta_addr=tag_array_2_s1_meta_addr_pipe_0; 
  assign tag_array_2_s1_meta_data=tag_array_2[tag_array_2_s1_meta_addr]; 
  assign tag_array_2_MPORT_data=metaArb_io_out_bits_data; 
  assign tag_array_2_MPORT_addr=metaArb_io_out_bits_idx; 
  assign tag_array_2_MPORT_mask=metaArb_io_out_bits_way_en[2]; 
  assign tag_array_2_MPORT_en=metaArb_io_out_valid&metaArb_io_out_bits_write; 
  assign tag_array_3_s1_meta_addr=tag_array_3_s1_meta_addr_pipe_0; 
  assign tag_array_3_s1_meta_data=tag_array_3[tag_array_3_s1_meta_addr]; 
  assign tag_array_3_MPORT_data=metaArb_io_out_bits_data; 
  assign tag_array_3_MPORT_addr=metaArb_io_out_bits_idx; 
  assign tag_array_3_MPORT_mask=metaArb_io_out_bits_way_en[3]; 
  assign tag_array_3_MPORT_en=metaArb_io_out_valid&metaArb_io_out_bits_write; 
  assign lfsr_lo={lfsr_prng_io_out_7,lfsr_prng_io_out_6,lfsr_prng_io_out_5,lfsr_prng_io_out_4,lfsr_prng_io_out_3,lfsr_prng_io_out_2,lfsr_prng_io_out_1,lfsr_prng_io_out_0}; 
  assign lfsr={lfsr_prng_io_out_15,lfsr_prng_io_out_14,lfsr_prng_io_out_13,lfsr_prng_io_out_12,lfsr_prng_io_out_11,lfsr_prng_io_out_10,lfsr_prng_io_out_9,lfsr_prng_io_out_8,lfsr_lo}; 
  assign s1_valid_x9=io_cpu_req_ready&io_cpu_req_valid; 
  assign _block_probe_for_core_progress_T=blockProbeAfterGrantCount>3'h0; 
  assign lrscValid=lrscCount>7'h3; 
  assign block_probe_for_core_progress=_block_probe_for_core_progress_T|lrscValid; 
  assign _releaseInFlight_T=s1_probe|s2_probe; 
  assign _releaseInFlight_T_1=release_state!=4'h0; 
  assign releaseInFlight=_releaseInFlight_T|_releaseInFlight_T_1; 
  assign _block_probe_for_pending_release_ack_T=auto_out_b_bits_address^release_ack_addr; 
  assign _block_probe_for_pending_release_ack_T_2=_block_probe_for_pending_release_ack_T[20:6]==15'h0; 
  assign block_probe_for_pending_release_ack=release_ack_wait&_block_probe_for_pending_release_ack_T_2; 
  assign _block_probe_for_ordering_T=releaseInFlight|block_probe_for_pending_release_ack; 
  assign block_probe_for_ordering=_block_probe_for_ordering_T|grantInProgress; 
  assign _bundleOut_0_b_ready_T=block_probe_for_core_progress|block_probe_for_ordering; 
  assign _bundleOut_0_b_ready_T_1=_bundleOut_0_b_ready_T|s1_valid; 
  assign _bundleOut_0_b_ready_T_2=_bundleOut_0_b_ready_T_1|s2_valid; 
  assign tl_out__b_ready=metaArb_io_in_6_ready&~_bundleOut_0_b_ready_T_2; 
  assign s1_probe_x12=tl_out__b_ready&auto_out_b_valid; 
  assign s1_valid_masked=s1_valid&~io_cpu_s1_kill; 
  assign s2_meta_error=|4'h0; 
  assign _T_118={probe_bits_param,s2_probe_state_state}; 
  assign _T_175=4'h3==_T_118; 
  assign _T_171=4'h2==_T_118; 
  assign _T_167=4'h1==_T_118; 
  assign _T_163=4'h0==_T_118; 
  assign _T_159=4'h7==_T_118; 
  assign _T_155=4'h6==_T_118; 
  assign _T_151=4'h5==_T_118; 
  assign _T_147=4'h4==_T_118; 
  assign _T_143=4'hb==_T_118; 
  assign _T_139=4'ha==_T_118; 
  assign _T_135=4'h9==_T_118; 
  assign _T_131=4'h8==_T_118; 
  assign _T_148=_T_147 ? 1'h0:_T_143; 
  assign _T_152=_T_151 ? 1'h0:_T_148; 
  assign _T_156=_T_155 ? 1'h0:_T_152; 
  assign _T_160=_T_159|_T_156; 
  assign _T_164=_T_163 ? 1'h0:_T_160; 
  assign _T_168=_T_167 ? 1'h0:_T_164; 
  assign _T_172=_T_171 ? 1'h0:_T_168; 
  assign s2_prb_ack_data=_T_175|_T_172; 
  assign _T_303=s2_probe_state_state>2'h0; 
  assign _last_T_2=counter_1==9'h1; 
  assign _T_308=release_state==4'h1; 
  assign _T_309=release_state==4'h6; 
  assign _T_311=_T_308|_T_309; 
  assign _T_310=release_state==4'h9; 
  assign _T_312=_T_311|_T_310; 
  assign _GEN_323=_T_310 ? 3'h6:3'h7; 
  assign _T_307=release_state==4'h2; 
  assign _T_306=release_state==4'h3; 
  assign _GEN_315=_T_307 ? 3'h5:3'h4; 
  assign tl_out__c_bits_opcode=_T_312 ? _GEN_323:_GEN_315; 
  assign beats1_opdata_1=tl_out__c_bits_opcode[0]; 
  assign tl_out__c_bits_size=_T_312 ? 4'h6:probe_bits_size; 
  assign _beats1_decode_T_5=27'hfff<<tl_out__c_bits_size; 
  assign beats1_decode_1=~_beats1_decode_T_5[11:3]; 
  assign beats1_1=beats1_opdata_1 ? beats1_decode_1:9'h0; 
  assign _last_T_3=beats1_1==9'h0; 
  assign c_last=_last_T_2|_last_T_3; 
  assign _T_305=release_state==4'h5; 
  assign c_first=counter_1==9'h0; 
  assign _bundleOut_0_c_valid_T_3=c_first&release_ack_wait; 
  assign _bundleOut_0_c_valid_T_5=s2_release_data_valid&~_bundleOut_0_c_valid_T_3; 
  assign _GEN_264=s2_prb_ack_data ? _bundleOut_0_c_valid_T_5:1'h1; 
  assign _GEN_274=s2_meta_error ? _bundleOut_0_c_valid_T_5:_GEN_264; 
  assign _GEN_285=s2_probe ? _GEN_274:_bundleOut_0_c_valid_T_5; 
  assign _GEN_302=_T_305|_GEN_285; 
  assign tl_out__c_valid=_T_306|_GEN_302; 
  assign _T_297=auto_out_c_ready&tl_out__c_valid; 
  assign releaseDone=c_last&_T_297; 
  assign _GEN_262=_T_303|~releaseDone; 
  assign _GEN_272=s2_prb_ack_data|_GEN_262; 
  assign probeNack=s2_meta_error|_GEN_272; 
  assign _s1_read_T=s1_req_cmd==5'h0; 
  assign _s1_read_T_1=s1_req_cmd==5'h6; 
  assign _s1_read_T_2=_s1_read_T|_s1_read_T_1; 
  assign _s1_read_T_3=s1_req_cmd==5'h7; 
  assign _s1_read_T_4=_s1_read_T_2|_s1_read_T_3; 
  assign _s1_read_T_5=s1_req_cmd==5'h4; 
  assign _s1_read_T_6=s1_req_cmd==5'h9; 
  assign _s1_read_T_9=_s1_read_T_5|_s1_read_T_6; 
  assign _s1_read_T_7=s1_req_cmd==5'ha; 
  assign _s1_read_T_10=_s1_read_T_9|_s1_read_T_7; 
  assign _s1_read_T_8=s1_req_cmd==5'hb; 
  assign _s1_read_T_11=_s1_read_T_10|_s1_read_T_8; 
  assign _s1_read_T_12=s1_req_cmd==5'h8; 
  assign _s1_read_T_13=s1_req_cmd==5'hc; 
  assign _s1_read_T_17=_s1_read_T_12|_s1_read_T_13; 
  assign _s1_read_T_14=s1_req_cmd==5'hd; 
  assign _s1_read_T_18=_s1_read_T_17|_s1_read_T_14; 
  assign _s1_read_T_15=s1_req_cmd==5'he; 
  assign _s1_read_T_19=_s1_read_T_18|_s1_read_T_15; 
  assign _s1_read_T_16=s1_req_cmd==5'hf; 
  assign _s1_read_T_20=_s1_read_T_19|_s1_read_T_16; 
  assign _s1_read_T_21=_s1_read_T_11|_s1_read_T_20; 
  assign s1_read=_s1_read_T_4|_s1_read_T_21; 
  assign _s2_write_T=s2_req_cmd==5'h1; 
  assign _s2_write_T_1=s2_req_cmd==5'h11; 
  assign _s2_write_T_2=_s2_write_T|_s2_write_T_1; 
  assign _s2_write_T_3=s2_req_cmd==5'h7; 
  assign _s2_write_T_4=_s2_write_T_2|_s2_write_T_3; 
  assign _s2_write_T_5=s2_req_cmd==5'h4; 
  assign _s2_write_T_6=s2_req_cmd==5'h9; 
  assign _s2_write_T_9=_s2_write_T_5|_s2_write_T_6; 
  assign _s2_write_T_7=s2_req_cmd==5'ha; 
  assign _s2_write_T_10=_s2_write_T_9|_s2_write_T_7; 
  assign _s2_write_T_8=s2_req_cmd==5'hb; 
  assign _s2_write_T_11=_s2_write_T_10|_s2_write_T_8; 
  assign _s2_write_T_12=s2_req_cmd==5'h8; 
  assign _s2_write_T_13=s2_req_cmd==5'hc; 
  assign _s2_write_T_17=_s2_write_T_12|_s2_write_T_13; 
  assign _s2_write_T_14=s2_req_cmd==5'hd; 
  assign _s2_write_T_18=_s2_write_T_17|_s2_write_T_14; 
  assign _s2_write_T_15=s2_req_cmd==5'he; 
  assign _s2_write_T_19=_s2_write_T_18|_s2_write_T_15; 
  assign _s2_write_T_16=s2_req_cmd==5'hf; 
  assign _s2_write_T_20=_s2_write_T_19|_s2_write_T_16; 
  assign _s2_write_T_21=_s2_write_T_11|_s2_write_T_20; 
  assign s2_write=_s2_write_T_4|_s2_write_T_21; 
  assign _pstore1_valid_likely_T=s2_valid&s2_write; 
  assign pstore1_valid_likely=_pstore1_valid_likely_T|pstore1_held; 
  assign s1_vaddr_hi=s1_req_addr[39:12]; 
  assign s1_vaddr_lo=s1_req_addr[11:0]; 
  assign s1_vaddr={s1_vaddr_hi,s1_vaddr_lo}; 
  assign _s1_hazard_T_2=pstore1_addr[11:3]==s1_vaddr[11:3]; 
  assign _s1_write_T=s1_req_cmd==5'h1; 
  assign _s1_write_T_1=s1_req_cmd==5'h11; 
  assign _s1_write_T_2=_s1_write_T|_s1_write_T_1; 
  assign _s1_write_T_4=_s1_write_T_2|_s1_read_T_3; 
  assign s1_write=_s1_write_T_4|_s1_read_T_21; 
  assign s1_hazard_hi_hi_hi=|pstore1_mask[7]; 
  assign s1_hazard_hi_hi_lo=|pstore1_mask[6]; 
  assign s1_hazard_hi_lo_hi=|pstore1_mask[5]; 
  assign s1_hazard_hi_lo_lo=|pstore1_mask[4]; 
  assign s1_hazard_lo_hi_hi=|pstore1_mask[3]; 
  assign s1_hazard_lo_hi_lo=|pstore1_mask[2]; 
  assign s1_hazard_lo_lo_hi=|pstore1_mask[1]; 
  assign s1_hazard_lo_lo_lo=|pstore1_mask[0]; 
  assign _s1_hazard_T_11={s1_hazard_hi_hi_hi,s1_hazard_hi_hi_lo,s1_hazard_hi_lo_hi,s1_hazard_hi_lo_lo,s1_hazard_lo_hi_hi,s1_hazard_lo_hi_lo,s1_hazard_lo_lo_hi,s1_hazard_lo_lo_lo}; 
  assign s1_hazard_hi_hi_hi_1=_s1_hazard_T_11[7]; 
  assign s1_hazard_hi_hi_lo_1=_s1_hazard_T_11[6]; 
  assign s1_hazard_hi_lo_hi_1=_s1_hazard_T_11[5]; 
  assign s1_hazard_hi_lo_lo_1=_s1_hazard_T_11[4]; 
  assign s1_hazard_lo_hi_hi_1=_s1_hazard_T_11[3]; 
  assign s1_hazard_lo_hi_lo_1=_s1_hazard_T_11[2]; 
  assign s1_hazard_lo_lo_hi_1=_s1_hazard_T_11[1]; 
  assign s1_hazard_lo_lo_lo_1=_s1_hazard_T_11[0]; 
  assign _s1_hazard_T_12={s1_hazard_hi_hi_hi_1,s1_hazard_hi_hi_lo_1,s1_hazard_hi_lo_hi_1,s1_hazard_hi_lo_lo_1,s1_hazard_lo_hi_hi_1,s1_hazard_lo_hi_lo_1,s1_hazard_lo_lo_hi_1,s1_hazard_lo_lo_lo_1}; 
  assign _s1_mask_xwr_upper_T_2=s1_req_size>=2'h1; 
  assign s1_mask_xwr_hi=s1_req_addr[0]|_s1_mask_xwr_upper_T_2; 
  assign s1_mask_xwr_lo=s1_req_addr[0] ? 1'h0:1'h1; 
  assign _s1_mask_xwr_T={s1_mask_xwr_hi,s1_mask_xwr_lo}; 
  assign _s1_mask_xwr_upper_T_5=s1_req_addr[1] ? _s1_mask_xwr_T:2'h0; 
  assign _s1_mask_xwr_upper_T_6=s1_req_size>=2'h2; 
  assign _s1_mask_xwr_upper_T_7=_s1_mask_xwr_upper_T_6 ? 2'h3:2'h0; 
  assign s1_mask_xwr_hi_1=_s1_mask_xwr_upper_T_5|_s1_mask_xwr_upper_T_7; 
  assign s1_mask_xwr_lo_1=s1_req_addr[1] ? 2'h0:_s1_mask_xwr_T; 
  assign _s1_mask_xwr_T_1={s1_mask_xwr_hi_1,s1_mask_xwr_lo_1}; 
  assign _s1_mask_xwr_upper_T_9=s1_req_addr[2] ? _s1_mask_xwr_T_1:4'h0; 
  assign _s1_mask_xwr_upper_T_10=s1_req_size>=2'h3; 
  assign _s1_mask_xwr_upper_T_11=_s1_mask_xwr_upper_T_10 ? 4'hf:4'h0; 
  assign s1_mask_xwr_hi_2=_s1_mask_xwr_upper_T_9|_s1_mask_xwr_upper_T_11; 
  assign s1_mask_xwr_lo_2=s1_req_addr[2] ? 4'h0:_s1_mask_xwr_T_1; 
  assign s1_mask_xwr={s1_mask_xwr_hi_2,s1_mask_xwr_lo_2}; 
  assign s1_hazard_hi_hi_hi_2=|s1_mask_xwr[7]; 
  assign s1_hazard_hi_hi_lo_2=|s1_mask_xwr[6]; 
  assign s1_hazard_hi_lo_hi_2=|s1_mask_xwr[5]; 
  assign s1_hazard_hi_lo_lo_2=|s1_mask_xwr[4]; 
  assign s1_hazard_lo_hi_hi_2=|s1_mask_xwr[3]; 
  assign s1_hazard_lo_hi_lo_2=|s1_mask_xwr[2]; 
  assign s1_hazard_lo_lo_hi_2=|s1_mask_xwr[1]; 
  assign s1_hazard_lo_lo_lo_2=|s1_mask_xwr[0]; 
  assign _s1_hazard_T_21={s1_hazard_hi_hi_hi_2,s1_hazard_hi_hi_lo_2,s1_hazard_hi_lo_hi_2,s1_hazard_hi_lo_lo_2,s1_hazard_lo_hi_hi_2,s1_hazard_lo_hi_lo_2,s1_hazard_lo_lo_hi_2,s1_hazard_lo_lo_lo_2}; 
  assign s1_hazard_hi_hi_hi_3=_s1_hazard_T_21[7]; 
  assign s1_hazard_hi_hi_lo_3=_s1_hazard_T_21[6]; 
  assign s1_hazard_hi_lo_hi_3=_s1_hazard_T_21[5]; 
  assign s1_hazard_hi_lo_lo_3=_s1_hazard_T_21[4]; 
  assign s1_hazard_lo_hi_hi_3=_s1_hazard_T_21[3]; 
  assign s1_hazard_lo_hi_lo_3=_s1_hazard_T_21[2]; 
  assign s1_hazard_lo_lo_hi_3=_s1_hazard_T_21[1]; 
  assign s1_hazard_lo_lo_lo_3=_s1_hazard_T_21[0]; 
  assign _s1_hazard_T_22={s1_hazard_hi_hi_hi_3,s1_hazard_hi_hi_lo_3,s1_hazard_hi_lo_hi_3,s1_hazard_hi_lo_lo_3,s1_hazard_lo_hi_hi_3,s1_hazard_lo_hi_lo_3,s1_hazard_lo_lo_hi_3,s1_hazard_lo_lo_lo_3}; 
  assign _s1_hazard_T_23=_s1_hazard_T_12&_s1_hazard_T_22; 
  assign _s1_hazard_T_24=|_s1_hazard_T_23; 
  assign _s1_hazard_T_25=pstore1_mask&s1_mask_xwr; 
  assign _s1_hazard_T_26=|_s1_hazard_T_25; 
  assign _s1_hazard_T_27=s1_write ? _s1_hazard_T_24:_s1_hazard_T_26; 
  assign _s1_hazard_T_28=_s1_hazard_T_2&_s1_hazard_T_27; 
  assign _s1_hazard_T_29=pstore1_valid_likely&_s1_hazard_T_28; 
  assign _s1_hazard_T_32=pstore2_addr[11:3]==s1_vaddr[11:3]; 
  assign s1_hazard_hi_hi_hi_4=|mask[7]; 
  assign s1_hazard_hi_hi_lo_4=|mask[6]; 
  assign s1_hazard_hi_lo_hi_4=|mask[5]; 
  assign s1_hazard_hi_lo_lo_4=|mask[4]; 
  assign s1_hazard_lo_hi_hi_4=|mask[3]; 
  assign s1_hazard_lo_hi_lo_4=|mask[2]; 
  assign s1_hazard_lo_lo_hi_4=|mask[1]; 
  assign s1_hazard_lo_lo_lo_4=|mask[0]; 
  assign _s1_hazard_T_41={s1_hazard_hi_hi_hi_4,s1_hazard_hi_hi_lo_4,s1_hazard_hi_lo_hi_4,s1_hazard_hi_lo_lo_4,s1_hazard_lo_hi_hi_4,s1_hazard_lo_hi_lo_4,s1_hazard_lo_lo_hi_4,s1_hazard_lo_lo_lo_4}; 
  assign s1_hazard_hi_hi_hi_5=_s1_hazard_T_41[7]; 
  assign s1_hazard_hi_hi_lo_5=_s1_hazard_T_41[6]; 
  assign s1_hazard_hi_lo_hi_5=_s1_hazard_T_41[5]; 
  assign s1_hazard_hi_lo_lo_5=_s1_hazard_T_41[4]; 
  assign s1_hazard_lo_hi_hi_5=_s1_hazard_T_41[3]; 
  assign s1_hazard_lo_hi_lo_5=_s1_hazard_T_41[2]; 
  assign s1_hazard_lo_lo_hi_5=_s1_hazard_T_41[1]; 
  assign s1_hazard_lo_lo_lo_5=_s1_hazard_T_41[0]; 
  assign _s1_hazard_T_42={s1_hazard_hi_hi_hi_5,s1_hazard_hi_hi_lo_5,s1_hazard_hi_lo_hi_5,s1_hazard_hi_lo_lo_5,s1_hazard_lo_hi_hi_5,s1_hazard_lo_hi_lo_5,s1_hazard_lo_lo_hi_5,s1_hazard_lo_lo_lo_5}; 
  assign _s1_hazard_T_53=_s1_hazard_T_42&_s1_hazard_T_22; 
  assign _s1_hazard_T_54=|_s1_hazard_T_53; 
  assign _s1_hazard_T_55=mask&s1_mask_xwr; 
  assign _s1_hazard_T_56=|_s1_hazard_T_55; 
  assign _s1_hazard_T_57=s1_write ? _s1_hazard_T_54:_s1_hazard_T_56; 
  assign _s1_hazard_T_58=_s1_hazard_T_32&_s1_hazard_T_57; 
  assign _s1_hazard_T_59=pstore2_valid&_s1_hazard_T_58; 
  assign s1_hazard=_s1_hazard_T_29|_s1_hazard_T_59; 
  assign s1_raw_hazard=s1_read&s1_hazard; 
  assign _T_262=s1_valid&s1_raw_hazard; 
  assign _s2_valid_no_xcpt_T={io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st,io_cpu_s2_xcpt_pf_ld,io_cpu_s2_xcpt_pf_st,io_cpu_s2_xcpt_ae_ld,io_cpu_s2_xcpt_ae_st}; 
  assign _s2_valid_no_xcpt_T_1=|_s2_valid_no_xcpt_T; 
  assign s2_valid_no_xcpt=s2_valid&~_s2_valid_no_xcpt_T_1; 
  assign s2_valid_masked=s2_valid_no_xcpt&s2_not_nacked_in_s1; 
  assign _s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1=s2_valid_masked&~s2_meta_error; 
  assign _c_cat_T_45=s2_req_cmd==5'h3; 
  assign _c_cat_T_46=s2_write|_c_cat_T_45; 
  assign _c_cat_T_47=s2_req_cmd==5'h6; 
  assign c_cat_lo=_c_cat_T_46|_c_cat_T_47; 
  assign _T_71={s2_write,c_cat_lo,s2_hit_state_state}; 
  assign _T_117=4'h3==_T_71; 
  assign _T_114=4'h2==_T_71; 
  assign _T_111=4'h1==_T_71; 
  assign _T_108=4'h7==_T_71; 
  assign _T_105=4'h6==_T_71; 
  assign _T_102=4'hf==_T_71; 
  assign _T_99=4'he==_T_71; 
  assign _T_96=4'h0==_T_71; 
  assign _T_93=4'h5==_T_71; 
  assign _T_90=4'h4==_T_71; 
  assign _T_87=4'hd==_T_71; 
  assign _T_84=4'hc==_T_71; 
  assign _T_103=_T_102|_T_99; 
  assign _T_106=_T_105|_T_103; 
  assign _T_109=_T_108|_T_106; 
  assign _T_112=_T_111|_T_109; 
  assign _T_115=_T_114|_T_112; 
  assign s2_hit=_T_117|_T_115; 
  assign s2_valid_hit_maybe_flush_pre_data_ecc_and_waw=_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1&s2_hit; 
  assign _s2_read_T=s2_req_cmd==5'h0; 
  assign _s2_read_T_2=_s2_read_T|_c_cat_T_47; 
  assign _s2_read_T_4=_s2_read_T_2|_s2_write_T_3; 
  assign s2_read=_s2_read_T_4|_s2_write_T_21; 
  assign s2_readwrite=s2_read|s2_write; 
  assign s2_valid_hit_pre_data_ecc_and_waw=s2_valid_hit_maybe_flush_pre_data_ecc_and_waw&s2_readwrite; 
  assign _T_86=_T_84 ? 2'h1:2'h0; 
  assign _T_89=_T_87 ? 2'h2:_T_86; 
  assign _T_92=_T_90 ? 2'h1:_T_89; 
  assign _T_95=_T_93 ? 2'h2:_T_92; 
  assign _T_98=_T_96 ? 2'h0:_T_95; 
  assign _T_101=_T_99 ? 2'h3:_T_98; 
  assign _T_104=_T_102 ? 2'h3:_T_101; 
  assign _T_107=_T_105 ? 2'h2:_T_104; 
  assign _T_110=_T_108 ? 2'h3:_T_107; 
  assign _T_113=_T_111 ? 2'h1:_T_110; 
  assign _T_116=_T_114 ? 2'h2:_T_113; 
  assign s2_grow_param=_T_117 ? 2'h3:_T_116; 
  assign _s2_update_meta_T=s2_hit_state_state==s2_grow_param; 
  assign s2_update_meta=~_s2_update_meta_T; 
  assign _T_241=s2_valid_hit_pre_data_ecc_and_waw&s2_update_meta; 
  assign _T_242=io_cpu_s2_nack|_T_241; 
  assign s1_readwrite=s1_read|s1_write; 
  assign _s1_flush_line_T=s1_req_cmd==5'h5; 
  assign s1_flush_line=_s1_flush_line_T&s1_req_size[0]; 
  assign _s1_cmd_uses_tlb_T=s1_readwrite|s1_flush_line; 
  assign _s1_cmd_uses_tlb_T_1=s1_req_cmd==5'h17; 
  assign s1_cmd_uses_tlb=_s1_cmd_uses_tlb_T|_s1_cmd_uses_tlb_T_1; 
  assign _T_13=s1_valid&s1_cmd_uses_tlb; 
  assign _T_14=_T_13&tlb_io_resp_miss; 
  assign _GEN_117=_T_242|_T_14; 
  assign _GEN_141=_T_262|_GEN_117; 
  assign _GEN_283=probeNack|_GEN_141; 
  assign s1_nack=s2_probe ? _GEN_283:_GEN_141; 
  assign s1_valid_not_nacked=s1_valid&~s1_nack; 
  assign s0_clk_en=metaArb_io_out_valid&~metaArb_io_out_bits_write; 
  assign s0_req_addr_hi=metaArb_io_out_bits_addr[39:6]; 
  assign s0_req_addr_lo=io_cpu_req_bits_addr[5:0]; 
  assign s0_req_addr={s0_req_addr_hi,s0_req_addr_lo}; 
  assign s0_req_phys=~metaArb_io_in_7_ready|io_cpu_req_bits_phys; 
  assign s1_sfence=s1_req_cmd==5'h14; 
  assign inWriteback=_T_308|_T_307; 
  assign _io_cpu_req_ready_T=release_state==4'h0; 
  assign _io_cpu_req_ready_T_2=_io_cpu_req_ready_T&~cached_grant_wait; 
  assign _io_cpu_req_ready_T_4=_io_cpu_req_ready_T_2&~s1_nack; 
  assign _s0_read_T=io_cpu_req_bits_cmd==5'h0; 
  assign _s0_read_T_1=io_cpu_req_bits_cmd==5'h6; 
  assign _s0_read_T_2=_s0_read_T|_s0_read_T_1; 
  assign _s0_read_T_3=io_cpu_req_bits_cmd==5'h7; 
  assign _s0_read_T_4=_s0_read_T_2|_s0_read_T_3; 
  assign _s0_read_T_5=io_cpu_req_bits_cmd==5'h4; 
  assign _s0_read_T_6=io_cpu_req_bits_cmd==5'h9; 
  assign _s0_read_T_7=io_cpu_req_bits_cmd==5'ha; 
  assign _s0_read_T_8=io_cpu_req_bits_cmd==5'hb; 
  assign _s0_read_T_9=_s0_read_T_5|_s0_read_T_6; 
  assign _s0_read_T_10=_s0_read_T_9|_s0_read_T_7; 
  assign _s0_read_T_11=_s0_read_T_10|_s0_read_T_8; 
  assign _s0_read_T_12=io_cpu_req_bits_cmd==5'h8; 
  assign _s0_read_T_13=io_cpu_req_bits_cmd==5'hc; 
  assign _s0_read_T_14=io_cpu_req_bits_cmd==5'hd; 
  assign _s0_read_T_15=io_cpu_req_bits_cmd==5'he; 
  assign _s0_read_T_16=io_cpu_req_bits_cmd==5'hf; 
  assign _s0_read_T_17=_s0_read_T_12|_s0_read_T_13; 
  assign _s0_read_T_18=_s0_read_T_17|_s0_read_T_14; 
  assign _s0_read_T_19=_s0_read_T_18|_s0_read_T_15; 
  assign _s0_read_T_20=_s0_read_T_19|_s0_read_T_16; 
  assign _s0_read_T_21=_s0_read_T_11|_s0_read_T_20; 
  assign s0_read=_s0_read_T_4|_s0_read_T_21; 
  assign _dataArb_io_in_3_valid_res_T=io_cpu_req_bits_cmd==5'h1; 
  assign _dataArb_io_in_3_valid_res_T_1=io_cpu_req_bits_cmd==5'h3; 
  assign _dataArb_io_in_3_valid_res_T_2=_dataArb_io_in_3_valid_res_T|_dataArb_io_in_3_valid_res_T_1; 
  assign res=~_dataArb_io_in_3_valid_res_T_2; 
  assign _dataArb_io_in_3_valid_T_24=io_cpu_req_bits_cmd==5'h11; 
  assign _dataArb_io_in_3_valid_T_25=_dataArb_io_in_3_valid_res_T|_dataArb_io_in_3_valid_T_24; 
  assign _dataArb_io_in_3_valid_T_27=_dataArb_io_in_3_valid_T_25|_s0_read_T_3; 
  assign _dataArb_io_in_3_valid_T_45=_dataArb_io_in_3_valid_T_27|_s0_read_T_21; 
  assign _dataArb_io_in_3_valid_T_49=_dataArb_io_in_3_valid_T_45&_dataArb_io_in_3_valid_T_24; 
  assign _dataArb_io_in_3_valid_T_50=s0_read|_dataArb_io_in_3_valid_T_49; 
  assign _dataArb_io_in_3_valid_T_52=~_dataArb_io_in_3_valid_T_50|res; 
  assign _dataArb_io_in_3_valid_T_54=_dataArb_io_in_3_valid_T_52|reset; 
  assign _dataArb_io_in_3_valid_T_56=io_cpu_req_valid&res; 
  assign dataArb_io_in_3_bits_addr_hi=io_cpu_req_bits_addr[39:12]; 
  assign dataArb_io_in_3_bits_addr_lo=io_cpu_req_bits_addr[11:0]; 
  assign _dataArb_io_in_3_bits_addr_T={dataArb_io_in_3_bits_addr_hi,dataArb_io_in_3_bits_addr_lo}; 
  assign _T_4=~dataArb_io_in_3_ready&s0_read; 
  assign _GEN_28=_T_4 ? 1'h0:_io_cpu_req_ready_T_4; 
  assign _s1_did_read_T_51=io_cpu_req_valid&_dataArb_io_in_3_valid_T_50; 
  assign _s1_did_read_T_52=dataArb_io_in_3_ready&_s1_did_read_T_51; 
  assign _GEN_31=metaArb_io_in_7_ready ? _GEN_28:1'h0; 
  assign _T_8=~tlb_io_req_ready&~tlb_io_ptw_resp_valid; 
  assign _T_10=_T_8&~io_cpu_req_bits_phys; 
  assign _GEN_32=_T_10 ? 1'h0:_GEN_31; 
  assign s1_paddr_hi=tlb_io_resp_paddr[31:12]; 
  assign s1_paddr={s1_paddr_hi,s1_vaddr_lo}; 
  assign _WIRE_2=tag_array_0_s1_meta_data; 
  assign s1_meta_uncorrected_0_tag=_WIRE_2[19:0]; 
  assign s1_meta_uncorrected_0_coh_state=_WIRE_2[21:20]; 
  assign _WIRE_3=tag_array_1_s1_meta_data; 
  assign s1_meta_uncorrected_1_tag=_WIRE_3[19:0]; 
  assign s1_meta_uncorrected_1_coh_state=_WIRE_3[21:20]; 
  assign _WIRE_4=tag_array_2_s1_meta_data; 
  assign s1_meta_uncorrected_2_tag=_WIRE_4[19:0]; 
  assign s1_meta_uncorrected_2_coh_state=_WIRE_4[21:20]; 
  assign _WIRE_5=tag_array_3_s1_meta_data; 
  assign s1_meta_uncorrected_3_tag=_WIRE_5[19:0]; 
  assign s1_meta_uncorrected_3_coh_state=_WIRE_5[21:20]; 
  assign s1_tag=s1_paddr[31:12]; 
  assign _T_32=s1_meta_uncorrected_0_coh_state>2'h0; 
  assign _T_33=s1_meta_uncorrected_0_tag==s1_tag; 
  assign lo_lo=_T_32&_T_33; 
  assign _T_34=s1_meta_uncorrected_1_coh_state>2'h0; 
  assign _T_35=s1_meta_uncorrected_1_tag==s1_tag; 
  assign lo_hi=_T_34&_T_35; 
  assign _T_36=s1_meta_uncorrected_2_coh_state>2'h0; 
  assign _T_37=s1_meta_uncorrected_2_tag==s1_tag; 
  assign hi_lo=_T_36&_T_37; 
  assign _T_38=s1_meta_uncorrected_3_coh_state>2'h0; 
  assign _T_39=s1_meta_uncorrected_3_tag==s1_tag; 
  assign hi_hi=_T_38&_T_39; 
  assign s1_meta_hit_way={hi_hi,hi_lo,lo_hi,lo_lo}; 
  assign _T_42=_T_33&~s1_flush_valid; 
  assign _T_43=_T_42 ? s1_meta_uncorrected_0_coh_state:2'h0; 
  assign _T_46=_T_35&~s1_flush_valid; 
  assign _T_47=_T_46 ? s1_meta_uncorrected_1_coh_state:2'h0; 
  assign _T_50=_T_37&~s1_flush_valid; 
  assign _T_51=_T_50 ? s1_meta_uncorrected_2_coh_state:2'h0; 
  assign _T_54=_T_39&~s1_flush_valid; 
  assign _T_55=_T_54 ? s1_meta_uncorrected_3_coh_state:2'h0; 
  assign _T_56=_T_43|_T_47; 
  assign _T_57=_T_56|_T_51; 
  assign s1_meta_hit_state_state=_T_57|_T_55; 
  assign s2_hit_valid=s2_hit_state_state>2'h0; 
  assign s2_victim_way=4'h1<<s2_victim_way_r; 
  assign s2_victim_or_hit_way=s2_hit_valid ? s2_hit_way:s2_victim_way; 
  assign releaseWay=_T_312 ? s2_victim_or_hit_way:s2_probe_way; 
  assign s1_data_way_x35=inWriteback ? releaseWay:s1_meta_hit_way; 
  assign tl_d_data_encoded_lo_lo_lo=auto_out_d_bits_data[7:0]; 
  assign tl_d_data_encoded_lo_lo_hi=auto_out_d_bits_data[15:8]; 
  assign tl_d_data_encoded_lo_hi_lo=auto_out_d_bits_data[23:16]; 
  assign tl_d_data_encoded_lo_hi_hi=auto_out_d_bits_data[31:24]; 
  assign tl_d_data_encoded_hi_lo_lo=auto_out_d_bits_data[39:32]; 
  assign tl_d_data_encoded_hi_lo_hi=auto_out_d_bits_data[47:40]; 
  assign tl_d_data_encoded_hi_hi_lo=auto_out_d_bits_data[55:48]; 
  assign tl_d_data_encoded_hi_hi_hi=auto_out_d_bits_data[63:56]; 
  assign tl_d_data_encoded_lo={tl_d_data_encoded_lo_hi_hi,tl_d_data_encoded_lo_hi_lo,tl_d_data_encoded_lo_lo_hi,tl_d_data_encoded_lo_lo_lo}; 
  assign tl_d_data_encoded_hi={tl_d_data_encoded_hi_hi_hi,tl_d_data_encoded_hi_hi_lo,tl_d_data_encoded_hi_lo_hi,tl_d_data_encoded_hi_lo_lo}; 
  assign _tl_d_data_encoded_T={tl_d_data_encoded_hi_hi_hi,tl_d_data_encoded_hi_hi_lo,tl_d_data_encoded_hi_lo_hi,tl_d_data_encoded_hi_lo_lo,tl_d_data_encoded_lo_hi_hi,tl_d_data_encoded_lo_hi_lo,tl_d_data_encoded_lo_lo_hi,tl_d_data_encoded_lo_lo_lo}; 
  assign _T_61=s1_valid_masked&_s1_write_T_1; 
  assign _T_65=&8'hff; 
  assign _T_66=~_T_61|_T_65; 
  assign _T_68=_T_66|reset; 
  assign s2_valid_x37=s1_valid_masked&~s1_sfence; 
  assign _s2_cmd_flush_all_T=s2_req_cmd==5'h5; 
  assign s2_cmd_flush_line=_s2_cmd_flush_all_T&s2_req_size[0]; 
  assign _T_70=s1_valid_not_nacked|s1_flush_valid; 
  assign _s2_pma_T_cacheable=tlb_io_resp_cacheable; 
  assign s2_vaddr_hi=s2_vaddr_r[39:12]; 
  assign s2_vaddr_lo=s2_req_addr[11:0]; 
  assign s2_vaddr={s2_vaddr_hi,s2_vaddr_lo}; 
  assign s1_meta_clk_en=_T_70|s1_probe; 
  assign s2_meta_corrected_0_tag=s2_meta_corrected_r[19:0]; 
  assign s2_meta_corrected_0_coh_state=s2_meta_corrected_r[21:20]; 
  assign s2_meta_corrected_1_tag=s2_meta_corrected_r_1[19:0]; 
  assign s2_meta_corrected_1_coh_state=s2_meta_corrected_r_1[21:20]; 
  assign s2_meta_corrected_2_tag=s2_meta_corrected_r_2[19:0]; 
  assign s2_meta_corrected_2_coh_state=s2_meta_corrected_r_2[21:20]; 
  assign s2_meta_corrected_3_tag=s2_meta_corrected_r_3[19:0]; 
  assign s2_meta_corrected_3_coh_state=s2_meta_corrected_r_3[21:20]; 
  assign s2_flush_valid=s2_flush_valid_pre_tag_ecc&~s2_meta_error; 
  assign _s2_data_en_T=s1_valid|inWriteback; 
  assign en=_s2_data_en_T|io_cpu_replay_next; 
  assign _s2_data_word_en_T=s1_did_read&s1_read_mask; 
  assign word_en=inWriteback|_s2_data_word_en_T; 
  assign s1_all_data_ways_0=data_io_resp_0; 
  assign s1_all_data_ways_1=data_io_resp_1; 
  assign s1_all_data_ways_2=data_io_resp_2; 
  assign s1_all_data_ways_3=data_io_resp_3; 
  assign s1_word_en=io_cpu_replay_next ? 1'h1:word_en; 
  assign grantIsUncachedData=auto_out_d_bits_opcode==3'h1; 
  assign _T_293=blockUncachedGrant|s1_valid; 
  assign _T_294=grantIsUncachedData&_T_293; 
  assign grantIsRefill=auto_out_d_bits_opcode==3'h5; 
  assign _T_292=grantIsRefill&~dataArb_io_in_1_ready; 
  assign _grantIsCached_T=auto_out_d_bits_opcode==3'h4; 
  assign grantIsCached=_grantIsCached_T|grantIsRefill; 
  assign d_first=counter==9'h0; 
  assign _bundleOut_0_d_ready_T_1=~d_first|auto_out_e_ready; 
  assign canAcceptCachedGrant=~_T_312; 
  assign _bundleOut_0_d_ready_T_2=_bundleOut_0_d_ready_T_1&canAcceptCachedGrant; 
  assign _bundleOut_0_d_ready_T_3=grantIsCached ? _bundleOut_0_d_ready_T_2:1'h1; 
  assign _GEN_233=_T_292 ? 1'h0:_bundleOut_0_d_ready_T_3; 
  assign tl_out__d_ready=_T_294 ? 1'h0:_GEN_233; 
  assign _T_271=tl_out__d_ready&auto_out_d_valid; 
  assign _T_267=auto_out_d_bits_opcode==3'h0; 
  assign _T_269=grantIsUncachedData|_T_267; 
  assign _T_268=auto_out_d_bits_opcode==3'h2; 
  assign grantIsUncached=_T_269|_T_268; 
  assign _GEN_189=grantIsUncachedData ? 5'h10:{1'b0,s1_data_way_x35}; 
  assign _GEN_198=grantIsUncached ? _GEN_189:{1'b0,s1_data_way_x35}; 
  assign _GEN_211=grantIsCached ? {1'b0,s1_data_way_x35}:_GEN_198; 
  assign s1_data_way=_T_271 ? _GEN_211:{1'b0,s1_data_way_x35}; 
  assign _s2_data_T_1=s1_word_en ? s1_data_way:5'h0; 
  assign _s2_data_T_7=_s2_data_T_1[0] ? s1_all_data_ways_0:64'h0; 
  assign _s2_data_T_8=_s2_data_T_1[1] ? s1_all_data_ways_1:64'h0; 
  assign _s2_data_T_9=_s2_data_T_1[2] ? s1_all_data_ways_2:64'h0; 
  assign _s2_data_T_10=_s2_data_T_1[3] ? s1_all_data_ways_3:64'h0; 
  assign _s2_data_T_11=_s2_data_T_1[4] ? _tl_d_data_encoded_T:64'h0; 
  assign _s2_data_T_12=_s2_data_T_7|_s2_data_T_8; 
  assign _s2_data_T_13=_s2_data_T_12|_s2_data_T_9; 
  assign _s2_data_T_14=_s2_data_T_13|_s2_data_T_10; 
  assign _s2_data_T_15=_s2_data_T_14|_s2_data_T_11; 
  assign s2_data_uncorrected_lo_lo_lo=s2_data[7:0]; 
  assign s2_data_uncorrected_lo_lo_hi=s2_data[15:8]; 
  assign s2_data_uncorrected_lo_hi_lo=s2_data[23:16]; 
  assign s2_data_uncorrected_lo_hi_hi=s2_data[31:24]; 
  assign s2_data_uncorrected_hi_lo_lo=s2_data[39:32]; 
  assign s2_data_uncorrected_hi_lo_hi=s2_data[47:40]; 
  assign s2_data_uncorrected_hi_hi_lo=s2_data[55:48]; 
  assign s2_data_uncorrected_hi_hi_hi=s2_data[63:56]; 
  assign s2_data_corrected_lo={s2_data_uncorrected_lo_hi_hi,s2_data_uncorrected_lo_hi_lo,s2_data_uncorrected_lo_lo_hi,s2_data_uncorrected_lo_lo_lo}; 
  assign s2_data_corrected_hi={s2_data_uncorrected_hi_hi_hi,s2_data_uncorrected_hi_hi_lo,s2_data_uncorrected_hi_lo_hi,s2_data_uncorrected_hi_lo_lo}; 
  assign s2_data_corrected={s2_data_uncorrected_hi_hi_hi,s2_data_uncorrected_hi_hi_lo,s2_data_uncorrected_hi_lo_hi,s2_data_uncorrected_hi_lo_lo,s2_data_uncorrected_lo_hi_hi,s2_data_uncorrected_lo_hi_lo,s2_data_uncorrected_lo_lo_hi,s2_data_uncorrected_lo_lo_lo}; 
  assign s2_valid_flush_line=s2_valid_hit_maybe_flush_pre_data_ecc_and_waw&s2_cmd_flush_line; 
  assign _s2_valid_miss_T=s2_valid_masked&s2_readwrite; 
  assign _s2_valid_miss_T_2=_s2_valid_miss_T&~s2_meta_error; 
  assign s2_valid_miss=_s2_valid_miss_T_2&~s2_hit; 
  assign s2_uncached=~s2_pma_cacheable; 
  assign _s2_valid_cached_miss_T_1=s2_valid_miss&~s2_uncached; 
  assign _s2_valid_cached_miss_T_2=|uncachedInFlight_0; 
  assign s2_valid_cached_miss=_s2_valid_cached_miss_T_1&~_s2_valid_cached_miss_T_2; 
  assign _s2_want_victimize_T=s2_valid_cached_miss|s2_valid_flush_line; 
  assign s2_want_victimize=_s2_want_victimize_T|s2_flush_valid; 
  assign _s2_valid_uncached_pending_T=s2_valid_miss&s2_uncached; 
  assign _s2_valid_uncached_pending_T_1=&uncachedInFlight_0; 
  assign s2_valid_uncached_pending=_s2_valid_uncached_pending_T&~_s2_valid_uncached_pending_T_1; 
  assign s1_victim_way=lfsr[1:0]; 
  assign _s2_victim_tag_T_6=s2_victim_way[0] ? s2_meta_corrected_0_tag:20'h0; 
  assign _s2_victim_tag_T_7=s2_victim_way[1] ? s2_meta_corrected_1_tag:20'h0; 
  assign _s2_victim_tag_T_8=s2_victim_way[2] ? s2_meta_corrected_2_tag:20'h0; 
  assign _s2_victim_tag_T_9=s2_victim_way[3] ? s2_meta_corrected_3_tag:20'h0; 
  assign _s2_victim_tag_T_10=_s2_victim_tag_T_6|_s2_victim_tag_T_7; 
  assign _s2_victim_tag_T_11=_s2_victim_tag_T_10|_s2_victim_tag_T_8; 
  assign _s2_victim_tag_T_12=_s2_victim_tag_T_11|_s2_victim_tag_T_9; 
  assign _s2_victim_tag_T_13=s2_victim_way[0] ? s2_meta_corrected_0_coh_state:2'h0; 
  assign _s2_victim_tag_T_14=s2_victim_way[1] ? s2_meta_corrected_1_coh_state:2'h0; 
  assign _s2_victim_tag_T_15=s2_victim_way[2] ? s2_meta_corrected_2_coh_state:2'h0; 
  assign _s2_victim_tag_T_16=s2_victim_way[3] ? s2_meta_corrected_3_coh_state:2'h0; 
  assign _s2_victim_tag_T_17=_s2_victim_tag_T_13|_s2_victim_tag_T_14; 
  assign _s2_victim_tag_T_18=_s2_victim_tag_T_17|_s2_victim_tag_T_15; 
  assign _s2_victim_tag_T_19=_s2_victim_tag_T_18|_s2_victim_tag_T_16; 
  assign s2_victim_tag=s2_valid_flush_line ? s2_req_addr[31:12]:_s2_victim_tag_T_12; 
  assign s2_victim_state_state=s2_hit_valid ? s2_hit_state_state:_s2_victim_tag_T_19; 
  assign _T_133=_T_131 ? 3'h5:3'h0; 
  assign _T_137=_T_135 ? 3'h2:_T_133; 
  assign _T_141=_T_139 ? 3'h1:_T_137; 
  assign _T_145=_T_143 ? 3'h1:_T_141; 
  assign _T_149=_T_147 ? 3'h5:_T_145; 
  assign _T_153=_T_151 ? 3'h4:_T_149; 
  assign _T_154=_T_151 ? 2'h1:2'h0; 
  assign _T_157=_T_155 ? 3'h0:_T_153; 
  assign _T_158=_T_155 ? 2'h1:_T_154; 
  assign _T_161=_T_159 ? 3'h0:_T_157; 
  assign _T_162=_T_159 ? 2'h1:_T_158; 
  assign _T_165=_T_163 ? 3'h5:_T_161; 
  assign _T_166=_T_163 ? 2'h0:_T_162; 
  assign _T_169=_T_167 ? 3'h4:_T_165; 
  assign _T_170=_T_167 ? 2'h1:_T_166; 
  assign _T_173=_T_171 ? 3'h3:_T_169; 
  assign _T_174=_T_171 ? 2'h2:_T_170; 
  assign s2_report_param=_T_175 ? 3'h3:_T_173; 
  assign probeNewCoh_state=_T_175 ? 2'h2:_T_174; 
  assign _T_182={2'h2,s2_victim_state_state}; 
  assign _T_195=4'h8==_T_182; 
  assign _T_197=_T_195 ? 3'h5:3'h0; 
  assign _T_199=4'h9==_T_182; 
  assign _T_201=_T_199 ? 3'h2:_T_197; 
  assign _T_203=4'ha==_T_182; 
  assign _T_205=_T_203 ? 3'h1:_T_201; 
  assign _T_207=4'hb==_T_182; 
  assign _T_209=_T_207 ? 3'h1:_T_205; 
  assign _T_211=4'h4==_T_182; 
  assign _T_212=_T_211 ? 1'h0:_T_207; 
  assign _T_213=_T_211 ? 3'h5:_T_209; 
  assign _T_215=4'h5==_T_182; 
  assign _T_216=_T_215 ? 1'h0:_T_212; 
  assign _T_217=_T_215 ? 3'h4:_T_213; 
  assign _T_218=_T_215 ? 2'h1:2'h0; 
  assign _T_219=4'h6==_T_182; 
  assign _T_220=_T_219 ? 1'h0:_T_216; 
  assign _T_221=_T_219 ? 3'h0:_T_217; 
  assign _T_222=_T_219 ? 2'h1:_T_218; 
  assign _T_223=4'h7==_T_182; 
  assign _T_224=_T_223|_T_220; 
  assign _T_225=_T_223 ? 3'h0:_T_221; 
  assign _T_226=_T_223 ? 2'h1:_T_222; 
  assign _T_227=4'h0==_T_182; 
  assign _T_228=_T_227 ? 1'h0:_T_224; 
  assign _T_229=_T_227 ? 3'h5:_T_225; 
  assign _T_230=_T_227 ? 2'h0:_T_226; 
  assign _T_231=4'h1==_T_182; 
  assign _T_232=_T_231 ? 1'h0:_T_228; 
  assign _T_233=_T_231 ? 3'h4:_T_229; 
  assign _T_234=_T_231 ? 2'h1:_T_230; 
  assign _T_235=4'h2==_T_182; 
  assign _T_236=_T_235 ? 1'h0:_T_232; 
  assign _T_237=_T_235 ? 3'h3:_T_233; 
  assign _T_238=_T_235 ? 2'h2:_T_234; 
  assign _T_239=4'h3==_T_182; 
  assign s2_victim_dirty=_T_239|_T_236; 
  assign s2_shrink_param=_T_239 ? 3'h3:_T_237; 
  assign voluntaryNewCoh_state=_T_239 ? 2'h2:_T_238; 
  assign s2_dont_nack_uncached=s2_valid_uncached_pending&auto_out_a_ready; 
  assign _s2_dont_nack_misc_T_10=s2_req_cmd==5'h17; 
  assign s2_dont_nack_misc=_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw_T_1&_s2_dont_nack_misc_T_10; 
  assign _io_cpu_s2_nack_T_1=s2_valid_no_xcpt&~s2_dont_nack_uncached; 
  assign _io_cpu_s2_nack_T_3=_io_cpu_s2_nack_T_1&~s2_dont_nack_misc; 
  assign _metaArb_io_in_1_valid_T=s2_valid_masked|s2_flush_valid_pre_tag_ecc; 
  assign _metaArb_io_in_1_valid_T_1=_metaArb_io_in_1_valid_T|s2_probe; 
  assign metaArb_io_in_1_bits_addr_lo={metaArb_io_in_1_bits_idx,6'h0}; 
  assign new_meta_coh_state=s2_meta_error ? 2'h0:s2_meta_corrected_3_coh_state; 
  assign metaArb_io_in_2_bits_addr_lo=s2_vaddr[11:0]; 
  assign metaArb_io_in_2_bits_data_meta_tag=s2_req_addr[31:12]; 
  assign _lrscBackingOff_T=lrscCount>7'h0; 
  assign lrscBackingOff=_lrscBackingOff_T&~lrscValid; 
  assign lrscAddrMatch=lrscAddr==s2_req_addr[39:6]; 
  assign _s2_sc_fail_T=lrscValid&lrscAddrMatch; 
  assign s2_sc_fail=_s2_write_T_3&~_s2_sc_fail_T; 
  assign _T_243=s2_valid_hit_pre_data_ecc_and_waw&_c_cat_T_47; 
  assign _T_245=_T_243&~cached_grant_wait; 
  assign _T_246=_T_245|s2_valid_cached_miss; 
  assign _lrscCount_T_2=lrscCount-7'h1; 
  assign _T_250=s2_valid_masked&lrscValid; 
  assign _pstore1_cmd_T=s1_valid_not_nacked&s1_write; 
  assign _pstore1_rmw_T_49=s1_write&_s1_write_T_1; 
  assign _pstore1_rmw_T_50=s1_read|_pstore1_rmw_T_49; 
  assign _pstore1_merge_T=s2_valid_hit_pre_data_ecc_and_waw&s2_write; 
  assign _pstore1_merge_T_2=_pstore1_merge_T&~s2_sc_fail; 
  assign pstore_drain_opportunistic=~_dataArb_io_in_3_valid_T_56; 
  assign pstore_drain_on_miss=releaseInFlight|pstore_drain_on_miss_REG; 
  assign pstore1_valid=_pstore1_merge_T_2|pstore1_held; 
  assign _pstore_drain_structural_T=pstore1_valid_likely&pstore2_valid; 
  assign _pstore_drain_structural_T_1=s1_valid&s1_write; 
  assign _pstore_drain_structural_T_2=_pstore_drain_structural_T_1|pstore1_rmw_r; 
  assign pstore_drain_structural=_pstore_drain_structural_T&_pstore_drain_structural_T_2; 
  assign _T_254=_pstore1_merge_T|pstore1_held; 
  assign _T_255=_T_254==pstore1_valid; 
  assign _T_256=pstore1_rmw_r|_T_255; 
  assign _T_258=_T_256|reset; 
  assign _pstore_drain_T_7=_T_254&~pstore1_rmw_r; 
  assign _pstore_drain_T_8=_pstore_drain_T_7|pstore2_valid; 
  assign _pstore_drain_T_9=pstore_drain_opportunistic|pstore_drain_on_miss; 
  assign _pstore_drain_T_10=_pstore_drain_T_8&_pstore_drain_T_9; 
  assign pstore_drain=pstore_drain_structural|_pstore_drain_T_10; 
  assign _pstore1_held_T_8=pstore1_valid&pstore2_valid; 
  assign _pstore1_held_T_10=_pstore1_held_T_8&~pstore_drain; 
  assign _advance_pstore1_T_1=pstore2_valid==pstore_drain; 
  assign advance_pstore1=pstore1_valid&_advance_pstore1_T_1; 
  assign _pstore2_valid_T_1=pstore2_valid&~pstore_drain; 
  assign _pstore2_valid_T_2=_pstore2_valid_T_1|advance_pstore1; 
  assign pstore1_storegen_data=amoalu_io_out; 
  assign pstore2_storegen_data={pstore2_storegen_data_hi_hi_hi,pstore2_storegen_data_hi_hi_lo,pstore2_storegen_data_hi_lo_hi,pstore2_storegen_data_hi_lo_lo,pstore2_storegen_data_lo_hi_hi,pstore2_storegen_data_lo_hi_lo,pstore2_storegen_data_lo_lo_hi,pstore2_storegen_data_lo_lo_lo}; 
  assign _dataArb_io_in_0_bits_addr_T=pstore2_valid ? pstore2_addr:pstore1_addr; 
  assign _dataArb_io_in_0_bits_wdata_T=pstore2_valid ? pstore2_storegen_data:pstore1_data; 
  assign dataArb_io_in_0_bits_wdata_lo_lo_lo=_dataArb_io_in_0_bits_wdata_T[7:0]; 
  assign dataArb_io_in_0_bits_wdata_lo_lo_hi=_dataArb_io_in_0_bits_wdata_T[15:8]; 
  assign dataArb_io_in_0_bits_wdata_lo_hi_lo=_dataArb_io_in_0_bits_wdata_T[23:16]; 
  assign dataArb_io_in_0_bits_wdata_lo_hi_hi=_dataArb_io_in_0_bits_wdata_T[31:24]; 
  assign dataArb_io_in_0_bits_wdata_hi_lo_lo=_dataArb_io_in_0_bits_wdata_T[39:32]; 
  assign dataArb_io_in_0_bits_wdata_hi_lo_hi=_dataArb_io_in_0_bits_wdata_T[47:40]; 
  assign dataArb_io_in_0_bits_wdata_hi_hi_lo=_dataArb_io_in_0_bits_wdata_T[55:48]; 
  assign dataArb_io_in_0_bits_wdata_hi_hi_hi=_dataArb_io_in_0_bits_wdata_T[63:56]; 
  assign dataArb_io_in_0_bits_wdata_lo={dataArb_io_in_0_bits_wdata_lo_hi_hi,dataArb_io_in_0_bits_wdata_lo_hi_lo,dataArb_io_in_0_bits_wdata_lo_lo_hi,dataArb_io_in_0_bits_wdata_lo_lo_lo}; 
  assign dataArb_io_in_0_bits_wdata_hi={dataArb_io_in_0_bits_wdata_hi_hi_hi,dataArb_io_in_0_bits_wdata_hi_hi_lo,dataArb_io_in_0_bits_wdata_hi_lo_hi,dataArb_io_in_0_bits_wdata_hi_lo_lo}; 
  assign _dataArb_io_in_0_bits_eccMask_T=pstore2_valid ? mask:pstore1_mask; 
  assign dataArb_io_in_0_bits_eccMask_lo_lo_lo=|_dataArb_io_in_0_bits_eccMask_T[0]; 
  assign dataArb_io_in_0_bits_eccMask_lo_lo_hi=|_dataArb_io_in_0_bits_eccMask_T[1]; 
  assign dataArb_io_in_0_bits_eccMask_lo_hi_lo=|_dataArb_io_in_0_bits_eccMask_T[2]; 
  assign dataArb_io_in_0_bits_eccMask_lo_hi_hi=|_dataArb_io_in_0_bits_eccMask_T[3]; 
  assign dataArb_io_in_0_bits_eccMask_hi_lo_lo=|_dataArb_io_in_0_bits_eccMask_T[4]; 
  assign dataArb_io_in_0_bits_eccMask_hi_lo_hi=|_dataArb_io_in_0_bits_eccMask_T[5]; 
  assign dataArb_io_in_0_bits_eccMask_hi_hi_lo=|_dataArb_io_in_0_bits_eccMask_T[6]; 
  assign dataArb_io_in_0_bits_eccMask_hi_hi_hi=|_dataArb_io_in_0_bits_eccMask_T[7]; 
  assign dataArb_io_in_0_bits_eccMask_lo={dataArb_io_in_0_bits_eccMask_lo_hi_hi,dataArb_io_in_0_bits_eccMask_lo_hi_lo,dataArb_io_in_0_bits_eccMask_lo_lo_hi,dataArb_io_in_0_bits_eccMask_lo_lo_lo}; 
  assign dataArb_io_in_0_bits_eccMask_hi={dataArb_io_in_0_bits_eccMask_hi_hi_hi,dataArb_io_in_0_bits_eccMask_hi_hi_lo,dataArb_io_in_0_bits_eccMask_hi_lo_hi,dataArb_io_in_0_bits_eccMask_hi_lo_lo}; 
  assign _a_source_T_1={~uncachedInFlight_0,1'h0}; 
  assign a_source=_a_source_T_1[0] ? 1'h0:1'h1; 
  assign acquire_address={s2_req_addr[39:6],6'h0}; 
  assign a_mask={15'b0,pstore1_mask}; 
  assign _get_a_mask_sizeOH_T={1'b0,s2_req_size}; 
  assign get_a_mask_sizeOH_shiftAmount=_get_a_mask_sizeOH_T[1:0]; 
  assign _get_a_mask_sizeOH_T_1=4'h1<<get_a_mask_sizeOH_shiftAmount; 
  assign get_a_mask_sizeOH=_get_a_mask_sizeOH_T_1[2:0]|3'h1; 
  assign _get_a_mask_T=s2_req_size>=2'h3; 
  assign get_a_mask_size=get_a_mask_sizeOH[2]; 
  assign get_a_mask_bit=s2_req_addr[2]; 
  assign get_a_mask_nbit=~get_a_mask_bit; 
  assign _get_a_mask_acc_T=get_a_mask_size&get_a_mask_nbit; 
  assign get_a_mask_acc=_get_a_mask_T|_get_a_mask_acc_T; 
  assign _get_a_mask_acc_T_1=get_a_mask_size&get_a_mask_bit; 
  assign get_a_mask_acc_1=_get_a_mask_T|_get_a_mask_acc_T_1; 
  assign get_a_mask_size_1=get_a_mask_sizeOH[1]; 
  assign get_a_mask_bit_1=s2_req_addr[1]; 
  assign get_a_mask_nbit_1=~get_a_mask_bit_1; 
  assign get_a_mask_eq_2=get_a_mask_nbit&get_a_mask_nbit_1; 
  assign _get_a_mask_acc_T_2=get_a_mask_size_1&get_a_mask_eq_2; 
  assign get_a_mask_acc_2=get_a_mask_acc|_get_a_mask_acc_T_2; 
  assign get_a_mask_eq_3=get_a_mask_nbit&get_a_mask_bit_1; 
  assign _get_a_mask_acc_T_3=get_a_mask_size_1&get_a_mask_eq_3; 
  assign get_a_mask_acc_3=get_a_mask_acc|_get_a_mask_acc_T_3; 
  assign get_a_mask_eq_4=get_a_mask_bit&get_a_mask_nbit_1; 
  assign _get_a_mask_acc_T_4=get_a_mask_size_1&get_a_mask_eq_4; 
  assign get_a_mask_acc_4=get_a_mask_acc_1|_get_a_mask_acc_T_4; 
  assign get_a_mask_eq_5=get_a_mask_bit&get_a_mask_bit_1; 
  assign _get_a_mask_acc_T_5=get_a_mask_size_1&get_a_mask_eq_5; 
  assign get_a_mask_acc_5=get_a_mask_acc_1|_get_a_mask_acc_T_5; 
  assign get_a_mask_size_2=get_a_mask_sizeOH[0]; 
  assign get_a_mask_bit_2=s2_req_addr[0]; 
  assign get_a_mask_nbit_2=~get_a_mask_bit_2; 
  assign get_a_mask_eq_6=get_a_mask_eq_2&get_a_mask_nbit_2; 
  assign _get_a_mask_acc_T_6=get_a_mask_size_2&get_a_mask_eq_6; 
  assign get_a_mask_lo_lo_lo=get_a_mask_acc_2|_get_a_mask_acc_T_6; 
  assign get_a_mask_eq_7=get_a_mask_eq_2&get_a_mask_bit_2; 
  assign _get_a_mask_acc_T_7=get_a_mask_size_2&get_a_mask_eq_7; 
  assign get_a_mask_lo_lo_hi=get_a_mask_acc_2|_get_a_mask_acc_T_7; 
  assign get_a_mask_eq_8=get_a_mask_eq_3&get_a_mask_nbit_2; 
  assign _get_a_mask_acc_T_8=get_a_mask_size_2&get_a_mask_eq_8; 
  assign get_a_mask_lo_hi_lo=get_a_mask_acc_3|_get_a_mask_acc_T_8; 
  assign get_a_mask_eq_9=get_a_mask_eq_3&get_a_mask_bit_2; 
  assign _get_a_mask_acc_T_9=get_a_mask_size_2&get_a_mask_eq_9; 
  assign get_a_mask_lo_hi_hi=get_a_mask_acc_3|_get_a_mask_acc_T_9; 
  assign get_a_mask_eq_10=get_a_mask_eq_4&get_a_mask_nbit_2; 
  assign _get_a_mask_acc_T_10=get_a_mask_size_2&get_a_mask_eq_10; 
  assign get_a_mask_hi_lo_lo=get_a_mask_acc_4|_get_a_mask_acc_T_10; 
  assign get_a_mask_eq_11=get_a_mask_eq_4&get_a_mask_bit_2; 
  assign _get_a_mask_acc_T_11=get_a_mask_size_2&get_a_mask_eq_11; 
  assign get_a_mask_hi_lo_hi=get_a_mask_acc_4|_get_a_mask_acc_T_11; 
  assign get_a_mask_eq_12=get_a_mask_eq_5&get_a_mask_nbit_2; 
  assign _get_a_mask_acc_T_12=get_a_mask_size_2&get_a_mask_eq_12; 
  assign get_a_mask_hi_hi_lo=get_a_mask_acc_5|_get_a_mask_acc_T_12; 
  assign get_a_mask_eq_13=get_a_mask_eq_5&get_a_mask_bit_2; 
  assign _get_a_mask_acc_T_13=get_a_mask_size_2&get_a_mask_eq_13; 
  assign get_a_mask_hi_hi_hi=get_a_mask_acc_5|_get_a_mask_acc_T_13; 
  assign get_mask={get_a_mask_hi_hi_hi,get_a_mask_hi_hi_lo,get_a_mask_hi_lo_hi,get_a_mask_hi_lo_lo,get_a_mask_lo_hi_hi,get_a_mask_lo_hi_lo,get_a_mask_lo_lo_hi,get_a_mask_lo_lo_lo}; 
  assign _atomics_T=5'h4==s2_req_cmd; 
  assign _atomics_T_1_opcode=_atomics_T ? 3'h3:3'h0; 
  assign atomics_a_size={2'b0,s2_req_size}; 
  assign _atomics_T_1_size=_atomics_T ? atomics_a_size:4'h0; 
  assign _atomics_T_1_source=_atomics_T&a_source; 
  assign atomics_a_address=s2_req_addr[31:0]; 
  assign _atomics_T_1_address=_atomics_T ? atomics_a_address:32'h0; 
  assign _atomics_T_1_mask=_atomics_T ? get_mask:8'h0; 
  assign _atomics_T_1_data=_atomics_T ? pstore1_data:64'h0; 
  assign _atomics_T_2=5'h9==s2_req_cmd; 
  assign _atomics_T_3_opcode=_atomics_T_2 ? 3'h3:_atomics_T_1_opcode; 
  assign _atomics_T_3_param=_atomics_T_2 ? 3'h0:_atomics_T_1_opcode; 
  assign _atomics_T_3_size=_atomics_T_2 ? atomics_a_size:_atomics_T_1_size; 
  assign _atomics_T_3_source=_atomics_T_2 ? a_source:_atomics_T_1_source; 
  assign _atomics_T_3_address=_atomics_T_2 ? atomics_a_address:_atomics_T_1_address; 
  assign _atomics_T_3_mask=_atomics_T_2 ? get_mask:_atomics_T_1_mask; 
  assign _atomics_T_3_data=_atomics_T_2 ? pstore1_data:_atomics_T_1_data; 
  assign _atomics_T_4=5'ha==s2_req_cmd; 
  assign _atomics_T_5_opcode=_atomics_T_4 ? 3'h3:_atomics_T_3_opcode; 
  assign _atomics_T_5_param=_atomics_T_4 ? 3'h1:_atomics_T_3_param; 
  assign _atomics_T_5_size=_atomics_T_4 ? atomics_a_size:_atomics_T_3_size; 
  assign _atomics_T_5_source=_atomics_T_4 ? a_source:_atomics_T_3_source; 
  assign _atomics_T_5_address=_atomics_T_4 ? atomics_a_address:_atomics_T_3_address; 
  assign _atomics_T_5_mask=_atomics_T_4 ? get_mask:_atomics_T_3_mask; 
  assign _atomics_T_5_data=_atomics_T_4 ? pstore1_data:_atomics_T_3_data; 
  assign _atomics_T_6=5'hb==s2_req_cmd; 
  assign _atomics_T_7_opcode=_atomics_T_6 ? 3'h3:_atomics_T_5_opcode; 
  assign _atomics_T_7_param=_atomics_T_6 ? 3'h2:_atomics_T_5_param; 
  assign _atomics_T_7_size=_atomics_T_6 ? atomics_a_size:_atomics_T_5_size; 
  assign _atomics_T_7_source=_atomics_T_6 ? a_source:_atomics_T_5_source; 
  assign _atomics_T_7_address=_atomics_T_6 ? atomics_a_address:_atomics_T_5_address; 
  assign _atomics_T_7_mask=_atomics_T_6 ? get_mask:_atomics_T_5_mask; 
  assign _atomics_T_7_data=_atomics_T_6 ? pstore1_data:_atomics_T_5_data; 
  assign _atomics_T_8=5'h8==s2_req_cmd; 
  assign _atomics_T_9_opcode=_atomics_T_8 ? 3'h2:_atomics_T_7_opcode; 
  assign _atomics_T_9_param=_atomics_T_8 ? 3'h4:_atomics_T_7_param; 
  assign _atomics_T_9_size=_atomics_T_8 ? atomics_a_size:_atomics_T_7_size; 
  assign _atomics_T_9_source=_atomics_T_8 ? a_source:_atomics_T_7_source; 
  assign _atomics_T_9_address=_atomics_T_8 ? atomics_a_address:_atomics_T_7_address; 
  assign _atomics_T_9_mask=_atomics_T_8 ? get_mask:_atomics_T_7_mask; 
  assign _atomics_T_9_data=_atomics_T_8 ? pstore1_data:_atomics_T_7_data; 
  assign _atomics_T_10=5'hc==s2_req_cmd; 
  assign _atomics_T_11_opcode=_atomics_T_10 ? 3'h2:_atomics_T_9_opcode; 
  assign _atomics_T_11_param=_atomics_T_10 ? 3'h0:_atomics_T_9_param; 
  assign _atomics_T_11_size=_atomics_T_10 ? atomics_a_size:_atomics_T_9_size; 
  assign _atomics_T_11_source=_atomics_T_10 ? a_source:_atomics_T_9_source; 
  assign _atomics_T_11_address=_atomics_T_10 ? atomics_a_address:_atomics_T_9_address; 
  assign _atomics_T_11_mask=_atomics_T_10 ? get_mask:_atomics_T_9_mask; 
  assign _atomics_T_11_data=_atomics_T_10 ? pstore1_data:_atomics_T_9_data; 
  assign _atomics_T_12=5'hd==s2_req_cmd; 
  assign _atomics_T_13_opcode=_atomics_T_12 ? 3'h2:_atomics_T_11_opcode; 
  assign _atomics_T_13_param=_atomics_T_12 ? 3'h1:_atomics_T_11_param; 
  assign _atomics_T_13_size=_atomics_T_12 ? atomics_a_size:_atomics_T_11_size; 
  assign _atomics_T_13_source=_atomics_T_12 ? a_source:_atomics_T_11_source; 
  assign _atomics_T_13_address=_atomics_T_12 ? atomics_a_address:_atomics_T_11_address; 
  assign _atomics_T_13_mask=_atomics_T_12 ? get_mask:_atomics_T_11_mask; 
  assign _atomics_T_13_data=_atomics_T_12 ? pstore1_data:_atomics_T_11_data; 
  assign _atomics_T_14=5'he==s2_req_cmd; 
  assign _atomics_T_15_opcode=_atomics_T_14 ? 3'h2:_atomics_T_13_opcode; 
  assign _atomics_T_15_param=_atomics_T_14 ? 3'h2:_atomics_T_13_param; 
  assign _atomics_T_15_size=_atomics_T_14 ? atomics_a_size:_atomics_T_13_size; 
  assign _atomics_T_15_source=_atomics_T_14 ? a_source:_atomics_T_13_source; 
  assign _atomics_T_15_address=_atomics_T_14 ? atomics_a_address:_atomics_T_13_address; 
  assign _atomics_T_15_mask=_atomics_T_14 ? get_mask:_atomics_T_13_mask; 
  assign _atomics_T_15_data=_atomics_T_14 ? pstore1_data:_atomics_T_13_data; 
  assign _atomics_T_16=5'hf==s2_req_cmd; 
  assign atomics_opcode=_atomics_T_16 ? 3'h2:_atomics_T_15_opcode; 
  assign atomics_param=_atomics_T_16 ? 3'h3:_atomics_T_15_param; 
  assign atomics_size=_atomics_T_16 ? atomics_a_size:_atomics_T_15_size; 
  assign atomics_source=_atomics_T_16 ? a_source:_atomics_T_15_source; 
  assign atomics_address=_atomics_T_16 ? atomics_a_address:_atomics_T_15_address; 
  assign atomics_mask=_atomics_T_16 ? get_mask:_atomics_T_15_mask; 
  assign atomics_data=_atomics_T_16 ? pstore1_data:_atomics_T_15_data; 
  assign _GEN_356={8'b0,release_ack_addr}; 
  assign _tl_out_a_valid_T_1=s2_req_addr^_GEN_356; 
  assign _tl_out_a_valid_T_3=_tl_out_a_valid_T_1[20:6]==15'h0; 
  assign _tl_out_a_valid_T_4=release_ack_wait&_tl_out_a_valid_T_3; 
  assign _tl_out_a_valid_T_6=s2_valid_cached_miss&~_tl_out_a_valid_T_4; 
  assign _tl_out_a_valid_T_12=_tl_out_a_valid_T_6&~s2_victim_dirty; 
  assign tl_out_a_valid=s2_valid_uncached_pending|_tl_out_a_valid_T_12; 
  assign _tl_out_a_bits_T_6_opcode=s2_read ? atomics_opcode:3'h0; 
  assign _tl_out_a_bits_T_6_param=s2_read ? atomics_param:3'h0; 
  assign _tl_out_a_bits_T_6_size=s2_read ? atomics_size:atomics_a_size; 
  assign _tl_out_a_bits_T_6_source=s2_read ? atomics_source:a_source; 
  assign _tl_out_a_bits_T_6_address=s2_read ? atomics_address:atomics_a_address; 
  assign _tl_out_a_bits_T_6_mask=s2_read ? atomics_mask:get_mask; 
  assign _tl_out_a_bits_T_6_data=s2_read ? atomics_data:pstore1_data; 
  assign _tl_out_a_bits_T_7_opcode=_s2_write_T_1 ? 3'h1:_tl_out_a_bits_T_6_opcode; 
  assign _tl_out_a_bits_T_7_param=_s2_write_T_1 ? 3'h0:_tl_out_a_bits_T_6_param; 
  assign _tl_out_a_bits_T_7_size=_s2_write_T_1 ? atomics_a_size:_tl_out_a_bits_T_6_size; 
  assign _tl_out_a_bits_T_7_source=_s2_write_T_1 ? a_source:_tl_out_a_bits_T_6_source; 
  assign _tl_out_a_bits_T_7_address=_s2_write_T_1 ? atomics_a_address:_tl_out_a_bits_T_6_address; 
  assign putpartial_mask=a_mask[7:0]; 
  assign _tl_out_a_bits_T_7_mask=_s2_write_T_1 ? putpartial_mask:_tl_out_a_bits_T_6_mask; 
  assign _tl_out_a_bits_T_7_data=_s2_write_T_1 ? pstore1_data:_tl_out_a_bits_T_6_data; 
  assign _tl_out_a_bits_T_8_opcode=s2_write ? _tl_out_a_bits_T_7_opcode:3'h4; 
  assign _tl_out_a_bits_T_8_param=s2_write ? _tl_out_a_bits_T_7_param:3'h0; 
  assign _tl_out_a_bits_T_8_size=s2_write ? _tl_out_a_bits_T_7_size:atomics_a_size; 
  assign _tl_out_a_bits_T_8_source=s2_write ? _tl_out_a_bits_T_7_source:a_source; 
  assign _tl_out_a_bits_T_8_address=s2_write ? _tl_out_a_bits_T_7_address:atomics_a_address; 
  assign _tl_out_a_bits_T_8_mask=s2_write ? _tl_out_a_bits_T_7_mask:get_mask; 
  assign _tl_out_a_bits_T_8_data=s2_write ? _tl_out_a_bits_T_7_data:64'h0; 
  assign tl_out_a_bits_a_param={1'b0,s2_grow_param}; 
  assign tl_out_a_bits_a_address=acquire_address[31:0]; 
  assign _a_sel_T=2'h1<<a_source; 
  assign a_sel=_a_sel_T[1]; 
  assign _T_263=auto_out_a_ready&tl_out_a_valid; 
  assign _GEN_142=a_sel|uncachedInFlight_0; 
  assign _beats1_decode_T_1=27'hfff<<auto_out_d_bits_size; 
  assign beats1_decode=~_beats1_decode_T_1[11:3]; 
  assign beats1_opdata=auto_out_d_bits_opcode[0]; 
  assign beats1=beats1_opdata ? beats1_decode:9'h0; 
  assign counter1=counter-9'h1; 
  assign _last_T=counter==9'h1; 
  assign _last_T_1=beats1==9'h0; 
  assign d_last=_last_T|_last_T_1; 
  assign d_done=d_last&_T_271; 
  assign count=beats1&~counter1; 
  assign d_address_inc={count,3'h0}; 
  assign grantIsVoluntary=auto_out_d_bits_opcode==3'h6; 
  assign _blockProbeAfterGrantCount_T_1=blockProbeAfterGrantCount-3'h1; 
  assign _uncachedRespIdxOH_T=2'h1<<auto_out_d_bits_source; 
  assign uncachedRespIdxOH=_uncachedRespIdxOH_T[1]; 
  assign _T_273=cached_grant_wait|reset; 
  assign _T_276=uncachedRespIdxOH&d_last; 
  assign _T_278=uncachedInFlight_0|reset; 
  assign dontCareBits={s1_paddr[31:3],3'h0}; 
  assign _GEN_357={29'b0,uncachedReqs_0_addr[2:0]}; 
  assign _s2_req_addr_T_1=dontCareBits|_GEN_357; 
  assign _T_281=release_ack_wait|reset; 
  assign _GEN_196=grantIsVoluntary ? 1'h0:release_ack_wait; 
  assign _GEN_205=grantIsUncached ? release_ack_wait:_GEN_196; 
  assign _GEN_209=grantIsCached&d_last; 
  assign _GEN_218=grantIsCached ? release_ack_wait:_GEN_205; 
  assign _GEN_231=_T_271 ? _GEN_218:release_ack_wait; 
  assign _bundleOut_0_e_valid_T=auto_out_d_valid&d_first; 
  assign _bundleOut_0_e_valid_T_1=_bundleOut_0_e_valid_T&grantIsCached; 
  assign _bundleOut_0_e_valid_T_2=_bundleOut_0_e_valid_T_1&canAcceptCachedGrant; 
  assign tl_out__e_valid=_T_292 ? 1'h0:_bundleOut_0_e_valid_T_2; 
  assign _T_283=auto_out_e_ready&tl_out__e_valid; 
  assign _T_285=_T_271&d_first; 
  assign _T_286=_T_285&grantIsCached; 
  assign _T_287=_T_283==_T_286; 
  assign _T_289=_T_287|reset; 
  assign _dataArb_io_in_1_valid_T=auto_out_d_valid&grantIsRefill; 
  assign _dataArb_io_in_1_valid_T_1=_dataArb_io_in_1_valid_T&canAcceptCachedGrant; 
  assign _dataArb_io_in_1_bits_addr_T_1={s2_vaddr[39:6],6'h0}; 
  assign _GEN_358={28'b0,d_address_inc}; 
  assign _dataArb_io_in_1_bits_addr_T_2=_dataArb_io_in_1_bits_addr_T_1|_GEN_358; 
  assign _metaArb_io_in_3_valid_T=grantIsCached&d_done; 
  assign _metaArb_io_in_3_bits_data_T_1={s2_write,c_cat_lo,auto_out_d_bits_param}; 
  assign _metaArb_io_in_3_bits_data_T_6=4'h1==_metaArb_io_in_3_bits_data_T_1; 
  assign _metaArb_io_in_3_bits_data_T_7=_metaArb_io_in_3_bits_data_T_6 ? 2'h1:2'h0; 
  assign _metaArb_io_in_3_bits_data_T_8=4'h0==_metaArb_io_in_3_bits_data_T_1; 
  assign _metaArb_io_in_3_bits_data_T_9=_metaArb_io_in_3_bits_data_T_8 ? 2'h2:_metaArb_io_in_3_bits_data_T_7; 
  assign _metaArb_io_in_3_bits_data_T_10=4'h4==_metaArb_io_in_3_bits_data_T_1; 
  assign _metaArb_io_in_3_bits_data_T_11=_metaArb_io_in_3_bits_data_T_10 ? 2'h2:_metaArb_io_in_3_bits_data_T_9; 
  assign _metaArb_io_in_3_bits_data_T_12=4'hc==_metaArb_io_in_3_bits_data_T_1; 
  assign metaArb_io_in_3_bits_data_meta_state=_metaArb_io_in_3_bits_data_T_12 ? 2'h3:_metaArb_io_in_3_bits_data_T_11; 
  assign _GEN_234=auto_out_d_valid ? 1'h0:_GEN_32; 
  assign _GEN_235=auto_out_d_valid|_dataArb_io_in_1_valid_T_1; 
  assign _GEN_236=auto_out_d_valid ? 1'h0:1'h1; 
  assign _metaArb_io_in_6_valid_T_1=~block_probe_for_core_progress|lrscBackingOff; 
  assign _metaArb_io_in_6_valid_T_2=auto_out_b_valid&_metaArb_io_in_6_valid_T_1; 
  assign metaArb_io_in_6_bits_addr_hi=io_cpu_req_bits_addr[39:32]; 
  assign _metaArb_io_in_6_bits_addr_T={metaArb_io_in_6_bits_addr_hi,auto_out_b_bits_address}; 
  assign counter1_1=counter_1-9'h1; 
  assign c_count=beats1_1&~counter1_1; 
  assign releaseRejected=s2_release_data_valid&~_T_297; 
  assign _releaseDataBeat_T={1'h0,c_count}; 
  assign _releaseDataBeat_T_1={1'h0,s2_release_data_valid}; 
  assign _GEN_359={1'b0,s1_release_data_valid}; 
  assign _releaseDataBeat_T_3=_GEN_359+_releaseDataBeat_T_1; 
  assign _releaseDataBeat_T_4=releaseRejected ? 2'h0:_releaseDataBeat_T_3; 
  assign _GEN_360={8'b0,_releaseDataBeat_T_4}; 
  assign releaseDataBeat=_releaseDataBeat_T+_GEN_360; 
  assign _T_298=s2_valid_flush_line|s2_flush_valid; 
  assign _T_299=_T_298|io_cpu_s2_nack; 
  assign _T_301=_T_299|reset; 
  assign discard_line=s2_valid_flush_line&s2_req_size[1]; 
  assign _release_state_T_1=s2_victim_dirty&~discard_line; 
  assign _release_state_T_13=_release_state_T_1 ? 4'h1:4'h6; 
  assign probe_bits_lo=s2_req_addr[11:6]; 
  assign _probe_bits_T_1={s2_victim_tag,probe_bits_lo}; 
  assign res_2_address={_probe_bits_T_1,6'h0}; 
  assign _GEN_244=s2_want_victimize ? _release_state_T_13:release_state; 
  assign _release_state_T_14=releaseDone ? 4'h7:4'h3; 
  assign _release_state_T_15=releaseDone ? 4'h0:4'h5; 
  assign _GEN_255=_T_303 ? s2_report_param:3'h5; 
  assign _GEN_261=_T_303 ? _release_state_T_14:_release_state_T_15; 
  assign _GEN_263=s2_prb_ack_data ? 4'h2:_GEN_261; 
  assign _GEN_266=s2_prb_ack_data ? 3'h5:_GEN_255; 
  assign _GEN_273=s2_meta_error ? 4'h4:_GEN_263; 
  assign _GEN_276=s2_meta_error ? 3'h5:_GEN_266; 
  assign _GEN_284=s2_probe ? _GEN_273:_GEN_244; 
  assign _GEN_287=s2_probe ? _GEN_276:3'h5; 
  assign _T_304=release_state==4'h4; 
  assign _metaArb_io_in_6_bits_addr_T_1={metaArb_io_in_6_bits_addr_hi,probe_bits_address}; 
  assign _GEN_294=metaArb_io_in_6_ready ? 4'h0:_GEN_284; 
  assign _GEN_295=metaArb_io_in_6_ready|s1_probe_x12; 
  assign _GEN_299=_T_304 ? _GEN_294:_GEN_284; 
  assign _GEN_301=releaseDone ? 4'h0:_GEN_299; 
  assign _GEN_303=_T_305 ? _GEN_301:_GEN_299; 
  assign _GEN_307=_T_306 ? s2_report_param:_GEN_287; 
  assign _GEN_316=_T_307 ? s2_report_param:_GEN_307; 
  assign _T_315=_T_297&c_first; 
  assign _GEN_331=_T_315|_GEN_231; 
  assign newCoh_state=_T_312 ? voluntaryNewCoh_state:probeNewCoh_state; 
  assign _dataArb_io_in_2_valid_T=releaseDataBeat<10'h8; 
  assign _dataArb_io_in_2_bits_addr_T_1={probe_bits_address[11:6],6'h0}; 
  assign _dataArb_io_in_2_bits_addr_T_3={releaseDataBeat[2:0],3'h0}; 
  assign _GEN_363={6'b0,_dataArb_io_in_2_bits_addr_T_3}; 
  assign _metaArb_io_in_4_valid_T_1=release_state==4'h7; 
  assign metaArb_io_in_4_bits_addr_lo=probe_bits_address[11:0]; 
  assign metaArb_io_in_4_bits_data_meta_tag=probe_bits_address[31:12]; 
  assign _T_316=metaArb_io_in_4_ready&metaArb_io_in_4_valid; 
  assign _io_cpu_ordered_T_4=s1_valid|s2_valid; 
  assign _io_cpu_ordered_T_5=_io_cpu_ordered_T_4|cached_grant_wait; 
  assign _io_cpu_ordered_T_7=_io_cpu_ordered_T_5|_s2_valid_cached_miss_T_2; 
  assign _s1_xcpt_valid_T_1=tlb_io_req_valid; 
  assign _T_321=~s2_valid_hit_pre_data_ecc_and_waw|reset; 
  assign io_cpu_resp_bits_data_shifted=get_a_mask_bit ? s2_data_corrected[63:32]:s2_data_corrected[31:0]; 
  assign _io_cpu_resp_bits_data_T=s2_req_size==2'h2; 
  assign _io_cpu_resp_bits_data_T_3=s2_req_signed&io_cpu_resp_bits_data_shifted[31]; 
  assign _io_cpu_resp_bits_data_T_5=_io_cpu_resp_bits_data_T_3 ? 32'hffffffff:32'h0; 
  assign io_cpu_resp_bits_data_hi=_io_cpu_resp_bits_data_T ? _io_cpu_resp_bits_data_T_5:s2_data_corrected[63:32]; 
  assign _io_cpu_resp_bits_data_T_7={io_cpu_resp_bits_data_hi,io_cpu_resp_bits_data_shifted}; 
  assign io_cpu_resp_bits_data_shifted_1=get_a_mask_bit_1 ? _io_cpu_resp_bits_data_T_7[31:16]:_io_cpu_resp_bits_data_T_7[15:0]; 
  assign _io_cpu_resp_bits_data_T_8=s2_req_size==2'h1; 
  assign _io_cpu_resp_bits_data_T_11=s2_req_signed&io_cpu_resp_bits_data_shifted_1[15]; 
  assign _io_cpu_resp_bits_data_T_13=_io_cpu_resp_bits_data_T_11 ? 48'hffffffffffff:48'h0; 
  assign io_cpu_resp_bits_data_hi_1=_io_cpu_resp_bits_data_T_8 ? _io_cpu_resp_bits_data_T_13:_io_cpu_resp_bits_data_T_7[63:16]; 
  assign _io_cpu_resp_bits_data_T_15={io_cpu_resp_bits_data_hi_1,io_cpu_resp_bits_data_shifted_1}; 
  assign io_cpu_resp_bits_data_shifted_2=get_a_mask_bit_2 ? _io_cpu_resp_bits_data_T_15[15:8]:_io_cpu_resp_bits_data_T_15[7:0]; 
  assign io_cpu_resp_bits_data_lo_2=_s2_write_T_3 ? 8'h0:io_cpu_resp_bits_data_shifted_2; 
  assign _io_cpu_resp_bits_data_T_16=s2_req_size==2'h0; 
  assign _io_cpu_resp_bits_data_T_17=_io_cpu_resp_bits_data_T_16|_s2_write_T_3; 
  assign _io_cpu_resp_bits_data_T_19=s2_req_signed&io_cpu_resp_bits_data_lo_2[7]; 
  assign _io_cpu_resp_bits_data_T_21=_io_cpu_resp_bits_data_T_19 ? 56'hffffffffffffff:56'h0; 
  assign io_cpu_resp_bits_data_hi_2=_io_cpu_resp_bits_data_T_17 ? _io_cpu_resp_bits_data_T_21:_io_cpu_resp_bits_data_T_15[63:8]; 
  assign _io_cpu_resp_bits_data_T_23={io_cpu_resp_bits_data_hi_2,io_cpu_resp_bits_data_lo_2}; 
  assign _GEN_364={63'b0,s2_sc_fail}; 
  assign _GEN_349=REG|resetting; 
  assign flushCounterNext=flushCounter+8'h1; 
  assign flushDone=flushCounterNext[8:6]==3'h4; 
  assign _s1_flush_valid_T=metaArb_io_in_5_ready&metaArb_io_in_5_valid; 
  assign _s1_flush_valid_T_2=_s1_flush_valid_T&~s1_flush_valid; 
  assign _s1_flush_valid_T_4=_s1_flush_valid_T_2&~s2_flush_valid_pre_tag_ecc; 
  assign _s1_flush_valid_T_6=_s1_flush_valid_T_4&_io_cpu_req_ready_T; 
  assign metaArb_io_in_5_bits_addr_lo={metaArb_io_in_5_bits_idx,6'h0}; 
  assign _GEN_351=resetting ? flushCounterNext:{1'b0,flushCounter}; 
  assign io_cpu_perf_release_counter1=io_cpu_perf_release_counter-9'h1; 
  assign io_cpu_perf_release_first=io_cpu_perf_release_counter==9'h0; 
  assign _io_cpu_perf_release_last_T=io_cpu_perf_release_counter==9'h1; 
  assign io_cpu_perf_release_last=_io_cpu_perf_release_last_T|_last_T_3; 
  assign auto_out_a_valid=s2_valid_uncached_pending|_tl_out_a_valid_T_12; 
  assign auto_out_a_bits_opcode=s2_uncached ? _tl_out_a_bits_T_8_opcode:3'h6; 
  assign auto_out_a_bits_param=s2_uncached ? _tl_out_a_bits_T_8_param:tl_out_a_bits_a_param; 
  assign auto_out_a_bits_size=s2_uncached ? _tl_out_a_bits_T_8_size:4'h6; 
  assign auto_out_a_bits_source=s2_uncached ? _tl_out_a_bits_T_8_source:1'h0; 
  assign auto_out_a_bits_address=s2_uncached ? _tl_out_a_bits_T_8_address:tl_out_a_bits_a_address; 
  assign auto_out_a_bits_mask=s2_uncached ? _tl_out_a_bits_T_8_mask:8'hff; 
  assign auto_out_a_bits_data=s2_uncached ? _tl_out_a_bits_T_8_data:64'h0; 
  assign auto_out_b_ready=metaArb_io_in_6_ready&~_bundleOut_0_b_ready_T_2; 
  assign auto_out_c_valid=_T_306|_GEN_302; 
  assign auto_out_c_bits_opcode=_T_312 ? _GEN_323:_GEN_315; 
  assign auto_out_c_bits_param=_T_312 ? s2_shrink_param:_GEN_316; 
  assign auto_out_c_bits_size=_T_312 ? 4'h6:probe_bits_size; 
  assign auto_out_c_bits_source=probe_bits_source; 
  assign auto_out_c_bits_address=probe_bits_address; 
  assign auto_out_c_bits_data={s2_data_corrected_hi,s2_data_corrected_lo}; 
  assign auto_out_d_ready=_T_294 ? 1'h0:_GEN_233; 
  assign auto_out_e_valid=_T_292 ? 1'h0:_bundleOut_0_e_valid_T_2; 
  assign auto_out_e_bits_sink=auto_out_d_bits_sink; 
  assign io_cpu_req_ready=_T_294 ? _GEN_234:_GEN_32; 
  assign io_cpu_s2_nack=_io_cpu_s2_nack_T_3&~s2_valid_hit_pre_data_ecc_and_waw; 
  assign io_cpu_resp_valid=s2_valid_hit_pre_data_ecc_and_waw|doUncachedResp; 
  assign io_cpu_resp_bits_tag=s2_req_tag; 
  assign io_cpu_resp_bits_size=s2_req_size; 
  assign io_cpu_resp_bits_data=_io_cpu_resp_bits_data_T_23|_GEN_364; 
  assign io_cpu_resp_bits_replay=doUncachedResp; 
  assign io_cpu_resp_bits_has_data=_s2_read_T_4|_s2_write_T_21; 
  assign io_cpu_resp_bits_data_word_bypass={io_cpu_resp_bits_data_hi,io_cpu_resp_bits_data_shifted}; 
  assign io_cpu_replay_next=_T_271&grantIsUncachedData; 
  assign io_cpu_s2_xcpt_ma_ld=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ma_ld; 
  assign io_cpu_s2_xcpt_ma_st=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ma_st; 
  assign io_cpu_s2_xcpt_pf_ld=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_pf_ld; 
  assign io_cpu_s2_xcpt_pf_st=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_pf_st; 
  assign io_cpu_s2_xcpt_ae_ld=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ae_ld; 
  assign io_cpu_s2_xcpt_ae_st=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ae_st; 
  assign io_cpu_ordered=~_io_cpu_ordered_T_7; 
  assign io_cpu_perf_release=io_cpu_perf_release_last&_T_297; 
  assign io_cpu_perf_grant=auto_out_d_valid&d_last; 
  assign io_ptw_req_valid=tlb_io_ptw_req_valid; 
  assign io_ptw_req_bits_bits_addr=tlb_io_ptw_req_bits_bits_addr; 
  assign tlb_clock=gated_clock; 
  assign tlb_reset=reset; 
  assign tlb_io_req_valid=s1_valid_masked&s1_cmd_uses_tlb; 
  assign tlb_io_req_bits_vaddr=s1_tlb_req_vaddr; 
  assign tlb_io_req_bits_passthrough=s1_tlb_req_passthrough; 
  assign tlb_io_req_bits_size=s1_tlb_req_size; 
  assign tlb_io_req_bits_cmd=s1_tlb_req_cmd; 
  assign tlb_io_sfence_valid=s1_valid_masked&s1_sfence; 
  assign tlb_io_sfence_bits_rs1=s1_req_size[0]; 
  assign tlb_io_sfence_bits_rs2=s1_req_size[1]; 
  assign tlb_io_sfence_bits_addr=s1_req_addr[38:0]; 
  assign tlb_io_ptw_req_ready=io_ptw_req_ready; 
  assign tlb_io_ptw_resp_valid=io_ptw_resp_valid; 
  assign tlb_io_ptw_resp_bits_ae=io_ptw_resp_bits_ae; 
  assign tlb_io_ptw_resp_bits_pte_ppn=io_ptw_resp_bits_pte_ppn; 
  assign tlb_io_ptw_resp_bits_pte_d=io_ptw_resp_bits_pte_d; 
  assign tlb_io_ptw_resp_bits_pte_a=io_ptw_resp_bits_pte_a; 
  assign tlb_io_ptw_resp_bits_pte_g=io_ptw_resp_bits_pte_g; 
  assign tlb_io_ptw_resp_bits_pte_u=io_ptw_resp_bits_pte_u; 
  assign tlb_io_ptw_resp_bits_pte_x=io_ptw_resp_bits_pte_x; 
  assign tlb_io_ptw_resp_bits_pte_w=io_ptw_resp_bits_pte_w; 
  assign tlb_io_ptw_resp_bits_pte_r=io_ptw_resp_bits_pte_r; 
  assign tlb_io_ptw_resp_bits_pte_v=io_ptw_resp_bits_pte_v; 
  assign tlb_io_ptw_resp_bits_level=io_ptw_resp_bits_level; 
  assign tlb_io_ptw_resp_bits_homogeneous=io_ptw_resp_bits_homogeneous; 
  assign tlb_io_ptw_ptbr_mode=io_ptw_ptbr_mode; 
  assign tlb_io_ptw_status_debug=io_ptw_status_debug; 
  assign tlb_io_ptw_status_dprv=io_ptw_status_dprv; 
  assign tlb_io_ptw_status_mxr=io_ptw_status_mxr; 
  assign tlb_io_ptw_status_sum=io_ptw_status_sum; 
  assign tlb_io_ptw_pmp_0_cfg_l=io_ptw_pmp_0_cfg_l; 
  assign tlb_io_ptw_pmp_0_cfg_a=io_ptw_pmp_0_cfg_a; 
  assign tlb_io_ptw_pmp_0_cfg_x=io_ptw_pmp_0_cfg_x; 
  assign tlb_io_ptw_pmp_0_cfg_w=io_ptw_pmp_0_cfg_w; 
  assign tlb_io_ptw_pmp_0_cfg_r=io_ptw_pmp_0_cfg_r; 
  assign tlb_io_ptw_pmp_0_addr=io_ptw_pmp_0_addr; 
  assign tlb_io_ptw_pmp_0_mask=io_ptw_pmp_0_mask; 
  assign tlb_io_ptw_pmp_1_cfg_l=io_ptw_pmp_1_cfg_l; 
  assign tlb_io_ptw_pmp_1_cfg_a=io_ptw_pmp_1_cfg_a; 
  assign tlb_io_ptw_pmp_1_cfg_x=io_ptw_pmp_1_cfg_x; 
  assign tlb_io_ptw_pmp_1_cfg_w=io_ptw_pmp_1_cfg_w; 
  assign tlb_io_ptw_pmp_1_cfg_r=io_ptw_pmp_1_cfg_r; 
  assign tlb_io_ptw_pmp_1_addr=io_ptw_pmp_1_addr; 
  assign tlb_io_ptw_pmp_1_mask=io_ptw_pmp_1_mask; 
  assign tlb_io_ptw_pmp_2_cfg_l=io_ptw_pmp_2_cfg_l; 
  assign tlb_io_ptw_pmp_2_cfg_a=io_ptw_pmp_2_cfg_a; 
  assign tlb_io_ptw_pmp_2_cfg_x=io_ptw_pmp_2_cfg_x; 
  assign tlb_io_ptw_pmp_2_cfg_w=io_ptw_pmp_2_cfg_w; 
  assign tlb_io_ptw_pmp_2_cfg_r=io_ptw_pmp_2_cfg_r; 
  assign tlb_io_ptw_pmp_2_addr=io_ptw_pmp_2_addr; 
  assign tlb_io_ptw_pmp_2_mask=io_ptw_pmp_2_mask; 
  assign tlb_io_ptw_pmp_3_cfg_l=io_ptw_pmp_3_cfg_l; 
  assign tlb_io_ptw_pmp_3_cfg_a=io_ptw_pmp_3_cfg_a; 
  assign tlb_io_ptw_pmp_3_cfg_x=io_ptw_pmp_3_cfg_x; 
  assign tlb_io_ptw_pmp_3_cfg_w=io_ptw_pmp_3_cfg_w; 
  assign tlb_io_ptw_pmp_3_cfg_r=io_ptw_pmp_3_cfg_r; 
  assign tlb_io_ptw_pmp_3_addr=io_ptw_pmp_3_addr; 
  assign tlb_io_ptw_pmp_3_mask=io_ptw_pmp_3_mask; 
  assign tlb_io_ptw_pmp_4_cfg_l=io_ptw_pmp_4_cfg_l; 
  assign tlb_io_ptw_pmp_4_cfg_a=io_ptw_pmp_4_cfg_a; 
  assign tlb_io_ptw_pmp_4_cfg_x=io_ptw_pmp_4_cfg_x; 
  assign tlb_io_ptw_pmp_4_cfg_w=io_ptw_pmp_4_cfg_w; 
  assign tlb_io_ptw_pmp_4_cfg_r=io_ptw_pmp_4_cfg_r; 
  assign tlb_io_ptw_pmp_4_addr=io_ptw_pmp_4_addr; 
  assign tlb_io_ptw_pmp_4_mask=io_ptw_pmp_4_mask; 
  assign tlb_io_ptw_pmp_5_cfg_l=io_ptw_pmp_5_cfg_l; 
  assign tlb_io_ptw_pmp_5_cfg_a=io_ptw_pmp_5_cfg_a; 
  assign tlb_io_ptw_pmp_5_cfg_x=io_ptw_pmp_5_cfg_x; 
  assign tlb_io_ptw_pmp_5_cfg_w=io_ptw_pmp_5_cfg_w; 
  assign tlb_io_ptw_pmp_5_cfg_r=io_ptw_pmp_5_cfg_r; 
  assign tlb_io_ptw_pmp_5_addr=io_ptw_pmp_5_addr; 
  assign tlb_io_ptw_pmp_5_mask=io_ptw_pmp_5_mask; 
  assign tlb_io_ptw_pmp_6_cfg_l=io_ptw_pmp_6_cfg_l; 
  assign tlb_io_ptw_pmp_6_cfg_a=io_ptw_pmp_6_cfg_a; 
  assign tlb_io_ptw_pmp_6_cfg_x=io_ptw_pmp_6_cfg_x; 
  assign tlb_io_ptw_pmp_6_cfg_w=io_ptw_pmp_6_cfg_w; 
  assign tlb_io_ptw_pmp_6_cfg_r=io_ptw_pmp_6_cfg_r; 
  assign tlb_io_ptw_pmp_6_addr=io_ptw_pmp_6_addr; 
  assign tlb_io_ptw_pmp_6_mask=io_ptw_pmp_6_mask; 
  assign tlb_io_ptw_pmp_7_cfg_l=io_ptw_pmp_7_cfg_l; 
  assign tlb_io_ptw_pmp_7_cfg_a=io_ptw_pmp_7_cfg_a; 
  assign tlb_io_ptw_pmp_7_cfg_x=io_ptw_pmp_7_cfg_x; 
  assign tlb_io_ptw_pmp_7_cfg_w=io_ptw_pmp_7_cfg_w; 
  assign tlb_io_ptw_pmp_7_cfg_r=io_ptw_pmp_7_cfg_r; 
  assign tlb_io_ptw_pmp_7_addr=io_ptw_pmp_7_addr; 
  assign tlb_io_ptw_pmp_7_mask=io_ptw_pmp_7_mask; 
  assign pma_checker_clock=gated_clock; 
  assign pma_checker_reset=reset; 
  assign pma_checker_io_req_valid=1'h0; 
  assign pma_checker_io_req_bits_vaddr=40'h0; 
  assign pma_checker_io_req_bits_passthrough=1'h1; 
  assign pma_checker_io_req_bits_size=s1_req_size; 
  assign pma_checker_io_req_bits_cmd=s1_req_cmd; 
  assign pma_checker_io_sfence_valid=1'h0; 
  assign pma_checker_io_sfence_bits_rs1=1'h0; 
  assign pma_checker_io_sfence_bits_rs2=1'h0; 
  assign pma_checker_io_sfence_bits_addr=39'h0; 
  assign pma_checker_io_ptw_req_ready=1'h0; 
  assign pma_checker_io_ptw_resp_valid=1'h0; 
  assign pma_checker_io_ptw_resp_bits_ae=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_ppn=54'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_d=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_a=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_g=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_u=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_x=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_w=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_r=1'h0; 
  assign pma_checker_io_ptw_resp_bits_pte_v=1'h0; 
  assign pma_checker_io_ptw_resp_bits_level=2'h0; 
  assign pma_checker_io_ptw_resp_bits_homogeneous=1'h0; 
  assign pma_checker_io_ptw_ptbr_mode=4'h0; 
  assign pma_checker_io_ptw_status_debug=1'h0; 
  assign pma_checker_io_ptw_status_dprv=2'h0; 
  assign pma_checker_io_ptw_status_mxr=1'h0; 
  assign pma_checker_io_ptw_status_sum=1'h0; 
  assign pma_checker_io_ptw_pmp_0_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_0_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_0_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_0_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_0_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_0_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_0_mask=32'h0; 
  assign pma_checker_io_ptw_pmp_1_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_1_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_1_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_1_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_1_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_1_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_1_mask=32'h0; 
  assign pma_checker_io_ptw_pmp_2_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_2_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_2_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_2_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_2_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_2_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_2_mask=32'h0; 
  assign pma_checker_io_ptw_pmp_3_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_3_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_3_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_3_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_3_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_3_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_3_mask=32'h0; 
  assign pma_checker_io_ptw_pmp_4_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_4_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_4_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_4_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_4_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_4_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_4_mask=32'h0; 
  assign pma_checker_io_ptw_pmp_5_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_5_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_5_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_5_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_5_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_5_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_5_mask=32'h0; 
  assign pma_checker_io_ptw_pmp_6_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_6_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_6_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_6_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_6_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_6_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_6_mask=32'h0; 
  assign pma_checker_io_ptw_pmp_7_cfg_l=1'h0; 
  assign pma_checker_io_ptw_pmp_7_cfg_a=2'h0; 
  assign pma_checker_io_ptw_pmp_7_cfg_x=1'h0; 
  assign pma_checker_io_ptw_pmp_7_cfg_w=1'h0; 
  assign pma_checker_io_ptw_pmp_7_cfg_r=1'h0; 
  assign pma_checker_io_ptw_pmp_7_addr=30'h0; 
  assign pma_checker_io_ptw_pmp_7_mask=32'h0; 
  assign lfsr_prng_clock=gated_clock; 
  assign lfsr_prng_reset=reset; 
  assign lfsr_prng_io_increment=_T_271&_GEN_209; 
  assign metaArb_io_in_0_valid=resetting; 
  assign metaArb_io_in_0_bits_addr=metaArb_io_in_5_bits_addr; 
  assign metaArb_io_in_0_bits_idx=metaArb_io_in_5_bits_idx; 
  assign metaArb_io_in_1_valid=s2_meta_error&_metaArb_io_in_1_valid_T_1; 
  assign metaArb_io_in_1_bits_addr={dataArb_io_in_3_bits_addr_hi,metaArb_io_in_1_bits_addr_lo}; 
  assign metaArb_io_in_1_bits_idx=s2_probe ? probe_bits_address[11:6]:s2_vaddr[11:6]; 
  assign metaArb_io_in_1_bits_data={new_meta_coh_state,s2_meta_corrected_3_tag}; 
  assign metaArb_io_in_2_valid=s2_valid_hit_pre_data_ecc_and_waw&s2_update_meta; 
  assign metaArb_io_in_2_bits_addr={dataArb_io_in_3_bits_addr_hi,metaArb_io_in_2_bits_addr_lo}; 
  assign metaArb_io_in_2_bits_idx=s2_vaddr[11:6]; 
  assign metaArb_io_in_2_bits_way_en=s2_hit_valid ? s2_hit_way:s2_victim_way; 
  assign metaArb_io_in_2_bits_data={s2_grow_param,metaArb_io_in_2_bits_data_meta_tag}; 
  assign metaArb_io_in_3_valid=_metaArb_io_in_3_valid_T&~auto_out_d_bits_denied; 
  assign metaArb_io_in_3_bits_addr={dataArb_io_in_3_bits_addr_hi,metaArb_io_in_2_bits_addr_lo}; 
  assign metaArb_io_in_3_bits_idx=s2_vaddr[11:6]; 
  assign metaArb_io_in_3_bits_way_en=refill_way; 
  assign metaArb_io_in_3_bits_data={metaArb_io_in_3_bits_data_meta_state,metaArb_io_in_2_bits_data_meta_tag}; 
  assign metaArb_io_in_4_valid=_T_309|_metaArb_io_in_4_valid_T_1; 
  assign metaArb_io_in_4_bits_addr={dataArb_io_in_3_bits_addr_hi,metaArb_io_in_4_bits_addr_lo}; 
  assign metaArb_io_in_4_bits_idx=probe_bits_address[11:6]; 
  assign metaArb_io_in_4_bits_way_en=_T_312 ? s2_victim_or_hit_way:s2_probe_way; 
  assign metaArb_io_in_4_bits_data={newCoh_state,metaArb_io_in_4_bits_data_meta_tag}; 
  assign metaArb_io_in_5_valid=1'h0; 
  assign metaArb_io_in_5_bits_addr={dataArb_io_in_3_bits_addr_hi,metaArb_io_in_5_bits_addr_lo}; 
  assign metaArb_io_in_5_bits_idx=flushCounter[5:0]; 
  assign metaArb_io_in_6_valid=_T_304|_metaArb_io_in_6_valid_T_2; 
  assign metaArb_io_in_6_bits_addr=_T_304 ? _metaArb_io_in_6_bits_addr_T_1:_metaArb_io_in_6_bits_addr_T; 
  assign metaArb_io_in_6_bits_idx=_T_304 ? probe_bits_address[11:6]:auto_out_b_bits_address[11:6]; 
  assign metaArb_io_in_6_bits_way_en=metaArb_io_in_4_bits_way_en; 
  assign metaArb_io_in_6_bits_data=metaArb_io_in_4_bits_data; 
  assign metaArb_io_in_7_valid=io_cpu_req_valid; 
  assign metaArb_io_in_7_bits_addr=io_cpu_req_bits_addr; 
  assign metaArb_io_in_7_bits_idx=dataArb_io_in_3_bits_addr[11:6]; 
  assign metaArb_io_in_7_bits_way_en=metaArb_io_in_4_bits_way_en; 
  assign metaArb_io_in_7_bits_data=metaArb_io_in_4_bits_data; 
  assign data_clock=gated_clock; 
  assign data_io_req_valid=dataArb_io_out_valid; 
  assign data_io_req_bits_addr=dataArb_io_out_bits_addr; 
  assign data_io_req_bits_write=dataArb_io_out_bits_write; 
  assign data_io_req_bits_wdata=dataArb_io_out_bits_wdata; 
  assign data_io_req_bits_eccMask=dataArb_io_out_bits_eccMask; 
  assign data_io_req_bits_way_en=dataArb_io_out_bits_way_en; 
  assign dataArb_io_in_0_valid=pstore_drain_structural|_pstore_drain_T_10; 
  assign dataArb_io_in_0_bits_addr=_dataArb_io_in_0_bits_addr_T[11:0]; 
  assign dataArb_io_in_0_bits_write=pstore_drain_structural|_pstore_drain_T_10; 
  assign dataArb_io_in_0_bits_wdata={dataArb_io_in_0_bits_wdata_hi,dataArb_io_in_0_bits_wdata_lo}; 
  assign dataArb_io_in_0_bits_eccMask={dataArb_io_in_0_bits_eccMask_hi,dataArb_io_in_0_bits_eccMask_lo}; 
  assign dataArb_io_in_0_bits_way_en=pstore2_valid ? pstore2_way:pstore1_way; 
  assign dataArb_io_in_1_valid=_T_294 ? _GEN_235:_dataArb_io_in_1_valid_T_1; 
  assign dataArb_io_in_1_bits_addr=_dataArb_io_in_1_bits_addr_T_2[11:0]; 
  assign dataArb_io_in_1_bits_write=_T_294 ? _GEN_236:1'h1; 
  assign dataArb_io_in_1_bits_wdata={tl_d_data_encoded_hi,tl_d_data_encoded_lo}; 
  assign dataArb_io_in_1_bits_way_en=refill_way; 
  assign dataArb_io_in_2_valid=inWriteback&_dataArb_io_in_2_valid_T; 
  assign dataArb_io_in_2_bits_addr=_dataArb_io_in_2_bits_addr_T_1|_GEN_363; 
  assign dataArb_io_in_2_bits_wdata=dataArb_io_in_1_bits_wdata; 
  assign dataArb_io_in_3_valid=io_cpu_req_valid&res; 
  assign dataArb_io_in_3_bits_addr=_dataArb_io_in_3_bits_addr_T[11:0]; 
  assign dataArb_io_in_3_bits_wdata=dataArb_io_in_1_bits_wdata; 
  assign dataArb_io_in_3_bits_wordMask=1'h1; 
  assign amoalu_io_mask=pstore1_mask; 
  assign amoalu_io_cmd=pstore1_cmd; 
  assign amoalu_io_lhs={s2_data_corrected_hi,s2_data_corrected_lo}; 
  assign amoalu_io_rhs=pstore1_data; 
  assign _GEN_367=_T_271&grantIsCached; 
  assign _GEN_370=_T_271&~grantIsCached; 
  assign _GEN_371=_GEN_370&grantIsUncached; 
  assign _GEN_372=_GEN_371&_T_276; 
  assign _GEN_380=_GEN_370&~grantIsUncached; 
  assign _GEN_381=_GEN_380&grantIsVoluntary; 
  assign DCache_cov_read_addr=DCache_state; 
  assign DCache_cov_read_data=DCache_cov[DCache_cov_read_addr]; 
  assign DCache_cov_write_data=1'h1; 
  assign DCache_cov_write_addr=DCache_state; 
  assign DCache_cov_write_mask=1'h1; 
  assign DCache_cov_write_en=1'h1; 
  assign mux_cond_0=s1_req_addr[0]; 
  assign mux_cond_1=get_a_mask_bit_2; 
  assign mux_cond_2=s1_req_addr[2]; 
  assign mux_cond_3=get_a_mask_bit; 
  assign mux_cond_4=get_a_mask_bit_1; 
  assign mux_cond_5=s1_req_addr[1]; 
  assign s2_req_size_shl={s2_req_size,3'h0}; 
  assign s2_req_size_pad={15'h0,s2_req_size_shl}; 
  assign pstore1_held_shl={pstore1_held,9'h0}; 
  assign pstore1_held_pad={10'h0,pstore1_held_shl}; 
  assign s2_req_signed_shl={s2_req_signed,5'h0}; 
  assign s2_req_signed_pad={14'h0,s2_req_signed_shl}; 
  assign pstore2_valid_shl={pstore2_valid,10'h0}; 
  assign pstore2_valid_pad={9'h0,pstore2_valid_shl}; 
  assign s1_flush_valid_shl={s1_flush_valid,17'h0}; 
  assign s1_flush_valid_pad={2'h0,s1_flush_valid_shl}; 
  assign uncachedInFlight_0_shl={uncachedInFlight_0,8'h0}; 
  assign uncachedInFlight_0_pad={11'h0,uncachedInFlight_0_shl}; 
  assign blockUncachedGrant_shl={blockUncachedGrant,18'h0}; 
  assign blockUncachedGrant_pad={1'h0,blockUncachedGrant_shl}; 
  assign probe_bits_param_shl={probe_bits_param,12'h0}; 
  assign probe_bits_param_pad={6'h0,probe_bits_param_shl}; 
  assign s2_flush_valid_pre_tag_ecc_shl={s2_flush_valid_pre_tag_ecc,16'h0}; 
  assign s2_flush_valid_pre_tag_ecc_pad={3'h0,s2_flush_valid_pre_tag_ecc_shl}; 
  assign s1_read_mask_shl={s1_read_mask,10'h0}; 
  assign s1_read_mask_pad={9'h0,s1_read_mask_shl}; 
  assign s2_victim_way_r_shl={s2_victim_way_r,12'h0}; 
  assign s2_victim_way_r_pad={6'h0,s2_victim_way_r_shl}; 
  assign s1_probe_shl={s1_probe,13'h0}; 
  assign s1_probe_pad={6'h0,s1_probe_shl}; 
  assign release_ack_wait_shl={release_ack_wait,2'h0}; 
  assign release_ack_wait_pad={17'h0,release_ack_wait_shl}; 
  assign s2_hit_state_state_shl={s2_hit_state_state,11'h0}; 
  assign s2_hit_state_state_pad={7'h0,s2_hit_state_state_shl}; 
  assign cached_grant_wait_shl={cached_grant_wait,15'h0}; 
  assign cached_grant_wait_pad={4'h0,cached_grant_wait_shl}; 
  assign s1_valid_shl={s1_valid,19'h0}; 
  assign s1_valid_pad=s1_valid_shl; 
  assign s2_pma_cacheable_shl={s2_pma_cacheable,18'h0}; 
  assign s2_pma_cacheable_pad={1'h0,s2_pma_cacheable_shl}; 
  assign s1_did_read_shl={s1_did_read,17'h0}; 
  assign s1_did_read_pad={2'h0,s1_did_read_shl}; 
  assign s2_probe_shl={s2_probe,19'h0}; 
  assign s2_probe_pad=s2_probe_shl; 
  assign s2_hit_way_shl={s2_hit_way,3'h0}; 
  assign s2_hit_way_pad={13'h0,s2_hit_way_shl}; 
  assign s2_not_nacked_in_s1_shl={s2_not_nacked_in_s1,9'h0}; 
  assign s2_not_nacked_in_s1_pad={10'h0,s2_not_nacked_in_s1_shl}; 
  assign s2_probe_state_state_shl={s2_probe_state_state,17'h0}; 
  assign s2_probe_state_state_pad={1'h0,s2_probe_state_state_shl}; 
  assign s1_req_size_shl={s1_req_size,3'h0}; 
  assign s1_req_size_pad={15'h0,s1_req_size_shl}; 
  assign pstore1_rmw_r_shl={pstore1_rmw_r,14'h0}; 
  assign pstore1_rmw_r_pad={5'h0,pstore1_rmw_r_shl}; 
  assign s2_release_data_valid_shl={s2_release_data_valid,7'h0}; 
  assign s2_release_data_valid_pad={12'h0,s2_release_data_valid_shl}; 
  assign s2_valid_shl={s2_valid,8'h0}; 
  assign s2_valid_pad={11'h0,s2_valid_shl}; 
  assign pstore_drain_on_miss_REG_shl={pstore_drain_on_miss_REG,19'h0}; 
  assign pstore_drain_on_miss_REG_pad=pstore_drain_on_miss_REG_shl; 
  assign resetting_shl={resetting,15'h0}; 
  assign resetting_pad={4'h0,resetting_shl}; 
  assign grantInProgress_shl={grantInProgress,19'h0}; 
  assign grantInProgress_pad=grantInProgress_shl; 
  assign s2_probe_way_shl={s2_probe_way,9'h0}; 
  assign s2_probe_way_pad={7'h0,s2_probe_way_shl}; 
  assign mux_cond_0_shl={mux_cond_0,11'h0}; 
  assign mux_cond_0_pad={8'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,1'h0}; 
  assign mux_cond_1_pad={18'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl={mux_cond_2,15'h0}; 
  assign mux_cond_2_pad={4'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,6'h0}; 
  assign mux_cond_3_pad={13'h0,mux_cond_3_shl}; 
  assign mux_cond_4_shl={mux_cond_4,7'h0}; 
  assign mux_cond_4_pad={12'h0,mux_cond_4_shl}; 
  assign mux_cond_5_shl={mux_cond_5,7'h0}; 
  assign mux_cond_5_pad={12'h0,mux_cond_5_shl}; 
  assign DCache_xor15=s2_req_size_pad^pstore1_held_pad; 
  assign DCache_xor16=s2_req_signed_pad^pstore2_valid_pad; 
  assign DCache_xor7=DCache_xor15^DCache_xor16; 
  assign DCache_xor17=s1_flush_valid_pad^uncachedInFlight_0_pad; 
  assign DCache_xor38=probe_bits_param_pad^s2_flush_valid_pre_tag_ecc_pad; 
  assign DCache_xor18=blockUncachedGrant_pad^DCache_xor38; 
  assign DCache_xor8=DCache_xor17^DCache_xor18; 
  assign DCache_xor3=DCache_xor7^DCache_xor8; 
  assign DCache_xor19=s1_read_mask_pad^s2_victim_way_r_pad; 
  assign DCache_xor20=s1_probe_pad^release_ack_wait_pad; 
  assign DCache_xor9=DCache_xor19^DCache_xor20; 
  assign DCache_xor21=s2_hit_state_state_pad^cached_grant_wait_pad; 
  assign DCache_xor46=s2_pma_cacheable_pad^s1_did_read_pad; 
  assign DCache_xor22=s1_valid_pad^DCache_xor46; 
  assign DCache_xor10=DCache_xor21^DCache_xor22; 
  assign DCache_xor4=DCache_xor9^DCache_xor10; 
  assign DCache_xor1=DCache_xor3^DCache_xor4; 
  assign DCache_xor23=s2_probe_pad^s2_hit_way_pad; 
  assign DCache_xor24=s2_not_nacked_in_s1_pad^s2_probe_state_state_pad; 
  assign DCache_xor11=DCache_xor23^DCache_xor24; 
  assign DCache_xor25=s1_req_size_pad^pstore1_rmw_r_pad; 
  assign DCache_xor54=s2_valid_pad^pstore_drain_on_miss_REG_pad; 
  assign DCache_xor26=s2_release_data_valid_pad^DCache_xor54; 
  assign DCache_xor12=DCache_xor25^DCache_xor26; 
  assign DCache_xor5=DCache_xor11^DCache_xor12; 
  assign DCache_xor27=resetting_pad^grantInProgress_pad; 
  assign DCache_xor28=s2_probe_way_pad^mux_cond_0_pad; 
  assign DCache_xor13=DCache_xor27^DCache_xor28; 
  assign DCache_xor29=mux_cond_1_pad^mux_cond_2_pad; 
  assign DCache_xor62=mux_cond_4_pad^mux_cond_5_pad; 
  assign DCache_xor30=mux_cond_3_pad^DCache_xor62; 
  assign DCache_xor14=DCache_xor29^DCache_xor30; 
  assign DCache_xor6=DCache_xor13^DCache_xor14; 
  assign DCache_xor2=DCache_xor5^DCache_xor6; 
  assign DCache_xor0=DCache_xor1^DCache_xor2; 
  assign data_sum=DCache_covSum+data_io_covSum; 
  assign tlb_sum=data_sum+tlb_io_covSum; 
  assign pma_checker_sum=tlb_sum+pma_checker_io_covSum; 
  assign metaArb_sum=pma_checker_sum+metaArb_io_covSum; 
  assign lfsr_prng_sum=metaArb_sum+lfsr_prng_io_covSum; 
  assign amoalu_sum=lfsr_prng_sum+amoalu_io_covSum; 
  assign dataArb_sum=amoalu_sum+dataArb_io_covSum; 
  assign io_covSum=dataArb_sum; 
  assign stopEn0=~_dataArb_io_in_3_valid_T_54; 
  assign stopEn1=~_T_68; 
  assign stopEn2=~_dataArb_io_in_3_valid_T_54; 
  assign stopEn3=~_T_258; 
  assign stopEn4=_GEN_367&~_T_273; 
  assign stopEn5=_GEN_372&~_T_278; 
  assign stopEn6=_GEN_381&~_T_281; 
  assign stopEn7=~_T_289; 
  assign stopEn8=s2_want_victimize&~_T_301; 
  assign stopEn9=doUncachedResp&~_T_321; 
  assign lfsr_prng_metaAssert_wire=lfsr_prng_metaAssert; 
  assign tlb_metaAssert_wire=tlb_metaAssert; 
  assign amoalu_metaAssert_wire=amoalu_metaAssert; 
  assign data_metaAssert_wire=data_metaAssert; 
  assign dataArb_metaAssert_wire=dataArb_metaAssert; 
  assign pma_checker_metaAssert_wire=pma_checker_metaAssert; 
  assign metaArb_metaAssert_wire=metaArb_metaAssert; 
  assign DCache_or7=stopEn0|stopEn1; 
  assign DCache_or8=stopEn2|stopEn3; 
  assign DCache_or3=DCache_or7|DCache_or8; 
  assign DCache_or9=stopEn4|stopEn5; 
  assign DCache_or10=stopEn6|stopEn7; 
  assign DCache_or4=DCache_or9|DCache_or10; 
  assign DCache_or1=DCache_or3|DCache_or4; 
  assign DCache_or11=stopEn8|stopEn9; 
  assign DCache_or12=dataArb_metaAssert_wire|tlb_metaAssert_wire; 
  assign DCache_or5=DCache_or11|DCache_or12; 
  assign DCache_or13=amoalu_metaAssert_wire|lfsr_prng_metaAssert_wire; 
  assign DCache_or30=pma_checker_metaAssert_wire|metaArb_metaAssert_wire; 
  assign DCache_or14=data_metaAssert_wire|DCache_or30; 
  assign DCache_or6=DCache_or13|DCache_or14; 
  assign DCache_or2=DCache_or5|DCache_or6; 
  assign DCache_or0=DCache_or1|DCache_or2; 
  assign metaAssert=DCache_or0; 
  assign data_metaReset=metaReset|data_halt; 
  assign tlb_metaReset=metaReset|tlb_halt; 
  assign pma_checker_metaReset=metaReset|pma_checker_halt; 
  assign lfsr_prng_metaReset=metaReset|lfsr_prng_halt; initial
    begin 
    end  
  always @( posedge gated_clock)
       begin 
         if (tag_array_0_MPORT_en&tag_array_0_MPORT_mask)
            begin 
              tag_array_0 [tag_array_0_MPORT_addr]<=tag_array_0_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_0_s1_meta_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_0_s1_meta_en_pipe_0 <=metaArb_io_out_valid&~metaArb_io_out_bits_write;
            end 
         if (metaReset)
            begin 
              tag_array_0_s1_meta_addr_pipe_0 <=6'h0;
            end 
          else 
            if (metaArb_io_out_valid&~metaArb_io_out_bits_write)
               begin 
                 tag_array_0_s1_meta_addr_pipe_0 <=metaArb_io_out_bits_idx;
               end 
         if (tag_array_1_MPORT_en&tag_array_1_MPORT_mask)
            begin 
              tag_array_1 [tag_array_1_MPORT_addr]<=tag_array_1_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_1_s1_meta_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_1_s1_meta_en_pipe_0 <=metaArb_io_out_valid&~metaArb_io_out_bits_write;
            end 
         if (metaReset)
            begin 
              tag_array_1_s1_meta_addr_pipe_0 <=6'h0;
            end 
          else 
            if (metaArb_io_out_valid&~metaArb_io_out_bits_write)
               begin 
                 tag_array_1_s1_meta_addr_pipe_0 <=metaArb_io_out_bits_idx;
               end 
         if (tag_array_2_MPORT_en&tag_array_2_MPORT_mask)
            begin 
              tag_array_2 [tag_array_2_MPORT_addr]<=tag_array_2_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_2_s1_meta_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_2_s1_meta_en_pipe_0 <=metaArb_io_out_valid&~metaArb_io_out_bits_write;
            end 
         if (metaReset)
            begin 
              tag_array_2_s1_meta_addr_pipe_0 <=6'h0;
            end 
          else 
            if (metaArb_io_out_valid&~metaArb_io_out_bits_write)
               begin 
                 tag_array_2_s1_meta_addr_pipe_0 <=metaArb_io_out_bits_idx;
               end 
         if (tag_array_3_MPORT_en&tag_array_3_MPORT_mask)
            begin 
              tag_array_3 [tag_array_3_MPORT_addr]<=tag_array_3_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_3_s1_meta_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_3_s1_meta_en_pipe_0 <=metaArb_io_out_valid&~metaArb_io_out_bits_write;
            end 
         if (metaReset)
            begin 
              tag_array_3_s1_meta_addr_pipe_0 <=6'h0;
            end 
          else 
            if (metaArb_io_out_valid&~metaArb_io_out_bits_write)
               begin 
                 tag_array_3_s1_meta_addr_pipe_0 <=metaArb_io_out_bits_idx;
               end 
         if (metaReset)
            begin 
              s1_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s1_valid <=1'h0;
               end 
             else 
               begin 
                 s1_valid <=s1_valid_x9;
               end 
         if (metaReset)
            begin 
              blockProbeAfterGrantCount <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 blockProbeAfterGrantCount <=3'h0;
               end 
             else 
               if (_T_271)
                  begin 
                    if (grantIsCached)
                       begin 
                         if (d_last)
                            begin 
                              blockProbeAfterGrantCount <=3'h7;
                            end 
                          else 
                            if (_block_probe_for_core_progress_T)
                               begin 
                                 blockProbeAfterGrantCount <=_blockProbeAfterGrantCount_T_1;
                               end 
                       end 
                     else 
                       if (_block_probe_for_core_progress_T)
                          begin 
                            blockProbeAfterGrantCount <=_blockProbeAfterGrantCount_T_1;
                          end 
                  end 
                else 
                  if (_block_probe_for_core_progress_T)
                     begin 
                       blockProbeAfterGrantCount <=_blockProbeAfterGrantCount_T_1;
                     end 
         if (metaReset)
            begin 
              lrscCount <=7'h0;
            end 
          else 
            if (reset)
               begin 
                 lrscCount <=7'h0;
               end 
             else 
               if (s1_probe)
                  begin 
                    lrscCount <=7'h0;
                  end 
                else 
                  if (_T_250)
                     begin 
                       lrscCount <=7'h3;
                     end 
                   else 
                     if (_lrscBackingOff_T)
                        begin 
                          lrscCount <=_lrscCount_T_2;
                        end 
                      else 
                        if (_T_246)
                           begin 
                             if (s2_hit)
                                begin 
                                  lrscCount <=7'h4f;
                                end 
                              else 
                                begin 
                                  lrscCount <=7'h0;
                                end 
                           end 
         if (metaReset)
            begin 
              s1_probe <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s1_probe <=1'h0;
               end 
             else 
               if (_T_304)
                  begin 
                    s1_probe <=_GEN_295;
                  end 
                else 
                  begin 
                    s1_probe <=s1_probe_x12;
                  end 
         if (metaReset)
            begin 
              s2_probe <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s2_probe <=1'h0;
               end 
             else 
               begin 
                 s2_probe <=s1_probe;
               end 
         if (metaReset)
            begin 
              release_state <=4'h0;
            end 
          else 
            if (reset)
               begin 
                 release_state <=4'h0;
               end 
             else 
               if (_T_316)
                  begin 
                    release_state <=4'h0;
                  end 
                else 
                  if (_T_312)
                     begin 
                       if (releaseDone)
                          begin 
                            release_state <=4'h6;
                          end 
                        else 
                          if (_T_307)
                             begin 
                               if (releaseDone)
                                  begin 
                                    release_state <=4'h7;
                                  end 
                                else 
                                  if (_T_306)
                                     begin 
                                       if (releaseDone)
                                          begin 
                                            release_state <=4'h7;
                                          end 
                                        else 
                                          if (_T_305)
                                             begin 
                                               if (releaseDone)
                                                  begin 
                                                    release_state <=4'h0;
                                                  end 
                                                else 
                                                  if (_T_304)
                                                     begin 
                                                       if (metaArb_io_in_6_ready)
                                                          begin 
                                                            release_state <=4'h0;
                                                          end 
                                                        else 
                                                          if (s2_probe)
                                                             begin 
                                                               if (s2_meta_error)
                                                                  begin 
                                                                    release_state <=4'h4;
                                                                  end 
                                                                else 
                                                                  if (s2_prb_ack_data)
                                                                     begin 
                                                                       release_state <=4'h2;
                                                                     end 
                                                                   else 
                                                                     if (_T_303)
                                                                        begin 
                                                                          if (releaseDone)
                                                                             begin 
                                                                               release_state <=4'h7;
                                                                             end 
                                                                           else 
                                                                             begin 
                                                                               release_state <=4'h3;
                                                                             end 
                                                                        end 
                                                                      else 
                                                                        if (releaseDone)
                                                                           begin 
                                                                             release_state <=4'h0;
                                                                           end 
                                                                         else 
                                                                           begin 
                                                                             release_state <=4'h5;
                                                                           end 
                                                             end 
                                                           else 
                                                             if (s2_want_victimize)
                                                                begin 
                                                                  if (_release_state_T_1)
                                                                     begin 
                                                                       release_state <=4'h1;
                                                                     end 
                                                                   else 
                                                                     begin 
                                                                       release_state <=4'h6;
                                                                     end 
                                                                end 
                                                     end 
                                                   else 
                                                     if (s2_probe)
                                                        begin 
                                                          if (s2_meta_error)
                                                             begin 
                                                               release_state <=4'h4;
                                                             end 
                                                           else 
                                                             if (s2_prb_ack_data)
                                                                begin 
                                                                  release_state <=4'h2;
                                                                end 
                                                              else 
                                                                if (_T_303)
                                                                   begin 
                                                                     if (releaseDone)
                                                                        begin 
                                                                          release_state <=4'h7;
                                                                        end 
                                                                      else 
                                                                        begin 
                                                                          release_state <=4'h3;
                                                                        end 
                                                                   end 
                                                                 else 
                                                                   if (releaseDone)
                                                                      begin 
                                                                        release_state <=4'h0;
                                                                      end 
                                                                    else 
                                                                      begin 
                                                                        release_state <=4'h5;
                                                                      end 
                                                        end 
                                                      else 
                                                        if (s2_want_victimize)
                                                           begin 
                                                             if (_release_state_T_1)
                                                                begin 
                                                                  release_state <=4'h1;
                                                                end 
                                                              else 
                                                                begin 
                                                                  release_state <=4'h6;
                                                                end 
                                                           end 
                                             end 
                                           else 
                                             if (_T_304)
                                                begin 
                                                  if (metaArb_io_in_6_ready)
                                                     begin 
                                                       release_state <=4'h0;
                                                     end 
                                                   else 
                                                     if (s2_probe)
                                                        begin 
                                                          if (s2_meta_error)
                                                             begin 
                                                               release_state <=4'h4;
                                                             end 
                                                           else 
                                                             if (s2_prb_ack_data)
                                                                begin 
                                                                  release_state <=4'h2;
                                                                end 
                                                              else 
                                                                if (_T_303)
                                                                   begin 
                                                                     if (releaseDone)
                                                                        begin 
                                                                          release_state <=4'h7;
                                                                        end 
                                                                      else 
                                                                        begin 
                                                                          release_state <=4'h3;
                                                                        end 
                                                                   end 
                                                                 else 
                                                                   if (releaseDone)
                                                                      begin 
                                                                        release_state <=4'h0;
                                                                      end 
                                                                    else 
                                                                      begin 
                                                                        release_state <=4'h5;
                                                                      end 
                                                        end 
                                                      else 
                                                        if (s2_want_victimize)
                                                           begin 
                                                             if (_release_state_T_1)
                                                                begin 
                                                                  release_state <=4'h1;
                                                                end 
                                                              else 
                                                                begin 
                                                                  release_state <=4'h6;
                                                                end 
                                                           end 
                                                end 
                                              else 
                                                if (s2_probe)
                                                   begin 
                                                     if (s2_meta_error)
                                                        begin 
                                                          release_state <=4'h4;
                                                        end 
                                                      else 
                                                        if (s2_prb_ack_data)
                                                           begin 
                                                             release_state <=4'h2;
                                                           end 
                                                         else 
                                                           if (_T_303)
                                                              begin 
                                                                if (releaseDone)
                                                                   begin 
                                                                     release_state <=4'h7;
                                                                   end 
                                                                 else 
                                                                   begin 
                                                                     release_state <=4'h3;
                                                                   end 
                                                              end 
                                                            else 
                                                              if (releaseDone)
                                                                 begin 
                                                                   release_state <=4'h0;
                                                                 end 
                                                               else 
                                                                 begin 
                                                                   release_state <=4'h5;
                                                                 end 
                                                   end 
                                                 else 
                                                   if (s2_want_victimize)
                                                      begin 
                                                        if (_release_state_T_1)
                                                           begin 
                                                             release_state <=4'h1;
                                                           end 
                                                         else 
                                                           begin 
                                                             release_state <=4'h6;
                                                           end 
                                                      end 
                                     end 
                                   else 
                                     if (_T_305)
                                        begin 
                                          if (releaseDone)
                                             begin 
                                               release_state <=4'h0;
                                             end 
                                           else 
                                             if (_T_304)
                                                begin 
                                                  if (metaArb_io_in_6_ready)
                                                     begin 
                                                       release_state <=4'h0;
                                                     end 
                                                   else 
                                                     begin 
                                                       release_state <=_GEN_284;
                                                     end 
                                                end 
                                              else 
                                                begin 
                                                  release_state <=_GEN_284;
                                                end 
                                        end 
                                      else 
                                        if (_T_304)
                                           begin 
                                             if (metaArb_io_in_6_ready)
                                                begin 
                                                  release_state <=4'h0;
                                                end 
                                              else 
                                                begin 
                                                  release_state <=_GEN_284;
                                                end 
                                           end 
                                         else 
                                           begin 
                                             release_state <=_GEN_284;
                                           end 
                             end 
                           else 
                             if (_T_306)
                                begin 
                                  if (releaseDone)
                                     begin 
                                       release_state <=4'h7;
                                     end 
                                   else 
                                     if (_T_305)
                                        begin 
                                          if (releaseDone)
                                             begin 
                                               release_state <=4'h0;
                                             end 
                                           else 
                                             begin 
                                               release_state <=_GEN_299;
                                             end 
                                        end 
                                      else 
                                        begin 
                                          release_state <=_GEN_299;
                                        end 
                                end 
                              else 
                                if (_T_305)
                                   begin 
                                     if (releaseDone)
                                        begin 
                                          release_state <=4'h0;
                                        end 
                                      else 
                                        begin 
                                          release_state <=_GEN_299;
                                        end 
                                   end 
                                 else 
                                   begin 
                                     release_state <=_GEN_299;
                                   end 
                     end 
                   else 
                     if (_T_307)
                        begin 
                          if (releaseDone)
                             begin 
                               release_state <=4'h7;
                             end 
                           else 
                             if (_T_306)
                                begin 
                                  if (releaseDone)
                                     begin 
                                       release_state <=4'h7;
                                     end 
                                   else 
                                     begin 
                                       release_state <=_GEN_303;
                                     end 
                                end 
                              else 
                                begin 
                                  release_state <=_GEN_303;
                                end 
                        end 
                      else 
                        if (_T_306)
                           begin 
                             if (releaseDone)
                                begin 
                                  release_state <=4'h7;
                                end 
                              else 
                                begin 
                                  release_state <=_GEN_303;
                                end 
                           end 
                         else 
                           begin 
                             release_state <=_GEN_303;
                           end 
         if (metaReset)
            begin 
              release_ack_wait <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 release_ack_wait <=1'h0;
               end 
             else 
               if (_T_312)
                  begin 
                    release_ack_wait <=_GEN_331;
                  end 
                else 
                  if (_T_271)
                     begin 
                       if (!(grantIsCached))
                          begin 
                            if (!(grantIsUncached))
                               begin 
                                 if (grantIsVoluntary)
                                    begin 
                                      release_ack_wait <=1'h0;
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              release_ack_addr <=32'h0;
            end 
          else 
            if (_T_312)
               begin 
                 if (_T_315)
                    begin 
                      release_ack_addr <=probe_bits_address;
                    end 
               end 
         if (metaReset)
            begin 
              grantInProgress <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 grantInProgress <=1'h0;
               end 
             else 
               if (_T_271)
                  begin 
                    if (grantIsCached)
                       begin 
                         if (d_last)
                            begin 
                              grantInProgress <=1'h0;
                            end 
                          else 
                            begin 
                              grantInProgress <=1'h1;
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              s2_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s2_valid <=1'h0;
               end 
             else 
               begin 
                 s2_valid <=s2_valid_x37;
               end 
         if (metaReset)
            begin 
              probe_bits_param <=2'h0;
            end 
          else 
            if (s2_want_victimize)
               begin 
                 probe_bits_param <=2'h0;
               end 
             else 
               if (s1_probe_x12)
                  begin 
                    probe_bits_param <=auto_out_b_bits_param;
                  end 
         if (metaReset)
            begin 
              probe_bits_size <=4'h0;
            end 
          else 
            if (s2_want_victimize)
               begin 
                 probe_bits_size <=4'h0;
               end 
             else 
               if (s1_probe_x12)
                  begin 
                    probe_bits_size <=auto_out_b_bits_size;
                  end 
         if (metaReset)
            begin 
              probe_bits_source <=1'h0;
            end 
          else 
            if (s2_want_victimize)
               begin 
                 probe_bits_source <=1'h0;
               end 
             else 
               if (s1_probe_x12)
                  begin 
                    probe_bits_source <=auto_out_b_bits_source;
                  end 
         if (metaReset)
            begin 
              probe_bits_address <=32'h0;
            end 
          else 
            if (s2_want_victimize)
               begin 
                 probe_bits_address <=res_2_address;
               end 
             else 
               if (s1_probe_x12)
                  begin 
                    probe_bits_address <=auto_out_b_bits_address;
                  end 
         if (metaReset)
            begin 
              s2_probe_state_state <=2'h0;
            end 
          else 
            if (s1_probe)
               begin 
                 s2_probe_state_state <=s1_meta_hit_state_state;
               end 
         if (metaReset)
            begin 
              counter_1 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 counter_1 <=9'h0;
               end 
             else 
               if (_T_297)
                  begin 
                    if (c_first)
                       begin 
                         if (beats1_opdata_1)
                            begin 
                              counter_1 <=beats1_decode_1;
                            end 
                          else 
                            begin 
                              counter_1 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         counter_1 <=counter1_1;
                       end 
                  end 
         if (metaReset)
            begin 
              s2_release_data_valid <=1'h0;
            end 
          else 
            begin 
              s2_release_data_valid <=s1_release_data_valid&~releaseRejected;
            end 
         if (metaReset)
            begin 
              s1_req_cmd <=5'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_req_cmd <=io_cpu_req_bits_cmd;
               end 
         if (metaReset)
            begin 
              s2_req_cmd <=5'h0;
            end 
          else 
            if (_T_271)
               begin 
                 if (grantIsCached)
                    begin 
                      if (_T_70)
                         begin 
                           s2_req_cmd <=s1_req_cmd;
                         end 
                    end 
                  else 
                    if (grantIsUncached)
                       begin 
                         if (grantIsUncachedData)
                            begin 
                              s2_req_cmd <=5'h0;
                            end 
                          else 
                            if (_T_70)
                               begin 
                                 s2_req_cmd <=s1_req_cmd;
                               end 
                       end 
                     else 
                       if (_T_70)
                          begin 
                            s2_req_cmd <=s1_req_cmd;
                          end 
               end 
             else 
               if (_T_70)
                  begin 
                    s2_req_cmd <=s1_req_cmd;
                  end 
         if (metaReset)
            begin 
              pstore1_held <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 pstore1_held <=1'h0;
               end 
             else 
               begin 
                 pstore1_held <=_pstore1_held_T_10;
               end 
         if (metaReset)
            begin 
              pstore1_addr <=40'h0;
            end 
          else 
            if (_pstore1_cmd_T)
               begin 
                 pstore1_addr <=s1_vaddr;
               end 
         if (metaReset)
            begin 
              s1_req_addr <=40'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_req_addr <=s0_req_addr;
               end 
         if (metaReset)
            begin 
              pstore1_mask <=8'h0;
            end 
          else 
            if (_pstore1_cmd_T)
               begin 
                 if (_s1_write_T_1)
                    begin 
                      pstore1_mask <=8'h0;
                    end 
                  else 
                    begin 
                      pstore1_mask <=s1_mask_xwr;
                    end 
               end 
         if (metaReset)
            begin 
              s1_req_size <=2'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_req_size <=io_cpu_req_bits_size;
               end 
         if (metaReset)
            begin 
              pstore2_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 pstore2_valid <=1'h0;
               end 
             else 
               begin 
                 pstore2_valid <=_pstore2_valid_T_2;
               end 
         if (metaReset)
            begin 
              pstore2_addr <=40'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_addr <=pstore1_addr;
               end 
         if (metaReset)
            begin 
              mask <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 mask <=pstore1_mask[7:0];
               end 
         if (metaReset)
            begin 
              s2_not_nacked_in_s1 <=1'h0;
            end 
          else 
            begin 
              s2_not_nacked_in_s1 <=~s1_nack;
            end 
         if (metaReset)
            begin 
              s2_hit_state_state <=2'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_hit_state_state <=s1_meta_hit_state_state;
               end 
         if (metaReset)
            begin 
              s1_req_tag <=7'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_req_tag <=io_cpu_req_bits_tag;
               end 
         if (metaReset)
            begin 
              s1_req_signed <=1'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_req_signed <=io_cpu_req_bits_signed;
               end 
         if (metaReset)
            begin 
              s1_tlb_req_vaddr <=40'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_tlb_req_vaddr <=s0_req_addr;
               end 
         if (metaReset)
            begin 
              s1_tlb_req_passthrough <=1'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_tlb_req_passthrough <=s0_req_phys;
               end 
         if (metaReset)
            begin 
              s1_tlb_req_size <=2'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_tlb_req_size <=io_cpu_req_bits_size;
               end 
         if (metaReset)
            begin 
              s1_tlb_req_cmd <=5'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_tlb_req_cmd <=io_cpu_req_bits_cmd;
               end 
         if (metaReset)
            begin 
              s1_flush_valid <=1'h0;
            end 
          else 
            begin 
              s1_flush_valid <=_s1_flush_valid_T_6&~release_ack_wait;
            end 
         if (metaReset)
            begin 
              cached_grant_wait <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 cached_grant_wait <=1'h0;
               end 
             else 
               if (_T_271)
                  begin 
                    if (grantIsCached)
                       begin 
                         if (d_last)
                            begin 
                              cached_grant_wait <=1'h0;
                            end 
                          else 
                            if (_T_263)
                               begin 
                                 if (!(s2_uncached))
                                    begin 
                                      cached_grant_wait <=1'h1;
                                    end 
                               end 
                       end 
                     else 
                       if (_T_263)
                          begin 
                            if (!(s2_uncached))
                               begin 
                                 cached_grant_wait <=1'h1;
                               end 
                          end 
                  end 
                else 
                  if (_T_263)
                     begin 
                       if (!(s2_uncached))
                          begin 
                            cached_grant_wait <=1'h1;
                          end 
                     end 
         if (metaReset)
            begin 
              resetting <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 resetting <=1'h0;
               end 
             else 
               if (resetting)
                  begin 
                    if (flushDone)
                       begin 
                         resetting <=1'h0;
                       end 
                     else 
                       begin 
                         resetting <=_GEN_349;
                       end 
                  end 
                else 
                  begin 
                    resetting <=_GEN_349;
                  end 
         if (metaReset)
            begin 
              flushCounter <=8'h0;
            end 
          else 
            if (reset)
               begin 
                 flushCounter <=8'hc0;
               end 
             else 
               begin 
                 flushCounter <=_GEN_351[7:0];
               end 
         if (metaReset)
            begin 
              refill_way <=4'h0;
            end 
          else 
            if (_T_263)
               begin 
                 if (!(s2_uncached))
                    begin 
                      if (s2_hit_valid)
                         begin 
                           refill_way <=s2_hit_way;
                         end 
                       else 
                         begin 
                           refill_way <=s2_victim_way;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              uncachedInFlight_0 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 uncachedInFlight_0 <=1'h0;
               end 
             else 
               if (_T_271)
                  begin 
                    if (grantIsCached)
                       begin 
                         if (_T_263)
                            begin 
                              if (s2_uncached)
                                 begin 
                                   uncachedInFlight_0 <=_GEN_142;
                                 end 
                            end 
                       end 
                     else 
                       if (grantIsUncached)
                          begin 
                            if (_T_276)
                               begin 
                                 uncachedInFlight_0 <=1'h0;
                               end 
                             else 
                               if (_T_263)
                                  begin 
                                    if (s2_uncached)
                                       begin 
                                         uncachedInFlight_0 <=_GEN_142;
                                       end 
                                  end 
                          end 
                        else 
                          if (_T_263)
                             begin 
                               if (s2_uncached)
                                  begin 
                                    uncachedInFlight_0 <=_GEN_142;
                                  end 
                             end 
                  end 
                else 
                  if (_T_263)
                     begin 
                       if (s2_uncached)
                          begin 
                            uncachedInFlight_0 <=_GEN_142;
                          end 
                     end 
         if (metaReset)
            begin 
              uncachedReqs_0_addr <=40'h0;
            end 
          else 
            if (_T_263)
               begin 
                 if (s2_uncached)
                    begin 
                      if (a_sel)
                         begin 
                           uncachedReqs_0_addr <=s2_req_addr;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              uncachedReqs_0_tag <=7'h0;
            end 
          else 
            if (_T_263)
               begin 
                 if (s2_uncached)
                    begin 
                      if (a_sel)
                         begin 
                           uncachedReqs_0_tag <=s2_req_tag;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              uncachedReqs_0_size <=2'h0;
            end 
          else 
            if (_T_263)
               begin 
                 if (s2_uncached)
                    begin 
                      if (a_sel)
                         begin 
                           uncachedReqs_0_size <=s2_req_size;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              uncachedReqs_0_signed <=1'h0;
            end 
          else 
            if (_T_263)
               begin 
                 if (s2_uncached)
                    begin 
                      if (a_sel)
                         begin 
                           uncachedReqs_0_signed <=s2_req_signed;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              s1_did_read <=1'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_did_read <=_s1_did_read_T_52;
               end 
         if (metaReset)
            begin 
              s1_read_mask <=1'h0;
            end 
          else 
            if (s0_clk_en)
               begin 
                 s1_read_mask <=dataArb_io_in_3_bits_wordMask;
               end 
         if (metaReset)
            begin 
              s2_hit_way <=4'h0;
            end 
          else 
            if (s1_valid_not_nacked)
               begin 
                 s2_hit_way <=s1_meta_hit_way;
               end 
         if (metaReset)
            begin 
              s2_victim_way_r <=2'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_victim_way_r <=s1_victim_way;
               end 
         if (metaReset)
            begin 
              s2_probe_way <=4'h0;
            end 
          else 
            if (s1_probe)
               begin 
                 s2_probe_way <=s1_meta_hit_way;
               end 
         if (metaReset)
            begin 
              s2_req_addr <=40'h0;
            end 
          else 
            if (_T_271)
               begin 
                 if (grantIsCached)
                    begin 
                      if (_T_70)
                         begin 
                           s2_req_addr <={8'b0,s1_paddr};
                         end 
                    end 
                  else 
                    if (grantIsUncached)
                       begin 
                         if (grantIsUncachedData)
                            begin 
                              s2_req_addr <={8'b0,_s2_req_addr_T_1};
                            end 
                          else 
                            if (_T_70)
                               begin 
                                 s2_req_addr <={8'b0,s1_paddr};
                               end 
                       end 
                     else 
                       if (_T_70)
                          begin 
                            s2_req_addr <={8'b0,s1_paddr};
                          end 
               end 
             else 
               if (_T_70)
                  begin 
                    s2_req_addr <={8'b0,s1_paddr};
                  end 
         if (metaReset)
            begin 
              s2_req_tag <=7'h0;
            end 
          else 
            if (_T_271)
               begin 
                 if (grantIsCached)
                    begin 
                      if (_T_70)
                         begin 
                           s2_req_tag <=s1_req_tag;
                         end 
                    end 
                  else 
                    if (grantIsUncached)
                       begin 
                         if (grantIsUncachedData)
                            begin 
                              s2_req_tag <=uncachedReqs_0_tag;
                            end 
                          else 
                            if (_T_70)
                               begin 
                                 s2_req_tag <=s1_req_tag;
                               end 
                       end 
                     else 
                       if (_T_70)
                          begin 
                            s2_req_tag <=s1_req_tag;
                          end 
               end 
             else 
               if (_T_70)
                  begin 
                    s2_req_tag <=s1_req_tag;
                  end 
         if (metaReset)
            begin 
              s2_req_size <=2'h0;
            end 
          else 
            if (_T_271)
               begin 
                 if (grantIsCached)
                    begin 
                      if (_T_70)
                         begin 
                           s2_req_size <=s1_req_size;
                         end 
                    end 
                  else 
                    if (grantIsUncached)
                       begin 
                         if (grantIsUncachedData)
                            begin 
                              s2_req_size <=uncachedReqs_0_size;
                            end 
                          else 
                            if (_T_70)
                               begin 
                                 s2_req_size <=s1_req_size;
                               end 
                       end 
                     else 
                       if (_T_70)
                          begin 
                            s2_req_size <=s1_req_size;
                          end 
               end 
             else 
               if (_T_70)
                  begin 
                    s2_req_size <=s1_req_size;
                  end 
         if (metaReset)
            begin 
              s2_req_signed <=1'h0;
            end 
          else 
            if (_T_271)
               begin 
                 if (grantIsCached)
                    begin 
                      if (_T_70)
                         begin 
                           s2_req_signed <=s1_req_signed;
                         end 
                    end 
                  else 
                    if (grantIsUncached)
                       begin 
                         if (grantIsUncachedData)
                            begin 
                              s2_req_signed <=uncachedReqs_0_signed;
                            end 
                          else 
                            if (_T_70)
                               begin 
                                 s2_req_signed <=s1_req_signed;
                               end 
                       end 
                     else 
                       if (_T_70)
                          begin 
                            s2_req_signed <=s1_req_signed;
                          end 
               end 
             else 
               if (_T_70)
                  begin 
                    s2_req_signed <=s1_req_signed;
                  end 
         if (metaReset)
            begin 
              s2_tlb_xcpt_pf_ld <=1'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_tlb_xcpt_pf_ld <=tlb_io_resp_pf_ld;
               end 
         if (metaReset)
            begin 
              s2_tlb_xcpt_pf_st <=1'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_tlb_xcpt_pf_st <=tlb_io_resp_pf_st;
               end 
         if (metaReset)
            begin 
              s2_tlb_xcpt_ae_ld <=1'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_tlb_xcpt_ae_ld <=tlb_io_resp_ae_ld;
               end 
         if (metaReset)
            begin 
              s2_tlb_xcpt_ae_st <=1'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_tlb_xcpt_ae_st <=tlb_io_resp_ae_st;
               end 
         if (metaReset)
            begin 
              s2_tlb_xcpt_ma_ld <=1'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_tlb_xcpt_ma_ld <=tlb_io_resp_ma_ld;
               end 
         if (metaReset)
            begin 
              s2_tlb_xcpt_ma_st <=1'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_tlb_xcpt_ma_st <=tlb_io_resp_ma_st;
               end 
         if (metaReset)
            begin 
              s2_pma_cacheable <=1'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_pma_cacheable <=_s2_pma_T_cacheable;
               end 
         if (metaReset)
            begin 
              s2_vaddr_r <=40'h0;
            end 
          else 
            if (_T_70)
               begin 
                 s2_vaddr_r <=s1_vaddr;
               end 
         if (metaReset)
            begin 
              s2_flush_valid_pre_tag_ecc <=1'h0;
            end 
          else 
            begin 
              s2_flush_valid_pre_tag_ecc <=s1_flush_valid;
            end 
         if (metaReset)
            begin 
              s2_meta_corrected_r <=22'h0;
            end 
          else 
            if (s1_meta_clk_en)
               begin 
                 s2_meta_corrected_r <=tag_array_0_s1_meta_data;
               end 
         if (metaReset)
            begin 
              s2_meta_corrected_r_1 <=22'h0;
            end 
          else 
            if (s1_meta_clk_en)
               begin 
                 s2_meta_corrected_r_1 <=tag_array_1_s1_meta_data;
               end 
         if (metaReset)
            begin 
              s2_meta_corrected_r_2 <=22'h0;
            end 
          else 
            if (s1_meta_clk_en)
               begin 
                 s2_meta_corrected_r_2 <=tag_array_2_s1_meta_data;
               end 
         if (metaReset)
            begin 
              s2_meta_corrected_r_3 <=22'h0;
            end 
          else 
            if (s1_meta_clk_en)
               begin 
                 s2_meta_corrected_r_3 <=tag_array_3_s1_meta_data;
               end 
         if (metaReset)
            begin 
              blockUncachedGrant <=1'h0;
            end 
          else 
            if (_T_294)
               begin 
                 if (auto_out_d_valid)
                    begin 
                      blockUncachedGrant <=~dataArb_io_in_1_ready;
                    end 
                  else 
                    begin 
                      blockUncachedGrant <=dataArb_io_out_valid;
                    end 
               end 
             else 
               begin 
                 blockUncachedGrant <=dataArb_io_out_valid;
               end 
         if (metaReset)
            begin 
              counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 counter <=9'h0;
               end 
             else 
               if (_T_271)
                  begin 
                    if (d_first)
                       begin 
                         if (beats1_opdata)
                            begin 
                              counter <=beats1_decode;
                            end 
                          else 
                            begin 
                              counter <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         counter <=counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              s2_data <=64'h0;
            end 
          else 
            if (en)
               begin 
                 s2_data <=_s2_data_T_15;
               end 
         if (metaReset)
            begin 
              lrscAddr <=34'h0;
            end 
          else 
            if (_T_246)
               begin 
                 lrscAddr <=s2_req_addr[39:6];
               end 
         if (metaReset)
            begin 
              pstore1_cmd <=5'h0;
            end 
          else 
            if (_pstore1_cmd_T)
               begin 
                 pstore1_cmd <=s1_req_cmd;
               end 
         if (metaReset)
            begin 
              pstore1_data <=64'h0;
            end 
          else 
            if (_pstore1_cmd_T)
               begin 
                 pstore1_data <=io_cpu_s1_data_data;
               end 
         if (metaReset)
            begin 
              pstore1_way <=4'h0;
            end 
          else 
            if (_pstore1_cmd_T)
               begin 
                 pstore1_way <=s1_meta_hit_way;
               end 
         if (metaReset)
            begin 
              pstore1_rmw_r <=1'h0;
            end 
          else 
            if (_pstore1_cmd_T)
               begin 
                 pstore1_rmw_r <=_pstore1_rmw_T_50;
               end 
         if (metaReset)
            begin 
              pstore_drain_on_miss_REG <=1'h0;
            end 
          else 
            begin 
              pstore_drain_on_miss_REG <=io_cpu_s2_nack;
            end 
         if (metaReset)
            begin 
              pstore2_way <=4'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_way <=pstore1_way;
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_lo_lo_lo <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_lo_lo_lo <=pstore1_storegen_data[7:0];
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_lo_lo_hi <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_lo_lo_hi <=pstore1_storegen_data[15:8];
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_lo_hi_lo <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_lo_hi_lo <=pstore1_storegen_data[23:16];
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_lo_hi_hi <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_lo_hi_hi <=pstore1_storegen_data[31:24];
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_hi_lo_lo <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_hi_lo_lo <=pstore1_storegen_data[39:32];
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_hi_lo_hi <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_hi_lo_hi <=pstore1_storegen_data[47:40];
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_hi_hi_lo <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_hi_hi_lo <=pstore1_storegen_data[55:48];
               end 
         if (metaReset)
            begin 
              pstore2_storegen_data_hi_hi_hi <=8'h0;
            end 
          else 
            if (advance_pstore1)
               begin 
                 pstore2_storegen_data_hi_hi_hi <=pstore1_storegen_data[63:56];
               end 
         if (metaReset)
            begin 
              s1_release_data_valid <=1'h0;
            end 
          else 
            begin 
              s1_release_data_valid <=dataArb_io_in_2_ready&dataArb_io_in_2_valid;
            end 
         if (metaReset)
            begin 
              io_cpu_s2_xcpt_REG <=1'h0;
            end 
          else 
            begin 
              io_cpu_s2_xcpt_REG <=_s1_xcpt_valid_T_1&~s1_nack;
            end 
         if (metaReset)
            begin 
              doUncachedResp <=1'h0;
            end 
          else 
            begin 
              doUncachedResp <=io_cpu_replay_next;
            end 
         if (metaReset)
            begin 
              REG <=1'h0;
            end 
          else 
            begin 
              REG <=reset;
            end 
         if (metaReset)
            begin 
              io_cpu_perf_release_counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 io_cpu_perf_release_counter <=9'h0;
               end 
             else 
               if (_T_297)
                  begin 
                    if (io_cpu_perf_release_first)
                       begin 
                         if (beats1_opdata_1)
                            begin 
                              io_cpu_perf_release_counter <=beats1_decode_1;
                            end 
                          else 
                            begin 
                              io_cpu_perf_release_counter <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         io_cpu_perf_release_counter <=io_cpu_perf_release_counter1;
                       end 
                  end 
         if (~_dataArb_io_in_3_valid_T_54)
            begin $display("Assertion failed\n    at DCache.scala:1154 assert(!needsRead(req) || res)\n");
            end 
         if (~_dataArb_io_in_3_valid_T_54)
            begin $display("fatal");
            end 
         if (~_T_68)
            begin $display("Assertion failed\n    at DCache.scala:300 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n");
            end 
         if (~_T_68)
            begin $display("fatal");
            end 
         if (~_dataArb_io_in_3_valid_T_54)
            begin $display("Assertion failed\n    at DCache.scala:1154 assert(!needsRead(req) || res)\n");
            end 
         if (~_dataArb_io_in_3_valid_T_54)
            begin $display("fatal");
            end 
         if (~_T_258)
            begin $display("Assertion failed\n    at DCache.scala:481 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n");
            end 
         if (~_T_258)
            begin $display("fatal");
            end 
         if (_GEN_367&~_T_273)
            begin $display("Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:648 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n");
            end 
         if (_GEN_367&~_T_273)
            begin $display("fatal");
            end 
         if (_GEN_372&~_T_278)
            begin $display("Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:658 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n");
            end 
         if (_GEN_372&~_T_278)
            begin $display("fatal");
            end 
         if (_GEN_381&~_T_281)
            begin $display("Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:679 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n");
            end 
         if (_GEN_381&~_T_281)
            begin $display("fatal");
            end 
         if (~_T_289)
            begin $display("Assertion failed\n    at DCache.scala:687 assert(tl_out.e.fire() === (tl_out.d.fire() && d_first && grantIsCached))\n");
            end 
         if (~_T_289)
            begin $display("fatal");
            end 
         if (s2_want_victimize&~_T_301)
            begin $display("Assertion failed\n    at DCache.scala:788 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n");
            end 
         if (s2_want_victimize&~_T_301)
            begin $display("fatal");
            end 
         if (doUncachedResp&~_T_321)
            begin $display("Assertion failed\n    at DCache.scala:920 assert(!s2_valid_hit)\n");
            end 
         if (doUncachedResp&~_T_321)
            begin $display("fatal");
            end 
         DCache_state <=DCache_xor0;
         if (!(DCache_cov_read_data))
            begin 
              DCache_covSum <=DCache_covSum+1'h1;
            end 
       end
  
  always @( posedge gated_clock)
       begin 
         if (DCache_cov_write_en&DCache_cov_write_mask)
            begin 
              DCache_cov [DCache_cov_write_addr]<=DCache_cov_write_data;
            end 
       end
  
endmodule
 
module Frontend (
  input gated_clock,
  input reset,
  input auto_icache_master_out_a_ready,
  output auto_icache_master_out_a_valid,
  output [31:0] auto_icache_master_out_a_bits_address,
  input auto_icache_master_out_d_valid,
  input [2:0] auto_icache_master_out_d_bits_opcode,
  input [3:0] auto_icache_master_out_d_bits_size,
  input [63:0] auto_icache_master_out_d_bits_data,
  input auto_icache_master_out_d_bits_corrupt,
  input [31:0] auto_reset_vector_sink_in,
  input io_cpu_might_request,
  input io_cpu_req_valid,
  input [39:0] io_cpu_req_bits_pc,
  input io_cpu_req_bits_speculative,
  input io_cpu_sfence_valid,
  input io_cpu_sfence_bits_rs1,
  input io_cpu_sfence_bits_rs2,
  input [38:0] io_cpu_sfence_bits_addr,
  input io_cpu_resp_ready,
  output io_cpu_resp_valid,
  output io_cpu_resp_bits_btb_taken,
  output io_cpu_resp_bits_btb_bridx,
  output [4:0] io_cpu_resp_bits_btb_entry,
  output [7:0] io_cpu_resp_bits_btb_bht_history,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output io_cpu_resp_bits_xcpt_pf_inst,
  output io_cpu_resp_bits_xcpt_ae_inst,
  output io_cpu_resp_bits_replay,
  input io_cpu_btb_update_valid,
  input [4:0] io_cpu_btb_update_bits_prediction_entry,
  input [38:0] io_cpu_btb_update_bits_pc,
  input io_cpu_btb_update_bits_isValid,
  input [38:0] io_cpu_btb_update_bits_br_pc,
  input [1:0] io_cpu_btb_update_bits_cfiType,
  input io_cpu_bht_update_valid,
  input [7:0] io_cpu_bht_update_bits_prediction_history,
  input [38:0] io_cpu_bht_update_bits_pc,
  input io_cpu_bht_update_bits_branch,
  input io_cpu_bht_update_bits_taken,
  input io_cpu_bht_update_bits_mispredict,
  input io_cpu_flush_icache,
  output [39:0] io_cpu_npc,
  input io_ptw_req_ready,
  output io_ptw_req_valid,
  output io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input io_ptw_resp_valid,
  input io_ptw_resp_bits_ae,
  input [53:0] io_ptw_resp_bits_pte_ppn,
  input io_ptw_resp_bits_pte_d,
  input io_ptw_resp_bits_pte_a,
  input io_ptw_resp_bits_pte_g,
  input io_ptw_resp_bits_pte_u,
  input io_ptw_resp_bits_pte_x,
  input io_ptw_resp_bits_pte_w,
  input io_ptw_resp_bits_pte_r,
  input io_ptw_resp_bits_pte_v,
  input [1:0] io_ptw_resp_bits_level,
  input io_ptw_resp_bits_homogeneous,
  input [3:0] io_ptw_ptbr_mode,
  input io_ptw_status_debug,
  input [1:0] io_ptw_status_prv,
  input io_ptw_pmp_0_cfg_l,
  input [1:0] io_ptw_pmp_0_cfg_a,
  input io_ptw_pmp_0_cfg_x,
  input io_ptw_pmp_0_cfg_w,
  input io_ptw_pmp_0_cfg_r,
  input [29:0] io_ptw_pmp_0_addr,
  input [31:0] io_ptw_pmp_0_mask,
  input io_ptw_pmp_1_cfg_l,
  input [1:0] io_ptw_pmp_1_cfg_a,
  input io_ptw_pmp_1_cfg_x,
  input io_ptw_pmp_1_cfg_w,
  input io_ptw_pmp_1_cfg_r,
  input [29:0] io_ptw_pmp_1_addr,
  input [31:0] io_ptw_pmp_1_mask,
  input io_ptw_pmp_2_cfg_l,
  input [1:0] io_ptw_pmp_2_cfg_a,
  input io_ptw_pmp_2_cfg_x,
  input io_ptw_pmp_2_cfg_w,
  input io_ptw_pmp_2_cfg_r,
  input [29:0] io_ptw_pmp_2_addr,
  input [31:0] io_ptw_pmp_2_mask,
  input io_ptw_pmp_3_cfg_l,
  input [1:0] io_ptw_pmp_3_cfg_a,
  input io_ptw_pmp_3_cfg_x,
  input io_ptw_pmp_3_cfg_w,
  input io_ptw_pmp_3_cfg_r,
  input [29:0] io_ptw_pmp_3_addr,
  input [31:0] io_ptw_pmp_3_mask,
  input io_ptw_pmp_4_cfg_l,
  input [1:0] io_ptw_pmp_4_cfg_a,
  input io_ptw_pmp_4_cfg_x,
  input io_ptw_pmp_4_cfg_w,
  input io_ptw_pmp_4_cfg_r,
  input [29:0] io_ptw_pmp_4_addr,
  input [31:0] io_ptw_pmp_4_mask,
  input io_ptw_pmp_5_cfg_l,
  input [1:0] io_ptw_pmp_5_cfg_a,
  input io_ptw_pmp_5_cfg_x,
  input io_ptw_pmp_5_cfg_w,
  input io_ptw_pmp_5_cfg_r,
  input [29:0] io_ptw_pmp_5_addr,
  input [31:0] io_ptw_pmp_5_mask,
  input io_ptw_pmp_6_cfg_l,
  input [1:0] io_ptw_pmp_6_cfg_a,
  input io_ptw_pmp_6_cfg_x,
  input io_ptw_pmp_6_cfg_w,
  input io_ptw_pmp_6_cfg_r,
  input [29:0] io_ptw_pmp_6_addr,
  input [31:0] io_ptw_pmp_6_mask,
  input io_ptw_pmp_7_cfg_l,
  input [1:0] io_ptw_pmp_7_cfg_a,
  input io_ptw_pmp_7_cfg_x,
  input io_ptw_pmp_7_cfg_w,
  input io_ptw_pmp_7_cfg_r,
  input [29:0] io_ptw_pmp_7_addr,
  input [31:0] io_ptw_pmp_7_mask,
  input [63:0] io_ptw_customCSRs_csrs_0_value,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input icache_halt,
  input fq_halt,
  input tlb_halt,
  input btb_halt) ; 
   wire icache_clock ;  
   wire icache_reset ;  
   wire icache_auto_master_out_a_ready ;  
   wire icache_auto_master_out_a_valid ;  
   wire [31:0] icache_auto_master_out_a_bits_address ;  
   wire icache_auto_master_out_d_valid ;  
   wire [2:0] icache_auto_master_out_d_bits_opcode ;  
   wire [3:0] icache_auto_master_out_d_bits_size ;  
   wire [63:0] icache_auto_master_out_d_bits_data ;  
   wire icache_auto_master_out_d_bits_corrupt ;  
   wire icache_io_req_ready ;  
   wire icache_io_req_valid ;  
   wire [38:0] icache_io_req_bits_addr ;  
   wire [31:0] icache_io_s1_paddr ;  
   wire icache_io_s1_kill ;  
   wire icache_io_s2_kill ;  
   wire icache_io_resp_valid ;  
   wire [31:0] icache_io_resp_bits_data ;  
   wire icache_io_resp_bits_replay ;  
   wire icache_io_resp_bits_ae ;  
   wire icache_io_invalidate ;  
   wire [29:0] icache_io_covSum ;  
   wire icache_metaAssert ;  
   wire icache_metaReset ;  
   wire icache_repl_way_v0_prng_halt ;  
   wire fq_clock ;  
   wire fq_reset ;  
   wire fq_io_enq_ready ;  
   wire fq_io_enq_valid ;  
   wire fq_io_enq_bits_btb_taken ;  
   wire fq_io_enq_bits_btb_bridx ;  
   wire [4:0] fq_io_enq_bits_btb_entry ;  
   wire [7:0] fq_io_enq_bits_btb_bht_history ;  
   wire [39:0] fq_io_enq_bits_pc ;  
   wire [31:0] fq_io_enq_bits_data ;  
   wire [1:0] fq_io_enq_bits_mask ;  
   wire fq_io_enq_bits_xcpt_pf_inst ;  
   wire fq_io_enq_bits_xcpt_ae_inst ;  
   wire fq_io_enq_bits_replay ;  
   wire fq_io_deq_ready ;  
   wire fq_io_deq_valid ;  
   wire fq_io_deq_bits_btb_taken ;  
   wire fq_io_deq_bits_btb_bridx ;  
   wire [4:0] fq_io_deq_bits_btb_entry ;  
   wire [7:0] fq_io_deq_bits_btb_bht_history ;  
   wire [39:0] fq_io_deq_bits_pc ;  
   wire [31:0] fq_io_deq_bits_data ;  
   wire fq_io_deq_bits_xcpt_pf_inst ;  
   wire fq_io_deq_bits_xcpt_ae_inst ;  
   wire fq_io_deq_bits_replay ;  
   wire [4:0] fq_io_mask ;  
   wire [29:0] fq_io_covSum ;  
   wire fq_metaAssert ;  
   wire fq_metaReset ;  
   wire tlb_clock ;  
   wire tlb_reset ;  
   wire tlb_io_req_ready ;  
   wire tlb_io_req_valid ;  
   wire [39:0] tlb_io_req_bits_vaddr ;  
   wire tlb_io_resp_miss ;  
   wire [31:0] tlb_io_resp_paddr ;  
   wire tlb_io_resp_pf_inst ;  
   wire tlb_io_resp_ae_inst ;  
   wire tlb_io_resp_cacheable ;  
   wire tlb_io_sfence_valid ;  
   wire tlb_io_sfence_bits_rs1 ;  
   wire tlb_io_sfence_bits_rs2 ;  
   wire [38:0] tlb_io_sfence_bits_addr ;  
   wire tlb_io_ptw_req_ready ;  
   wire tlb_io_ptw_req_valid ;  
   wire tlb_io_ptw_req_bits_valid ;  
   wire [26:0] tlb_io_ptw_req_bits_bits_addr ;  
   wire tlb_io_ptw_resp_valid ;  
   wire tlb_io_ptw_resp_bits_ae ;  
   wire [53:0] tlb_io_ptw_resp_bits_pte_ppn ;  
   wire tlb_io_ptw_resp_bits_pte_d ;  
   wire tlb_io_ptw_resp_bits_pte_a ;  
   wire tlb_io_ptw_resp_bits_pte_g ;  
   wire tlb_io_ptw_resp_bits_pte_u ;  
   wire tlb_io_ptw_resp_bits_pte_x ;  
   wire tlb_io_ptw_resp_bits_pte_w ;  
   wire tlb_io_ptw_resp_bits_pte_r ;  
   wire tlb_io_ptw_resp_bits_pte_v ;  
   wire [1:0] tlb_io_ptw_resp_bits_level ;  
   wire tlb_io_ptw_resp_bits_homogeneous ;  
   wire [3:0] tlb_io_ptw_ptbr_mode ;  
   wire tlb_io_ptw_status_debug ;  
   wire [1:0] tlb_io_ptw_status_prv ;  
   wire tlb_io_ptw_pmp_0_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_0_cfg_a ;  
   wire tlb_io_ptw_pmp_0_cfg_x ;  
   wire tlb_io_ptw_pmp_0_cfg_w ;  
   wire tlb_io_ptw_pmp_0_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_0_addr ;  
   wire [31:0] tlb_io_ptw_pmp_0_mask ;  
   wire tlb_io_ptw_pmp_1_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_1_cfg_a ;  
   wire tlb_io_ptw_pmp_1_cfg_x ;  
   wire tlb_io_ptw_pmp_1_cfg_w ;  
   wire tlb_io_ptw_pmp_1_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_1_addr ;  
   wire [31:0] tlb_io_ptw_pmp_1_mask ;  
   wire tlb_io_ptw_pmp_2_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_2_cfg_a ;  
   wire tlb_io_ptw_pmp_2_cfg_x ;  
   wire tlb_io_ptw_pmp_2_cfg_w ;  
   wire tlb_io_ptw_pmp_2_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_2_addr ;  
   wire [31:0] tlb_io_ptw_pmp_2_mask ;  
   wire tlb_io_ptw_pmp_3_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_3_cfg_a ;  
   wire tlb_io_ptw_pmp_3_cfg_x ;  
   wire tlb_io_ptw_pmp_3_cfg_w ;  
   wire tlb_io_ptw_pmp_3_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_3_addr ;  
   wire [31:0] tlb_io_ptw_pmp_3_mask ;  
   wire tlb_io_ptw_pmp_4_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_4_cfg_a ;  
   wire tlb_io_ptw_pmp_4_cfg_x ;  
   wire tlb_io_ptw_pmp_4_cfg_w ;  
   wire tlb_io_ptw_pmp_4_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_4_addr ;  
   wire [31:0] tlb_io_ptw_pmp_4_mask ;  
   wire tlb_io_ptw_pmp_5_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_5_cfg_a ;  
   wire tlb_io_ptw_pmp_5_cfg_x ;  
   wire tlb_io_ptw_pmp_5_cfg_w ;  
   wire tlb_io_ptw_pmp_5_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_5_addr ;  
   wire [31:0] tlb_io_ptw_pmp_5_mask ;  
   wire tlb_io_ptw_pmp_6_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_6_cfg_a ;  
   wire tlb_io_ptw_pmp_6_cfg_x ;  
   wire tlb_io_ptw_pmp_6_cfg_w ;  
   wire tlb_io_ptw_pmp_6_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_6_addr ;  
   wire [31:0] tlb_io_ptw_pmp_6_mask ;  
   wire tlb_io_ptw_pmp_7_cfg_l ;  
   wire [1:0] tlb_io_ptw_pmp_7_cfg_a ;  
   wire tlb_io_ptw_pmp_7_cfg_x ;  
   wire tlb_io_ptw_pmp_7_cfg_w ;  
   wire tlb_io_ptw_pmp_7_cfg_r ;  
   wire [29:0] tlb_io_ptw_pmp_7_addr ;  
   wire [31:0] tlb_io_ptw_pmp_7_mask ;  
   wire tlb_io_kill ;  
   wire [29:0] tlb_io_covSum ;  
   wire tlb_metaAssert ;  
   wire tlb_metaReset ;  
   wire btb_clock ;  
   wire btb_reset ;  
   wire [38:0] btb_io_req_bits_addr ;  
   wire btb_io_resp_valid ;  
   wire btb_io_resp_bits_taken ;  
   wire btb_io_resp_bits_bridx ;  
   wire [38:0] btb_io_resp_bits_target ;  
   wire [4:0] btb_io_resp_bits_entry ;  
   wire [7:0] btb_io_resp_bits_bht_history ;  
   wire btb_io_resp_bits_bht_value ;  
   wire btb_io_btb_update_valid ;  
   wire [4:0] btb_io_btb_update_bits_prediction_entry ;  
   wire [38:0] btb_io_btb_update_bits_pc ;  
   wire btb_io_btb_update_bits_isValid ;  
   wire [38:0] btb_io_btb_update_bits_br_pc ;  
   wire [1:0] btb_io_btb_update_bits_cfiType ;  
   wire btb_io_bht_update_valid ;  
   wire [7:0] btb_io_bht_update_bits_prediction_history ;  
   wire [38:0] btb_io_bht_update_bits_pc ;  
   wire btb_io_bht_update_bits_branch ;  
   wire btb_io_bht_update_bits_taken ;  
   wire btb_io_bht_update_bits_mispredict ;  
   wire btb_io_bht_advance_valid ;  
   wire btb_io_bht_advance_bits_bht_value ;  
   wire btb_io_ras_update_valid ;  
   wire [1:0] btb_io_ras_update_bits_cfiType ;  
   wire [38:0] btb_io_ras_update_bits_returnAddr ;  
   wire btb_io_ras_head_valid ;  
   wire [38:0] btb_io_ras_head_bits ;  
   wire btb_io_flush ;  
   wire [29:0] btb_io_covSum ;  
   wire btb_metaAssert ;  
   wire btb_metaReset ;  
   wire _T_2 ;  
   wire _T_3 ;  
   wire _T_4 ;  
   wire _T_5 ;  
   wire _T_7 ;  
   wire _T_9 ;  
   reg s1_valid ;  
   reg [31:0] _RAND_0 ;  
   reg s2_valid ;  
   reg [31:0] _RAND_1 ;  
   wire _s0_fq_has_space_T_6 ;  
   wire _s0_fq_has_space_T_7 ;  
   wire _s0_fq_has_space_T_8 ;  
   wire _s0_fq_has_space_T_13 ;  
   wire _s0_fq_has_space_T_14 ;  
   wire s0_fq_has_space ;  
   wire s0_valid ;  
   reg [39:0] s1_pc ;  
   reg [63:0] _RAND_2 ;  
   reg s1_speculative ;  
   reg [31:0] _RAND_3 ;  
   wire [31:0] _s2_pc_T_1 ;  
   reg [39:0] s2_pc ;  
   reg [63:0] _RAND_4 ;  
   reg s2_btb_resp_valid ;  
   reg [31:0] _RAND_5 ;  
   reg s2_btb_resp_bits_taken ;  
   reg [31:0] _RAND_6 ;  
   reg s2_btb_resp_bits_bridx ;  
   reg [31:0] _RAND_7 ;  
   reg [4:0] s2_btb_resp_bits_entry ;  
   reg [31:0] _RAND_8 ;  
   reg [7:0] s2_btb_resp_bits_bht_history ;  
   reg [31:0] _RAND_9 ;  
   reg s2_btb_resp_bits_bht_value ;  
   reg [31:0] _RAND_10 ;  
   wire s2_btb_taken ;  
   reg s2_tlb_resp_miss ;  
   reg [31:0] _RAND_11 ;  
   reg s2_tlb_resp_pf_inst ;  
   reg [31:0] _RAND_12 ;  
   reg s2_tlb_resp_ae_inst ;  
   reg [31:0] _RAND_13 ;  
   reg s2_tlb_resp_cacheable ;  
   reg [31:0] _RAND_14 ;  
   wire s2_xcpt ;  
   reg s2_speculative ;  
   reg [31:0] _RAND_15 ;  
   reg s2_partial_insn_valid ;  
   reg [31:0] _RAND_16 ;  
   reg [15:0] s2_partial_insn ;  
   reg [31:0] _RAND_17 ;  
   reg wrong_path ;  
   reg [31:0] _RAND_18 ;  
   wire [39:0] _s1_base_pc_T_1 ;  
   wire [39:0] s1_base_pc ;  
   wire [39:0] ntpc ;  
   wire _s2_replay_T ;  
   wire _s2_replay_T_2 ;  
   reg s2_replay_REG ;  
   reg [31:0] _RAND_19 ;  
   wire s2_replay ;  
   wire _s2_replay_T_4 ;  
   wire _taken_prevRVI_T_1 ;  
   wire taken_prevRVI ;  
   wire [15:0] taken_bits ;  
   wire [31:0] taken_rviBits ;  
   wire taken_rviJump ;  
   wire taken_rviJALR ;  
   wire _taken_taken_T ;  
   wire taken_rviBranch ;  
   wire _taken_taken_T_1 ;  
   wire _taken_taken_T_2 ;  
   wire _taken_taken_T_3 ;  
   wire taken_valid ;  
   wire [15:0] _taken_rvcJump_T ;  
   wire taken_rvcJump ;  
   wire [15:0] _taken_rvcJALR_T ;  
   wire _taken_rvcJALR_T_1 ;  
   wire _taken_rvcJALR_T_3 ;  
   wire taken_rvcJALR ;  
   wire _taken_taken_T_4 ;  
   wire _taken_rvcJR_T_1 ;  
   wire taken_rvcJR ;  
   wire _taken_taken_T_5 ;  
   wire _taken_rvcBranch_T_1 ;  
   wire _taken_rvcBranch_T_3 ;  
   wire taken_rvcBranch ;  
   wire _taken_taken_T_6 ;  
   wire _taken_taken_T_7 ;  
   wire _taken_taken_T_8 ;  
   wire taken_taken ;  
   wire taken_idx ;  
   wire _taken_prevRVI_T_4 ;  
   wire taken_prevRVI_1 ;  
   wire [15:0] taken_bits_1 ;  
   wire [31:0] taken_rviBits_1 ;  
   wire taken_rviJALR_1 ;  
   wire _taken_rviReturn_T_8 ;  
   wire [4:0] _taken_rviReturn_T_10 ;  
   wire _taken_rviReturn_T_11 ;  
   wire taken_rviReturn_1 ;  
   wire _taken_predictReturn_T_3 ;  
   wire taken_valid_1 ;  
   wire [15:0] _taken_rvcJR_T_4 ;  
   wire _taken_rvcJR_T_5 ;  
   wire _taken_rvcJR_T_7 ;  
   wire taken_rvcJR_1 ;  
   wire [4:0] _taken_rvcReturn_T_4 ;  
   wire _taken_rvcReturn_T_5 ;  
   wire taken_rvcReturn_1 ;  
   wire _taken_predictReturn_T_4 ;  
   wire _taken_predictReturn_T_5 ;  
   wire taken_predictReturn_1 ;  
   wire _taken_T_45 ;  
   wire _taken_rviReturn_T_2 ;  
   wire [4:0] _taken_rviReturn_T_4 ;  
   wire _taken_rviReturn_T_5 ;  
   wire taken_rviReturn ;  
   wire _taken_predictReturn_T ;  
   wire [4:0] _taken_rvcReturn_T_1 ;  
   wire _taken_rvcReturn_T_2 ;  
   wire taken_rvcReturn ;  
   wire _taken_predictReturn_T_1 ;  
   wire _taken_predictReturn_T_2 ;  
   wire taken_predictReturn ;  
   wire _taken_T_16 ;  
   wire _GEN_45 ;  
   wire _GEN_78 ;  
   wire _GEN_81 ;  
   wire useRAS ;  
   wire taken_rviBranch_1 ;  
   wire _taken_predictBranch_T_3 ;  
   wire [15:0] _taken_rvcBranch_T_4 ;  
   wire _taken_rvcBranch_T_5 ;  
   wire _taken_rvcBranch_T_7 ;  
   wire taken_rvcBranch_1 ;  
   wire _taken_predictBranch_T_4 ;  
   wire _taken_predictBranch_T_5 ;  
   wire taken_predictBranch_1 ;  
   wire taken_rviJump_1 ;  
   wire _taken_predictJump_T_2 ;  
   wire taken_rvcJump_1 ;  
   wire _taken_predictJump_T_3 ;  
   wire taken_predictJump_1 ;  
   wire _taken_T_46 ;  
   wire _taken_T_47 ;  
   wire [39:0] _s2_base_pc_T_1 ;  
   wire [39:0] s2_base_pc ;  
   wire [39:0] taken_pc_1 ;  
   wire [39:0] _taken_npc_T_6 ;  
   wire [39:0] _taken_npc_T_8 ;  
   wire taken_rviImm_sign_2 ;  
   wire taken_rviImm_hi_hi_hi_2 ;  
   wire [10:0] taken_rviImm_hi_hi_lo_2 ;  
   wire [7:0] taken_rviImm_hi_lo_hi_2 ;  
   wire taken_rviImm_hi_lo_lo_2 ;  
   wire [5:0] taken_rviImm_lo_hi_hi_2 ;  
   wire [3:0] taken_rviImm_lo_hi_lo_2 ;  
   wire [31:0] _taken_rviImm_T_7 ;  
   wire [7:0] taken_rviImm_hi_lo_hi_3 ;  
   wire taken_rviImm_hi_lo_lo_3 ;  
   wire [31:0] _taken_rviImm_T_9 ;  
   wire [31:0] taken_rviImm_1 ;  
   wire [4:0] taken_rvcImm_hi_hi_hi_2 ;  
   wire [1:0] taken_rvcImm_hi_hi_lo_2 ;  
   wire taken_rvcImm_hi_lo_2 ;  
   wire [1:0] taken_rvcImm_lo_hi_hi_2 ;  
   wire [1:0] taken_rvcImm_lo_hi_lo_2 ;  
   wire [12:0] _taken_rvcImm_T_13 ;  
   wire [9:0] taken_rvcImm_hi_hi_hi_hi_1 ;  
   wire taken_rvcImm_hi_hi_hi_lo_1 ;  
   wire [1:0] taken_rvcImm_hi_hi_lo_3 ;  
   wire taken_rvcImm_hi_lo_hi_1 ;  
   wire taken_rvcImm_hi_lo_lo_1 ;  
   wire taken_rvcImm_lo_hi_lo_3 ;  
   wire [2:0] taken_rvcImm_lo_lo_hi_1 ;  
   wire [20:0] _taken_rvcImm_T_17 ;  
   wire [20:0] taken_rvcImm_1 ;  
   wire [31:0] _taken_npc_T_9 ;  
   wire [39:0] _GEN_127 ;  
   wire [39:0] _taken_predicted_npc_T_1 ;  
   wire _taken_predictBranch_T ;  
   wire _taken_predictBranch_T_1 ;  
   wire _taken_predictBranch_T_2 ;  
   wire taken_predictBranch ;  
   wire _taken_predictJump_T ;  
   wire _taken_predictJump_T_1 ;  
   wire taken_predictJump ;  
   wire _taken_T_17 ;  
   wire _taken_T_18 ;  
   wire [39:0] _taken_npc_T ;  
   wire taken_rviImm_sign ;  
   wire taken_rviImm_hi_hi_hi ;  
   wire [10:0] taken_rviImm_hi_hi_lo ;  
   wire [7:0] taken_rviImm_hi_lo_hi ;  
   wire taken_rviImm_hi_lo_lo ;  
   wire [5:0] taken_rviImm_lo_hi_hi ;  
   wire [3:0] taken_rviImm_lo_hi_lo ;  
   wire [31:0] _taken_rviImm_T_2 ;  
   wire [7:0] taken_rviImm_hi_lo_hi_1 ;  
   wire taken_rviImm_hi_lo_lo_1 ;  
   wire [31:0] _taken_rviImm_T_4 ;  
   wire [31:0] taken_rviImm ;  
   wire [32:0] _taken_npc_T_1 ;  
   wire [4:0] taken_rvcImm_hi_hi_hi ;  
   wire [1:0] taken_rvcImm_hi_hi_lo ;  
   wire taken_rvcImm_hi_lo ;  
   wire [1:0] taken_rvcImm_lo_hi_hi ;  
   wire [1:0] taken_rvcImm_lo_hi_lo ;  
   wire [12:0] _taken_rvcImm_T_4 ;  
   wire [9:0] taken_rvcImm_hi_hi_hi_hi ;  
   wire taken_rvcImm_hi_hi_hi_lo ;  
   wire [1:0] taken_rvcImm_hi_hi_lo_1 ;  
   wire taken_rvcImm_hi_lo_hi ;  
   wire taken_rvcImm_hi_lo_lo ;  
   wire taken_rvcImm_lo_hi_lo_1 ;  
   wire [2:0] taken_rvcImm_lo_lo_hi ;  
   wire [20:0] _taken_rvcImm_T_8 ;  
   wire [20:0] taken_rvcImm ;  
   wire [32:0] _taken_npc_T_2 ;  
   wire [39:0] _GEN_128 ;  
   wire [39:0] _taken_predicted_npc_T ;  
   wire predicted_taken ;  
   wire predicted_npc_hi ;  
   wire [39:0] _predicted_npc_T ;  
   wire [39:0] _GEN_28 ;  
   wire [39:0] _GEN_43 ;  
   wire [39:0] _GEN_46 ;  
   wire [39:0] _GEN_79 ;  
   wire [39:0] _GEN_82 ;  
   wire [39:0] _GEN_99 ;  
   wire [39:0] predicted_npc ;  
   wire [39:0] npc ;  
   wire _s0_speculative_T_1 ;  
   wire _s0_speculative_T_2 ;  
   wire s0_speculative ;  
   wire _taken_taken_T_9 ;  
   wire _taken_taken_T_10 ;  
   wire _taken_taken_T_11 ;  
   wire _taken_taken_T_12 ;  
   wire _taken_rvcJALR_T_5 ;  
   wire taken_rvcJALR_1 ;  
   wire _taken_taken_T_13 ;  
   wire _taken_taken_T_14 ;  
   wire _taken_taken_T_15 ;  
   wire _taken_taken_T_16 ;  
   wire _taken_taken_T_17 ;  
   wire taken_taken_1 ;  
   wire taken ;  
   wire _GEN_116 ;  
   wire _GEN_120 ;  
   wire s2_redirect ;  
   wire _GEN_0 ;  
   wire _icache_io_s1_kill_T ;  
   wire s2_can_speculatively_refill ;  
   wire _icache_io_s2_kill_T_1 ;  
   reg fq_io_enq_valid_REG ;  
   reg [31:0] _RAND_20 ;  
   wire _fq_io_enq_valid_T ;  
   wire _fq_io_enq_valid_T_2 ;  
   wire _fq_io_enq_valid_T_3 ;  
   wire [39:0] _io_cpu_npc_T ;  
   wire [39:0] _io_cpu_npc_T_2 ;  
   wire [2:0] _fq_io_enq_bits_mask_T_1 ;  
   wire _fq_io_enq_bits_replay_T_1 ;  
   wire _fq_io_enq_bits_replay_T_3 ;  
   wire _fq_io_enq_bits_replay_T_4 ;  
   wire _T_13 ;  
   wire _T_15 ;  
   wire _T_18 ;  
   wire _T_20 ;  
   wire fetch_bubble_likely ;  
   wire _btb_io_btb_update_valid_T_2 ;  
   wire _btb_io_btb_update_valid_T_3 ;  
   wire _taken_T_53 ;  
   wire _taken_T_54 ;  
   wire _taken_T_55 ;  
   wire _taken_T_56 ;  
   wire _taken_T_24 ;  
   wire _taken_T_25 ;  
   wire _taken_T_26 ;  
   wire _taken_T_27 ;  
   wire _GEN_92 ;  
   wire updateBTB ;  
   wire _btb_io_btb_update_valid_T_4 ;  
   wire [1:0] _btb_io_btb_update_bits_br_pc_T ;  
   wire [39:0] _GEN_129 ;  
   wire [39:0] _btb_io_btb_update_bits_br_pc_T_1 ;  
   wire [39:0] _GEN_36 ;  
   wire [39:0] _GEN_37 ;  
   wire [1:0] after_idx ;  
   wire [2:0] _btb_io_ras_update_bits_returnAddr_T ;  
   wire [39:0] _GEN_130 ;  
   wire [39:0] _btb_io_ras_update_bits_returnAddr_T_2 ;  
   wire _taken_rviCall_T ;  
   wire taken_rviCall ;  
   wire _taken_T ;  
   wire _taken_T_2 ;  
   wire _taken_T_3 ;  
   wire _taken_T_5 ;  
   wire _GEN_39 ;  
   wire _GEN_40 ;  
   wire _taken_btb_io_ras_update_valid_T_3 ;  
   wire _taken_btb_io_ras_update_valid_T_4 ;  
   wire _taken_btb_io_ras_update_valid_T_5 ;  
   wire _taken_btb_io_ras_update_valid_T_6 ;  
   wire _taken_btb_io_ras_update_valid_T_7 ;  
   wire _taken_btb_io_ras_update_valid_T_8 ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T_1 ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T_2 ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T_5 ;  
   wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_6 ;  
   wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_7 ;  
   wire _taken_T_9 ;  
   wire _taken_T_11 ;  
   wire _taken_T_13 ;  
   wire _taken_T_15 ;  
   wire _GEN_41 ;  
   wire _GEN_44 ;  
   wire _GEN_47 ;  
   wire taken_rvc_1 ;  
   wire _taken_rviCall_T_2 ;  
   wire taken_rviCall_1 ;  
   wire _taken_T_31 ;  
   wire _taken_T_32 ;  
   wire _taken_T_34 ;  
   wire _GEN_76 ;  
   wire _taken_btb_io_ras_update_valid_T_12 ;  
   wire _taken_btb_io_ras_update_valid_T_13 ;  
   wire _taken_btb_io_ras_update_valid_T_14 ;  
   wire _taken_btb_io_ras_update_valid_T_15 ;  
   wire _taken_btb_io_ras_update_valid_T_16 ;  
   wire _taken_btb_io_ras_update_valid_T_17 ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T_8 ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T_9 ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T_10 ;  
   wire _taken_btb_io_ras_update_bits_cfiType_T_13 ;  
   wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_14 ;  
   wire [1:0] _taken_btb_io_ras_update_bits_cfiType_T_15 ;  
   wire _taken_T_38 ;  
   wire _taken_T_40 ;  
   wire _taken_T_42 ;  
   wire _taken_T_44 ;  
   wire _GEN_77 ;  
   wire _GEN_83 ;  
   wire _taken_T_59 ;  
   wire _taken_T_61 ;  
   wire [15:0] _taken_lo_T ;  
   wire _T_25 ;  
   wire _T_26 ;  
   wire _GEN_117 ;  
   wire _GEN_118 ;  
   wire [4:0] _GEN_119 ;  
   wire _T_31 ;  
   wire _T_33 ;  
   reg [5:0] Frontend_state ;  
   reg [31:0] _RAND_21 ;  
   reg Frontend_cov[0:63] ;  
   reg [31:0] _RAND_22 ;  
   wire Frontend_cov_read_data ;  
   wire [5:0] Frontend_cov_read_addr ;  
   wire Frontend_cov_write_data ;  
   wire [5:0] Frontend_cov_write_addr ;  
   wire Frontend_cov_write_mask ;  
   wire Frontend_cov_write_en ;  
   reg [29:0] Frontend_covSum ;  
   reg [31:0] _RAND_23 ;  
   wire s2_partial_insn_valid_shl ;  
   wire [5:0] s2_partial_insn_valid_pad ;  
   wire [1:0] s2_btb_resp_valid_shl ;  
   wire [5:0] s2_btb_resp_valid_pad ;  
   wire [2:0] s2_replay_REG_shl ;  
   wire [5:0] s2_replay_REG_pad ;  
   wire [3:0] s2_btb_resp_bits_bht_value_shl ;  
   wire [5:0] s2_btb_resp_bits_bht_value_pad ;  
   wire [4:0] s2_valid_shl ;  
   wire [5:0] s2_valid_pad ;  
   wire [5:0] s2_btb_resp_bits_taken_shl ;  
   wire [5:0] s2_btb_resp_bits_taken_pad ;  
   wire [5:0] Frontend_xor4 ;  
   wire [5:0] Frontend_xor1 ;  
   wire [5:0] Frontend_xor6 ;  
   wire [5:0] Frontend_xor2 ;  
   wire [5:0] Frontend_xor0 ;  
   wire [29:0] icache_sum ;  
   wire [29:0] fq_sum ;  
   wire [29:0] tlb_sum ;  
   wire [29:0] btb_sum ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire stopEn2 ;  
   wire icache_metaAssert_wire ;  
   wire fq_metaAssert_wire ;  
   wire tlb_metaAssert_wire ;  
   wire btb_metaAssert_wire ;  
   wire Frontend_or4 ;  
   wire Frontend_or1 ;  
   wire Frontend_or5 ;  
   wire Frontend_or6 ;  
   wire Frontend_or2 ;  
   wire Frontend_or0 ;  
  ICache icache(.clock(icache_clock),.reset(icache_reset),.auto_master_out_a_ready(icache_auto_master_out_a_ready),.auto_master_out_a_valid(icache_auto_master_out_a_valid),.auto_master_out_a_bits_address(icache_auto_master_out_a_bits_address),.auto_master_out_d_valid(icache_auto_master_out_d_valid),.auto_master_out_d_bits_opcode(icache_auto_master_out_d_bits_opcode),.auto_master_out_d_bits_size(icache_auto_master_out_d_bits_size),.auto_master_out_d_bits_data(icache_auto_master_out_d_bits_data),.auto_master_out_d_bits_corrupt(icache_auto_master_out_d_bits_corrupt),.io_req_ready(icache_io_req_ready),.io_req_valid(icache_io_req_valid),.io_req_bits_addr(icache_io_req_bits_addr),.io_s1_paddr(icache_io_s1_paddr),.io_s1_kill(icache_io_s1_kill),.io_s2_kill(icache_io_s2_kill),.io_resp_valid(icache_io_resp_valid),.io_resp_bits_data(icache_io_resp_bits_data),.io_resp_bits_replay(icache_io_resp_bits_replay),.io_resp_bits_ae(icache_io_resp_bits_ae),.io_invalidate(icache_io_invalidate),.io_covSum(icache_io_covSum),.metaAssert(icache_metaAssert),.metaReset(icache_metaReset),.repl_way_v0_prng_halt(icache_repl_way_v0_prng_halt)); 
  ShiftQueue fq(.clock(fq_clock),.reset(fq_reset),.io_enq_ready(fq_io_enq_ready),.io_enq_valid(fq_io_enq_valid),.io_enq_bits_btb_taken(fq_io_enq_bits_btb_taken),.io_enq_bits_btb_bridx(fq_io_enq_bits_btb_bridx),.io_enq_bits_btb_entry(fq_io_enq_bits_btb_entry),.io_enq_bits_btb_bht_history(fq_io_enq_bits_btb_bht_history),.io_enq_bits_pc(fq_io_enq_bits_pc),.io_enq_bits_data(fq_io_enq_bits_data),.io_enq_bits_mask(fq_io_enq_bits_mask),.io_enq_bits_xcpt_pf_inst(fq_io_enq_bits_xcpt_pf_inst),.io_enq_bits_xcpt_ae_inst(fq_io_enq_bits_xcpt_ae_inst),.io_enq_bits_replay(fq_io_enq_bits_replay),.io_deq_ready(fq_io_deq_ready),.io_deq_valid(fq_io_deq_valid),.io_deq_bits_btb_taken(fq_io_deq_bits_btb_taken),.io_deq_bits_btb_bridx(fq_io_deq_bits_btb_bridx),.io_deq_bits_btb_entry(fq_io_deq_bits_btb_entry),.io_deq_bits_btb_bht_history(fq_io_deq_bits_btb_bht_history),.io_deq_bits_pc(fq_io_deq_bits_pc),.io_deq_bits_data(fq_io_deq_bits_data),.io_deq_bits_xcpt_pf_inst(fq_io_deq_bits_xcpt_pf_inst),.io_deq_bits_xcpt_ae_inst(fq_io_deq_bits_xcpt_ae_inst),.io_deq_bits_replay(fq_io_deq_bits_replay),.io_mask(fq_io_mask),.io_covSum(fq_io_covSum),.metaAssert(fq_metaAssert),.metaReset(fq_metaReset)); 
  TLB_1 tlb(.clock(tlb_clock),.reset(tlb_reset),.io_req_ready(tlb_io_req_ready),.io_req_valid(tlb_io_req_valid),.io_req_bits_vaddr(tlb_io_req_bits_vaddr),.io_resp_miss(tlb_io_resp_miss),.io_resp_paddr(tlb_io_resp_paddr),.io_resp_pf_inst(tlb_io_resp_pf_inst),.io_resp_ae_inst(tlb_io_resp_ae_inst),.io_resp_cacheable(tlb_io_resp_cacheable),.io_sfence_valid(tlb_io_sfence_valid),.io_sfence_bits_rs1(tlb_io_sfence_bits_rs1),.io_sfence_bits_rs2(tlb_io_sfence_bits_rs2),.io_sfence_bits_addr(tlb_io_sfence_bits_addr),.io_ptw_req_ready(tlb_io_ptw_req_ready),.io_ptw_req_valid(tlb_io_ptw_req_valid),.io_ptw_req_bits_valid(tlb_io_ptw_req_bits_valid),.io_ptw_req_bits_bits_addr(tlb_io_ptw_req_bits_bits_addr),.io_ptw_resp_valid(tlb_io_ptw_resp_valid),.io_ptw_resp_bits_ae(tlb_io_ptw_resp_bits_ae),.io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),.io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),.io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),.io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),.io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),.io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),.io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),.io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),.io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),.io_ptw_resp_bits_level(tlb_io_ptw_resp_bits_level),.io_ptw_resp_bits_homogeneous(tlb_io_ptw_resp_bits_homogeneous),.io_ptw_ptbr_mode(tlb_io_ptw_ptbr_mode),.io_ptw_status_debug(tlb_io_ptw_status_debug),.io_ptw_status_prv(tlb_io_ptw_status_prv),.io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),.io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),.io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),.io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),.io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),.io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),.io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),.io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),.io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),.io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),.io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),.io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),.io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),.io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),.io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),.io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),.io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),.io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),.io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),.io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),.io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),.io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),.io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),.io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),.io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),.io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),.io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),.io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),.io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),.io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),.io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),.io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),.io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),.io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),.io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),.io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),.io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),.io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),.io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),.io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),.io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),.io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),.io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),.io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),.io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),.io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),.io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),.io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),.io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),.io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),.io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),.io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),.io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),.io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),.io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),.io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask),.io_kill(tlb_io_kill),.io_covSum(tlb_io_covSum),.metaAssert(tlb_metaAssert),.metaReset(tlb_metaReset)); 
  BTB btb(.clock(btb_clock),.reset(btb_reset),.io_req_bits_addr(btb_io_req_bits_addr),.io_resp_valid(btb_io_resp_valid),.io_resp_bits_taken(btb_io_resp_bits_taken),.io_resp_bits_bridx(btb_io_resp_bits_bridx),.io_resp_bits_target(btb_io_resp_bits_target),.io_resp_bits_entry(btb_io_resp_bits_entry),.io_resp_bits_bht_history(btb_io_resp_bits_bht_history),.io_resp_bits_bht_value(btb_io_resp_bits_bht_value),.io_btb_update_valid(btb_io_btb_update_valid),.io_btb_update_bits_prediction_entry(btb_io_btb_update_bits_prediction_entry),.io_btb_update_bits_pc(btb_io_btb_update_bits_pc),.io_btb_update_bits_isValid(btb_io_btb_update_bits_isValid),.io_btb_update_bits_br_pc(btb_io_btb_update_bits_br_pc),.io_btb_update_bits_cfiType(btb_io_btb_update_bits_cfiType),.io_bht_update_valid(btb_io_bht_update_valid),.io_bht_update_bits_prediction_history(btb_io_bht_update_bits_prediction_history),.io_bht_update_bits_pc(btb_io_bht_update_bits_pc),.io_bht_update_bits_branch(btb_io_bht_update_bits_branch),.io_bht_update_bits_taken(btb_io_bht_update_bits_taken),.io_bht_update_bits_mispredict(btb_io_bht_update_bits_mispredict),.io_bht_advance_valid(btb_io_bht_advance_valid),.io_bht_advance_bits_bht_value(btb_io_bht_advance_bits_bht_value),.io_ras_update_valid(btb_io_ras_update_valid),.io_ras_update_bits_cfiType(btb_io_ras_update_bits_cfiType),.io_ras_update_bits_returnAddr(btb_io_ras_update_bits_returnAddr),.io_ras_head_valid(btb_io_ras_head_valid),.io_ras_head_bits(btb_io_ras_head_bits),.io_flush(btb_io_flush),.io_covSum(btb_io_covSum),.metaAssert(btb_metaAssert),.metaReset(btb_metaReset)); 
  assign _T_2=io_cpu_req_valid|io_cpu_sfence_valid; 
  assign _T_3=_T_2|io_cpu_flush_icache; 
  assign _T_4=_T_3|io_cpu_bht_update_valid; 
  assign _T_5=_T_4|io_cpu_btb_update_valid; 
  assign _T_7=~_T_5|io_cpu_might_request; 
  assign _T_9=_T_7|reset; 
  assign _s0_fq_has_space_T_6=~s1_valid|~s2_valid; 
  assign _s0_fq_has_space_T_7=~fq_io_mask[3]&_s0_fq_has_space_T_6; 
  assign _s0_fq_has_space_T_8=~fq_io_mask[2]|_s0_fq_has_space_T_7; 
  assign _s0_fq_has_space_T_13=~s1_valid&~s2_valid; 
  assign _s0_fq_has_space_T_14=~fq_io_mask[4]&_s0_fq_has_space_T_13; 
  assign s0_fq_has_space=_s0_fq_has_space_T_8|_s0_fq_has_space_T_14; 
  assign s0_valid=io_cpu_req_valid|s0_fq_has_space; 
  assign _s2_pc_T_1=~auto_reset_vector_sink_in|32'h1; 
  assign s2_btb_taken=s2_btb_resp_valid&s2_btb_resp_bits_taken; 
  assign s2_xcpt=s2_tlb_resp_ae_inst|s2_tlb_resp_pf_inst; 
  assign _s1_base_pc_T_1=~s1_pc|40'h3; 
  assign s1_base_pc=~_s1_base_pc_T_1; 
  assign ntpc=s1_base_pc+40'h4; 
  assign _s2_replay_T=fq_io_enq_ready&fq_io_enq_valid; 
  assign _s2_replay_T_2=s2_valid&~_s2_replay_T; 
  assign s2_replay=_s2_replay_T_2|s2_replay_REG; 
  assign _s2_replay_T_4=s2_replay&~s0_valid; 
  assign _taken_prevRVI_T_1=s2_partial_insn[1:0]!=2'h3; 
  assign taken_prevRVI=s2_partial_insn_valid&~_taken_prevRVI_T_1; 
  assign taken_bits=fq_io_enq_bits_data[15:0]; 
  assign taken_rviBits={taken_bits,s2_partial_insn}; 
  assign taken_rviJump=taken_rviBits[6:0]==7'h6f; 
  assign taken_rviJALR=taken_rviBits[6:0]==7'h67; 
  assign _taken_taken_T=taken_rviJump|taken_rviJALR; 
  assign taken_rviBranch=taken_rviBits[6:0]==7'h63; 
  assign _taken_taken_T_1=taken_rviBranch&s2_btb_resp_bits_bht_value; 
  assign _taken_taken_T_2=_taken_taken_T|_taken_taken_T_1; 
  assign _taken_taken_T_3=taken_prevRVI&_taken_taken_T_2; 
  assign taken_valid=fq_io_enq_bits_mask[0]&~taken_prevRVI; 
  assign _taken_rvcJump_T=taken_bits&16'he003; 
  assign taken_rvcJump=16'ha001==_taken_rvcJump_T; 
  assign _taken_rvcJALR_T=taken_bits&16'hf003; 
  assign _taken_rvcJALR_T_1=16'h9002==_taken_rvcJALR_T; 
  assign _taken_rvcJALR_T_3=taken_bits[6:2]==5'h0; 
  assign taken_rvcJALR=_taken_rvcJALR_T_1&_taken_rvcJALR_T_3; 
  assign _taken_taken_T_4=taken_rvcJump|taken_rvcJALR; 
  assign _taken_rvcJR_T_1=16'h8002==_taken_rvcJALR_T; 
  assign taken_rvcJR=_taken_rvcJR_T_1&_taken_rvcJALR_T_3; 
  assign _taken_taken_T_5=_taken_taken_T_4|taken_rvcJR; 
  assign _taken_rvcBranch_T_1=16'hc001==_taken_rvcJump_T; 
  assign _taken_rvcBranch_T_3=16'he001==_taken_rvcJump_T; 
  assign taken_rvcBranch=_taken_rvcBranch_T_1|_taken_rvcBranch_T_3; 
  assign _taken_taken_T_6=taken_rvcBranch&s2_btb_resp_bits_bht_value; 
  assign _taken_taken_T_7=_taken_taken_T_5|_taken_taken_T_6; 
  assign _taken_taken_T_8=taken_valid&_taken_taken_T_7; 
  assign taken_taken=_taken_taken_T_3|_taken_taken_T_8; 
  assign taken_idx=~taken_taken; 
  assign _taken_prevRVI_T_4=taken_bits[1:0]!=2'h3; 
  assign taken_prevRVI_1=taken_valid&~_taken_prevRVI_T_4; 
  assign taken_bits_1=fq_io_enq_bits_data[31:16]; 
  assign taken_rviBits_1={taken_bits_1,taken_bits}; 
  assign taken_rviJALR_1=taken_rviBits_1[6:0]==7'h67; 
  assign _taken_rviReturn_T_8=taken_rviJALR_1&~taken_rviBits_1[7]; 
  assign _taken_rviReturn_T_10=taken_rviBits_1[19:15]&5'h1b; 
  assign _taken_rviReturn_T_11=5'h1==_taken_rviReturn_T_10; 
  assign taken_rviReturn_1=_taken_rviReturn_T_8&_taken_rviReturn_T_11; 
  assign _taken_predictReturn_T_3=taken_prevRVI_1&taken_rviReturn_1; 
  assign taken_valid_1=fq_io_enq_bits_mask[1]&~taken_prevRVI_1; 
  assign _taken_rvcJR_T_4=taken_bits_1&16'hf003; 
  assign _taken_rvcJR_T_5=16'h8002==_taken_rvcJR_T_4; 
  assign _taken_rvcJR_T_7=taken_bits_1[6:2]==5'h0; 
  assign taken_rvcJR_1=_taken_rvcJR_T_5&_taken_rvcJR_T_7; 
  assign _taken_rvcReturn_T_4=taken_bits_1[11:7]&5'h1b; 
  assign _taken_rvcReturn_T_5=5'h1==_taken_rvcReturn_T_4; 
  assign taken_rvcReturn_1=taken_rvcJR_1&_taken_rvcReturn_T_5; 
  assign _taken_predictReturn_T_4=taken_valid_1&taken_rvcReturn_1; 
  assign _taken_predictReturn_T_5=_taken_predictReturn_T_3|_taken_predictReturn_T_4; 
  assign taken_predictReturn_1=btb_io_ras_head_valid&_taken_predictReturn_T_5; 
  assign _taken_T_45=s2_valid&taken_predictReturn_1; 
  assign _taken_rviReturn_T_2=taken_rviJALR&~taken_rviBits[7]; 
  assign _taken_rviReturn_T_4=taken_rviBits[19:15]&5'h1b; 
  assign _taken_rviReturn_T_5=5'h1==_taken_rviReturn_T_4; 
  assign taken_rviReturn=_taken_rviReturn_T_2&_taken_rviReturn_T_5; 
  assign _taken_predictReturn_T=taken_prevRVI&taken_rviReturn; 
  assign _taken_rvcReturn_T_1=taken_bits[11:7]&5'h1b; 
  assign _taken_rvcReturn_T_2=5'h1==_taken_rvcReturn_T_1; 
  assign taken_rvcReturn=taken_rvcJR&_taken_rvcReturn_T_2; 
  assign _taken_predictReturn_T_1=taken_valid&taken_rvcReturn; 
  assign _taken_predictReturn_T_2=_taken_predictReturn_T|_taken_predictReturn_T_1; 
  assign taken_predictReturn=btb_io_ras_head_valid&_taken_predictReturn_T_2; 
  assign _taken_T_16=s2_valid&taken_predictReturn; 
  assign _GEN_45=~s2_btb_taken&_taken_T_16; 
  assign _GEN_78=_taken_T_45|_GEN_45; 
  assign _GEN_81=s2_btb_taken ? _GEN_45:_GEN_78; 
  assign useRAS=taken_idx ? _GEN_81:_GEN_45; 
  assign taken_rviBranch_1=taken_rviBits_1[6:0]==7'h63; 
  assign _taken_predictBranch_T_3=taken_prevRVI_1&taken_rviBranch_1; 
  assign _taken_rvcBranch_T_4=taken_bits_1&16'he003; 
  assign _taken_rvcBranch_T_5=16'hc001==_taken_rvcBranch_T_4; 
  assign _taken_rvcBranch_T_7=16'he001==_taken_rvcBranch_T_4; 
  assign taken_rvcBranch_1=_taken_rvcBranch_T_5|_taken_rvcBranch_T_7; 
  assign _taken_predictBranch_T_4=taken_valid_1&taken_rvcBranch_1; 
  assign _taken_predictBranch_T_5=_taken_predictBranch_T_3|_taken_predictBranch_T_4; 
  assign taken_predictBranch_1=s2_btb_resp_bits_bht_value&_taken_predictBranch_T_5; 
  assign taken_rviJump_1=taken_rviBits_1[6:0]==7'h6f; 
  assign _taken_predictJump_T_2=taken_prevRVI_1&taken_rviJump_1; 
  assign taken_rvcJump_1=16'ha001==_taken_rvcBranch_T_4; 
  assign _taken_predictJump_T_3=taken_valid_1&taken_rvcJump_1; 
  assign taken_predictJump_1=_taken_predictJump_T_2|_taken_predictJump_T_3; 
  assign _taken_T_46=taken_predictBranch_1|taken_predictJump_1; 
  assign _taken_T_47=s2_valid&_taken_T_46; 
  assign _s2_base_pc_T_1=~s2_pc|40'h3; 
  assign s2_base_pc=~_s2_base_pc_T_1; 
  assign taken_pc_1=s2_base_pc|40'h2; 
  assign _taken_npc_T_6=taken_pc_1-40'h2; 
  assign _taken_npc_T_8=taken_prevRVI_1 ? _taken_npc_T_6:taken_pc_1; 
  assign taken_rviImm_sign_2=taken_rviBits_1[31]; 
  assign taken_rviImm_hi_hi_hi_2=taken_rviBits_1[31]; 
  assign taken_rviImm_hi_hi_lo_2={11{taken_rviImm_sign_2}}; 
  assign taken_rviImm_hi_lo_hi_2=taken_rviBits_1[19:12]; 
  assign taken_rviImm_hi_lo_lo_2=taken_rviBits_1[20]; 
  assign taken_rviImm_lo_hi_hi_2=taken_rviBits_1[30:25]; 
  assign taken_rviImm_lo_hi_lo_2=taken_rviBits_1[24:21]; 
  assign _taken_rviImm_T_7={taken_rviImm_hi_hi_hi_2,taken_rviImm_hi_hi_lo_2,taken_rviImm_hi_lo_hi_2,taken_rviImm_hi_lo_lo_2,taken_rviImm_lo_hi_hi_2,taken_rviImm_lo_hi_lo_2,1'h0}; 
  assign taken_rviImm_hi_lo_hi_3={8{taken_rviImm_sign_2}}; 
  assign taken_rviImm_hi_lo_lo_3=taken_rviBits_1[7]; 
  assign _taken_rviImm_T_9={taken_rviImm_hi_hi_hi_2,taken_rviImm_hi_hi_lo_2,taken_rviImm_hi_lo_hi_3,taken_rviImm_hi_lo_lo_3,taken_rviImm_lo_hi_hi_2,taken_rviBits_1[11:8],1'h0}; 
  assign taken_rviImm_1=taken_rviBits_1[3] ? $signed(_taken_rviImm_T_7):$signed(_taken_rviImm_T_9); 
  assign taken_rvcImm_hi_hi_hi_2=taken_bits_1[12] ? 5'h1f:5'h0; 
  assign taken_rvcImm_hi_hi_lo_2=taken_bits_1[6:5]; 
  assign taken_rvcImm_hi_lo_2=taken_bits_1[2]; 
  assign taken_rvcImm_lo_hi_hi_2=taken_bits_1[11:10]; 
  assign taken_rvcImm_lo_hi_lo_2=taken_bits_1[4:3]; 
  assign _taken_rvcImm_T_13={taken_rvcImm_hi_hi_hi_2,taken_rvcImm_hi_hi_lo_2,taken_rvcImm_hi_lo_2,taken_rvcImm_lo_hi_hi_2,taken_rvcImm_lo_hi_lo_2,1'h0}; 
  assign taken_rvcImm_hi_hi_hi_hi_1=taken_bits_1[12] ? 10'h3ff:10'h0; 
  assign taken_rvcImm_hi_hi_hi_lo_1=taken_bits_1[8]; 
  assign taken_rvcImm_hi_hi_lo_3=taken_bits_1[10:9]; 
  assign taken_rvcImm_hi_lo_hi_1=taken_bits_1[6]; 
  assign taken_rvcImm_hi_lo_lo_1=taken_bits_1[7]; 
  assign taken_rvcImm_lo_hi_lo_3=taken_bits_1[11]; 
  assign taken_rvcImm_lo_lo_hi_1=taken_bits_1[5:3]; 
  assign _taken_rvcImm_T_17={taken_rvcImm_hi_hi_hi_hi_1,taken_rvcImm_hi_hi_hi_lo_1,taken_rvcImm_hi_hi_lo_3,taken_rvcImm_hi_lo_hi_1,taken_rvcImm_hi_lo_lo_1,taken_rvcImm_hi_lo_2,taken_rvcImm_lo_hi_lo_3,taken_rvcImm_lo_lo_hi_1,1'h0}; 
  assign taken_rvcImm_1=taken_bits_1[14] ? $signed({{8{_taken_rvcImm_T_13[12]}},_taken_rvcImm_T_13}):$signed(_taken_rvcImm_T_17); 
  assign _taken_npc_T_9=taken_prevRVI_1 ? $signed(taken_rviImm_1):$signed({{11{taken_rvcImm_1[20]}},taken_rvcImm_1}); 
  assign _GEN_127={{8{_taken_npc_T_9[31]}},_taken_npc_T_9}; 
  assign _taken_predicted_npc_T_1=$signed(_taken_npc_T_8)+$signed(_GEN_127); 
  assign _taken_predictBranch_T=taken_prevRVI&taken_rviBranch; 
  assign _taken_predictBranch_T_1=taken_valid&taken_rvcBranch; 
  assign _taken_predictBranch_T_2=_taken_predictBranch_T|_taken_predictBranch_T_1; 
  assign taken_predictBranch=s2_btb_resp_bits_bht_value&_taken_predictBranch_T_2; 
  assign _taken_predictJump_T=taken_prevRVI&taken_rviJump; 
  assign _taken_predictJump_T_1=taken_valid&taken_rvcJump; 
  assign taken_predictJump=_taken_predictJump_T|_taken_predictJump_T_1; 
  assign _taken_T_17=taken_predictBranch|taken_predictJump; 
  assign _taken_T_18=s2_valid&_taken_T_17; 
  assign _taken_npc_T=~_s2_base_pc_T_1; 
  assign taken_rviImm_sign=taken_rviBits[31]; 
  assign taken_rviImm_hi_hi_hi=taken_rviBits[31]; 
  assign taken_rviImm_hi_hi_lo={11{taken_rviImm_sign}}; 
  assign taken_rviImm_hi_lo_hi=taken_rviBits[19:12]; 
  assign taken_rviImm_hi_lo_lo=taken_rviBits[20]; 
  assign taken_rviImm_lo_hi_hi=taken_rviBits[30:25]; 
  assign taken_rviImm_lo_hi_lo=taken_rviBits[24:21]; 
  assign _taken_rviImm_T_2={taken_rviImm_hi_hi_hi,taken_rviImm_hi_hi_lo,taken_rviImm_hi_lo_hi,taken_rviImm_hi_lo_lo,taken_rviImm_lo_hi_hi,taken_rviImm_lo_hi_lo,1'h0}; 
  assign taken_rviImm_hi_lo_hi_1={8{taken_rviImm_sign}}; 
  assign taken_rviImm_hi_lo_lo_1=taken_rviBits[7]; 
  assign _taken_rviImm_T_4={taken_rviImm_hi_hi_hi,taken_rviImm_hi_hi_lo,taken_rviImm_hi_lo_hi_1,taken_rviImm_hi_lo_lo_1,taken_rviImm_lo_hi_hi,taken_rviBits[11:8],1'h0}; 
  assign taken_rviImm=taken_rviBits[3] ? $signed(_taken_rviImm_T_2):$signed(_taken_rviImm_T_4); 
  assign _taken_npc_T_1=$signed(taken_rviImm)-32'sh2; 
  assign taken_rvcImm_hi_hi_hi=taken_bits[12] ? 5'h1f:5'h0; 
  assign taken_rvcImm_hi_hi_lo=taken_bits[6:5]; 
  assign taken_rvcImm_hi_lo=taken_bits[2]; 
  assign taken_rvcImm_lo_hi_hi=taken_bits[11:10]; 
  assign taken_rvcImm_lo_hi_lo=taken_bits[4:3]; 
  assign _taken_rvcImm_T_4={taken_rvcImm_hi_hi_hi,taken_rvcImm_hi_hi_lo,taken_rvcImm_hi_lo,taken_rvcImm_lo_hi_hi,taken_rvcImm_lo_hi_lo,1'h0}; 
  assign taken_rvcImm_hi_hi_hi_hi=taken_bits[12] ? 10'h3ff:10'h0; 
  assign taken_rvcImm_hi_hi_hi_lo=taken_bits[8]; 
  assign taken_rvcImm_hi_hi_lo_1=taken_bits[10:9]; 
  assign taken_rvcImm_hi_lo_hi=taken_bits[6]; 
  assign taken_rvcImm_hi_lo_lo=taken_bits[7]; 
  assign taken_rvcImm_lo_hi_lo_1=taken_bits[11]; 
  assign taken_rvcImm_lo_lo_hi=taken_bits[5:3]; 
  assign _taken_rvcImm_T_8={taken_rvcImm_hi_hi_hi_hi,taken_rvcImm_hi_hi_hi_lo,taken_rvcImm_hi_hi_lo_1,taken_rvcImm_hi_lo_hi,taken_rvcImm_hi_lo_lo,taken_rvcImm_hi_lo,taken_rvcImm_lo_hi_lo_1,taken_rvcImm_lo_lo_hi,1'h0}; 
  assign taken_rvcImm=taken_bits[14] ? $signed({{8{_taken_rvcImm_T_4[12]}},_taken_rvcImm_T_4}):$signed(_taken_rvcImm_T_8); 
  assign _taken_npc_T_2=taken_prevRVI ? $signed(_taken_npc_T_1):$signed({{12{taken_rvcImm[20]}},taken_rvcImm}); 
  assign _GEN_128={{7{_taken_npc_T_2[32]}},_taken_npc_T_2}; 
  assign _taken_predicted_npc_T=$signed(_taken_npc_T)+$signed(_GEN_128); 
  assign predicted_taken=btb_io_resp_valid&btb_io_resp_bits_taken; 
  assign predicted_npc_hi=btb_io_resp_bits_target[38]; 
  assign _predicted_npc_T={predicted_npc_hi,btb_io_resp_bits_target}; 
  assign _GEN_28=predicted_taken ? _predicted_npc_T:ntpc; 
  assign _GEN_43=_taken_T_18 ? _taken_predicted_npc_T:_GEN_28; 
  assign _GEN_46=s2_btb_taken ? _GEN_28:_GEN_43; 
  assign _GEN_79=_taken_T_47 ? _taken_predicted_npc_T_1:_GEN_46; 
  assign _GEN_82=s2_btb_taken ? _GEN_46:_GEN_79; 
  assign _GEN_99=taken_idx ? _GEN_82:_GEN_46; 
  assign predicted_npc=useRAS ? {1'b0,btb_io_ras_head_bits}:_GEN_99; 
  assign npc=s2_replay ? s2_pc:predicted_npc; 
  assign _s0_speculative_T_1=s2_valid&~s2_speculative; 
  assign _s0_speculative_T_2=s1_speculative|_s0_speculative_T_1; 
  assign s0_speculative=_s0_speculative_T_2|predicted_taken; 
  assign _taken_taken_T_9=taken_rviJump_1|taken_rviJALR_1; 
  assign _taken_taken_T_10=taken_rviBranch_1&s2_btb_resp_bits_bht_value; 
  assign _taken_taken_T_11=_taken_taken_T_9|_taken_taken_T_10; 
  assign _taken_taken_T_12=taken_prevRVI_1&_taken_taken_T_11; 
  assign _taken_rvcJALR_T_5=16'h9002==_taken_rvcJR_T_4; 
  assign taken_rvcJALR_1=_taken_rvcJALR_T_5&_taken_rvcJR_T_7; 
  assign _taken_taken_T_13=taken_rvcJump_1|taken_rvcJALR_1; 
  assign _taken_taken_T_14=_taken_taken_T_13|taken_rvcJR_1; 
  assign _taken_taken_T_15=taken_rvcBranch_1&s2_btb_resp_bits_bht_value; 
  assign _taken_taken_T_16=_taken_taken_T_14|_taken_taken_T_15; 
  assign _taken_taken_T_17=taken_valid_1&_taken_taken_T_16; 
  assign taken_taken_1=_taken_taken_T_12|_taken_taken_T_17; 
  assign taken=taken_taken|taken_taken_1; 
  assign _GEN_116=_s2_replay_T|io_cpu_req_valid; 
  assign _GEN_120=taken ? _GEN_116:io_cpu_req_valid; 
  assign s2_redirect=s2_btb_taken ? io_cpu_req_valid:_GEN_120; 
  assign _GEN_0=~s2_replay&~s2_redirect; 
  assign _icache_io_s1_kill_T=s2_redirect|tlb_io_resp_miss; 
  assign s2_can_speculatively_refill=s2_tlb_resp_cacheable&~io_ptw_customCSRs_csrs_0_value[3]; 
  assign _icache_io_s2_kill_T_1=s2_speculative&~s2_can_speculatively_refill; 
  assign _fq_io_enq_valid_T=fq_io_enq_valid_REG&s2_valid; 
  assign _fq_io_enq_valid_T_2=~s2_tlb_resp_miss&icache_io_s2_kill; 
  assign _fq_io_enq_valid_T_3=icache_io_resp_valid|_fq_io_enq_valid_T_2; 
  assign _io_cpu_npc_T=io_cpu_req_valid ? io_cpu_req_bits_pc:npc; 
  assign _io_cpu_npc_T_2=~_io_cpu_npc_T|40'h1; 
  assign _fq_io_enq_bits_mask_T_1=3'h3<<s2_pc[1]; 
  assign _fq_io_enq_bits_replay_T_1=icache_io_s2_kill&~icache_io_resp_valid; 
  assign _fq_io_enq_bits_replay_T_3=_fq_io_enq_bits_replay_T_1&~s2_xcpt; 
  assign _fq_io_enq_bits_replay_T_4=icache_io_resp_bits_replay|_fq_io_enq_bits_replay_T_3; 
  assign _T_13=s2_speculative&io_ptw_customCSRs_csrs_0_value[3]; 
  assign _T_15=_T_13&~icache_io_s2_kill; 
  assign _T_18=~_T_15|reset; 
  assign _T_20=icache_io_resp_valid&icache_io_resp_bits_ae; 
  assign fetch_bubble_likely=~fq_io_mask[1]; 
  assign _btb_io_btb_update_valid_T_2=_s2_replay_T&~wrong_path; 
  assign _btb_io_btb_update_valid_T_3=_btb_io_btb_update_valid_T_2&fetch_bubble_likely; 
  assign _taken_T_53=taken_predictBranch_1&s2_btb_resp_bits_bht_value; 
  assign _taken_T_54=_taken_T_53|taken_predictJump_1; 
  assign _taken_T_55=_taken_T_54|taken_predictReturn_1; 
  assign _taken_T_56=~s2_btb_resp_valid&_taken_T_55; 
  assign _taken_T_24=taken_predictBranch&s2_btb_resp_bits_bht_value; 
  assign _taken_T_25=_taken_T_24|taken_predictJump; 
  assign _taken_T_26=_taken_T_25|taken_predictReturn; 
  assign _taken_T_27=~s2_btb_resp_valid&_taken_T_26; 
  assign _GEN_92=_taken_T_56|_taken_T_27; 
  assign updateBTB=taken_idx ? _GEN_92:_taken_T_27; 
  assign _btb_io_btb_update_valid_T_4=_btb_io_btb_update_valid_T_3&updateBTB; 
  assign _btb_io_btb_update_bits_br_pc_T={taken_idx,1'h0}; 
  assign _GEN_129={38'b0,_btb_io_btb_update_bits_br_pc_T}; 
  assign _btb_io_btb_update_bits_br_pc_T_1=s2_base_pc|_GEN_129; 
  assign _GEN_36=io_cpu_btb_update_valid ? {1'b0,io_cpu_btb_update_bits_br_pc}:_btb_io_btb_update_bits_br_pc_T_1; 
  assign _GEN_37=io_cpu_btb_update_valid ? {1'b0,io_cpu_btb_update_bits_pc}:s2_base_pc; 
  assign after_idx=taken_idx ? 2'h2:2'h1; 
  assign _btb_io_ras_update_bits_returnAddr_T={after_idx,1'h0}; 
  assign _GEN_130={37'b0,_btb_io_ras_update_bits_returnAddr_T}; 
  assign _btb_io_ras_update_bits_returnAddr_T_2=s2_base_pc+_GEN_130; 
  assign _taken_rviCall_T=taken_rviJALR|taken_rviJump; 
  assign taken_rviCall=_taken_rviCall_T&taken_rviBits[7]; 
  assign _taken_T=s2_valid&s2_btb_resp_valid; 
  assign _taken_T_2=_taken_T&~s2_btb_resp_bits_bridx; 
  assign _taken_T_3=_taken_T_2&taken_valid; 
  assign _taken_T_5=_taken_T_3&~_taken_prevRVI_T_4; 
  assign _GEN_39=_taken_T_5|_fq_io_enq_bits_replay_T_4; 
  assign _GEN_40=_taken_T_5|wrong_path; 
  assign _taken_btb_io_ras_update_valid_T_3=taken_rviCall|taken_rviReturn; 
  assign _taken_btb_io_ras_update_valid_T_4=taken_prevRVI&_taken_btb_io_ras_update_valid_T_3; 
  assign _taken_btb_io_ras_update_valid_T_5=taken_rvcJALR|taken_rvcReturn; 
  assign _taken_btb_io_ras_update_valid_T_6=taken_valid&_taken_btb_io_ras_update_valid_T_5; 
  assign _taken_btb_io_ras_update_valid_T_7=_taken_btb_io_ras_update_valid_T_4|_taken_btb_io_ras_update_valid_T_6; 
  assign _taken_btb_io_ras_update_valid_T_8=_btb_io_btb_update_valid_T_2&_taken_btb_io_ras_update_valid_T_7; 
  assign _taken_btb_io_ras_update_bits_cfiType_T=taken_prevRVI ? taken_rviReturn:taken_rvcReturn; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_1=taken_prevRVI ? taken_rviCall:taken_rvcJALR; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_2=taken_prevRVI ? taken_rviBranch:taken_rvcBranch; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_5=_taken_btb_io_ras_update_bits_cfiType_T_2 ? 1'h0:1'h1; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_6=_taken_btb_io_ras_update_bits_cfiType_T_1 ? 2'h2:{1'b0,_taken_btb_io_ras_update_bits_cfiType_T_5}; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_7=_taken_btb_io_ras_update_bits_cfiType_T ? 2'h3:_taken_btb_io_ras_update_bits_cfiType_T_6; 
  assign _taken_T_9=_s2_replay_T&taken_taken; 
  assign _taken_T_11=_taken_T_9&~taken_predictBranch; 
  assign _taken_T_13=_taken_T_11&~taken_predictJump; 
  assign _taken_T_15=_taken_T_13&~taken_predictReturn; 
  assign _GEN_41=_taken_T_15|_GEN_40; 
  assign _GEN_44=s2_btb_taken ? _GEN_40:_GEN_41; 
  assign _GEN_47=_taken_predictBranch_T_2&_btb_io_btb_update_valid_T_2; 
  assign taken_rvc_1=taken_bits_1[1:0]!=2'h3; 
  assign _taken_rviCall_T_2=taken_rviJALR_1|taken_rviJump_1; 
  assign taken_rviCall_1=_taken_rviCall_T_2&taken_rviBits_1[7]; 
  assign _taken_T_31=_taken_T&s2_btb_resp_bits_bridx; 
  assign _taken_T_32=_taken_T_31&taken_valid_1; 
  assign _taken_T_34=_taken_T_32&~taken_rvc_1; 
  assign _GEN_76=_taken_T_34|_GEN_44; 
  assign _taken_btb_io_ras_update_valid_T_12=taken_rviCall_1|taken_rviReturn_1; 
  assign _taken_btb_io_ras_update_valid_T_13=taken_prevRVI_1&_taken_btb_io_ras_update_valid_T_12; 
  assign _taken_btb_io_ras_update_valid_T_14=taken_rvcJALR_1|taken_rvcReturn_1; 
  assign _taken_btb_io_ras_update_valid_T_15=taken_valid_1&_taken_btb_io_ras_update_valid_T_14; 
  assign _taken_btb_io_ras_update_valid_T_16=_taken_btb_io_ras_update_valid_T_13|_taken_btb_io_ras_update_valid_T_15; 
  assign _taken_btb_io_ras_update_valid_T_17=_btb_io_btb_update_valid_T_2&_taken_btb_io_ras_update_valid_T_16; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_8=taken_prevRVI_1 ? taken_rviReturn_1:taken_rvcReturn_1; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_9=taken_prevRVI_1 ? taken_rviCall_1:taken_rvcJALR_1; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_10=taken_prevRVI_1 ? taken_rviBranch_1:taken_rvcBranch_1; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_13=_taken_btb_io_ras_update_bits_cfiType_T_10 ? 1'h0:1'h1; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_14=_taken_btb_io_ras_update_bits_cfiType_T_9 ? 2'h2:{1'b0,_taken_btb_io_ras_update_bits_cfiType_T_13}; 
  assign _taken_btb_io_ras_update_bits_cfiType_T_15=_taken_btb_io_ras_update_bits_cfiType_T_8 ? 2'h3:_taken_btb_io_ras_update_bits_cfiType_T_14; 
  assign _taken_T_38=_s2_replay_T&taken_taken_1; 
  assign _taken_T_40=_taken_T_38&~taken_predictBranch_1; 
  assign _taken_T_42=_taken_T_40&~taken_predictJump_1; 
  assign _taken_T_44=_taken_T_42&~taken_predictReturn_1; 
  assign _GEN_77=_taken_T_44|_GEN_76; 
  assign _GEN_83=_taken_predictBranch_T_5 ? _btb_io_btb_update_valid_T_2:_GEN_47; 
  assign _taken_T_59=taken_valid_1&taken_idx; 
  assign _taken_T_61=_taken_T_59&~taken_rvc_1; 
  assign _taken_lo_T=taken_bits_1|16'h3; 
  assign _T_25=s2_btb_taken|taken; 
  assign _T_26=_s2_replay_T&_T_25; 
  assign _GEN_117=taken ? taken_idx:s2_btb_resp_bits_bridx; 
  assign _GEN_118=taken|s2_btb_taken; 
  assign _GEN_119=taken ? 5'h1c:s2_btb_resp_bits_entry; 
  assign _T_31=~s2_partial_insn_valid|fq_io_enq_bits_mask[0]; 
  assign _T_33=_T_31|reset; 
  assign auto_icache_master_out_a_valid=icache_auto_master_out_a_valid; 
  assign auto_icache_master_out_a_bits_address=icache_auto_master_out_a_bits_address; 
  assign io_cpu_resp_valid=fq_io_deq_valid; 
  assign io_cpu_resp_bits_btb_taken=fq_io_deq_bits_btb_taken; 
  assign io_cpu_resp_bits_btb_bridx=fq_io_deq_bits_btb_bridx; 
  assign io_cpu_resp_bits_btb_entry=fq_io_deq_bits_btb_entry; 
  assign io_cpu_resp_bits_btb_bht_history=fq_io_deq_bits_btb_bht_history; 
  assign io_cpu_resp_bits_pc=fq_io_deq_bits_pc; 
  assign io_cpu_resp_bits_data=fq_io_deq_bits_data; 
  assign io_cpu_resp_bits_xcpt_pf_inst=fq_io_deq_bits_xcpt_pf_inst; 
  assign io_cpu_resp_bits_xcpt_ae_inst=fq_io_deq_bits_xcpt_ae_inst; 
  assign io_cpu_resp_bits_replay=fq_io_deq_bits_replay; 
  assign io_cpu_npc=~_io_cpu_npc_T_2; 
  assign io_ptw_req_valid=tlb_io_ptw_req_valid; 
  assign io_ptw_req_bits_valid=tlb_io_ptw_req_bits_valid; 
  assign io_ptw_req_bits_bits_addr=tlb_io_ptw_req_bits_bits_addr; 
  assign icache_clock=gated_clock; 
  assign icache_reset=reset; 
  assign icache_auto_master_out_a_ready=auto_icache_master_out_a_ready; 
  assign icache_auto_master_out_d_valid=auto_icache_master_out_d_valid; 
  assign icache_auto_master_out_d_bits_opcode=auto_icache_master_out_d_bits_opcode; 
  assign icache_auto_master_out_d_bits_size=auto_icache_master_out_d_bits_size; 
  assign icache_auto_master_out_d_bits_data=auto_icache_master_out_d_bits_data; 
  assign icache_auto_master_out_d_bits_corrupt=auto_icache_master_out_d_bits_corrupt; 
  assign icache_io_req_valid=io_cpu_req_valid|s0_fq_has_space; 
  assign icache_io_req_bits_addr=io_cpu_npc[38:0]; 
  assign icache_io_s1_paddr=tlb_io_resp_paddr; 
  assign icache_io_s1_kill=_icache_io_s1_kill_T|s2_replay; 
  assign icache_io_s2_kill=_icache_io_s2_kill_T_1|s2_xcpt; 
  assign icache_io_invalidate=io_cpu_flush_icache; 
  assign fq_clock=gated_clock; 
  assign fq_reset=reset|io_cpu_req_valid; 
  assign fq_io_enq_valid=_fq_io_enq_valid_T&_fq_io_enq_valid_T_3; 
  assign fq_io_enq_bits_btb_taken=s2_btb_taken ? s2_btb_taken:_GEN_118; 
  assign fq_io_enq_bits_btb_bridx=s2_btb_taken ? s2_btb_resp_bits_bridx:_GEN_117; 
  assign fq_io_enq_bits_btb_entry=s2_btb_taken ? s2_btb_resp_bits_entry:_GEN_119; 
  assign fq_io_enq_bits_btb_bht_history=s2_btb_resp_bits_bht_history; 
  assign fq_io_enq_bits_pc=s2_pc; 
  assign fq_io_enq_bits_data=icache_io_resp_bits_data; 
  assign fq_io_enq_bits_mask=_fq_io_enq_bits_mask_T_1[1:0]; 
  assign fq_io_enq_bits_xcpt_pf_inst=s2_tlb_resp_pf_inst; 
  assign fq_io_enq_bits_xcpt_ae_inst=_T_20|s2_tlb_resp_ae_inst; 
  assign fq_io_enq_bits_replay=_taken_T_34|_GEN_39; 
  assign fq_io_deq_ready=io_cpu_resp_ready; 
  assign tlb_clock=gated_clock; 
  assign tlb_reset=reset; 
  assign tlb_io_req_valid=s1_valid&~s2_replay; 
  assign tlb_io_req_bits_vaddr=s1_pc; 
  assign tlb_io_sfence_valid=io_cpu_sfence_valid; 
  assign tlb_io_sfence_bits_rs1=io_cpu_sfence_bits_rs1; 
  assign tlb_io_sfence_bits_rs2=io_cpu_sfence_bits_rs2; 
  assign tlb_io_sfence_bits_addr=io_cpu_sfence_bits_addr; 
  assign tlb_io_ptw_req_ready=io_ptw_req_ready; 
  assign tlb_io_ptw_resp_valid=io_ptw_resp_valid; 
  assign tlb_io_ptw_resp_bits_ae=io_ptw_resp_bits_ae; 
  assign tlb_io_ptw_resp_bits_pte_ppn=io_ptw_resp_bits_pte_ppn; 
  assign tlb_io_ptw_resp_bits_pte_d=io_ptw_resp_bits_pte_d; 
  assign tlb_io_ptw_resp_bits_pte_a=io_ptw_resp_bits_pte_a; 
  assign tlb_io_ptw_resp_bits_pte_g=io_ptw_resp_bits_pte_g; 
  assign tlb_io_ptw_resp_bits_pte_u=io_ptw_resp_bits_pte_u; 
  assign tlb_io_ptw_resp_bits_pte_x=io_ptw_resp_bits_pte_x; 
  assign tlb_io_ptw_resp_bits_pte_w=io_ptw_resp_bits_pte_w; 
  assign tlb_io_ptw_resp_bits_pte_r=io_ptw_resp_bits_pte_r; 
  assign tlb_io_ptw_resp_bits_pte_v=io_ptw_resp_bits_pte_v; 
  assign tlb_io_ptw_resp_bits_level=io_ptw_resp_bits_level; 
  assign tlb_io_ptw_resp_bits_homogeneous=io_ptw_resp_bits_homogeneous; 
  assign tlb_io_ptw_ptbr_mode=io_ptw_ptbr_mode; 
  assign tlb_io_ptw_status_debug=io_ptw_status_debug; 
  assign tlb_io_ptw_status_prv=io_ptw_status_prv; 
  assign tlb_io_ptw_pmp_0_cfg_l=io_ptw_pmp_0_cfg_l; 
  assign tlb_io_ptw_pmp_0_cfg_a=io_ptw_pmp_0_cfg_a; 
  assign tlb_io_ptw_pmp_0_cfg_x=io_ptw_pmp_0_cfg_x; 
  assign tlb_io_ptw_pmp_0_cfg_w=io_ptw_pmp_0_cfg_w; 
  assign tlb_io_ptw_pmp_0_cfg_r=io_ptw_pmp_0_cfg_r; 
  assign tlb_io_ptw_pmp_0_addr=io_ptw_pmp_0_addr; 
  assign tlb_io_ptw_pmp_0_mask=io_ptw_pmp_0_mask; 
  assign tlb_io_ptw_pmp_1_cfg_l=io_ptw_pmp_1_cfg_l; 
  assign tlb_io_ptw_pmp_1_cfg_a=io_ptw_pmp_1_cfg_a; 
  assign tlb_io_ptw_pmp_1_cfg_x=io_ptw_pmp_1_cfg_x; 
  assign tlb_io_ptw_pmp_1_cfg_w=io_ptw_pmp_1_cfg_w; 
  assign tlb_io_ptw_pmp_1_cfg_r=io_ptw_pmp_1_cfg_r; 
  assign tlb_io_ptw_pmp_1_addr=io_ptw_pmp_1_addr; 
  assign tlb_io_ptw_pmp_1_mask=io_ptw_pmp_1_mask; 
  assign tlb_io_ptw_pmp_2_cfg_l=io_ptw_pmp_2_cfg_l; 
  assign tlb_io_ptw_pmp_2_cfg_a=io_ptw_pmp_2_cfg_a; 
  assign tlb_io_ptw_pmp_2_cfg_x=io_ptw_pmp_2_cfg_x; 
  assign tlb_io_ptw_pmp_2_cfg_w=io_ptw_pmp_2_cfg_w; 
  assign tlb_io_ptw_pmp_2_cfg_r=io_ptw_pmp_2_cfg_r; 
  assign tlb_io_ptw_pmp_2_addr=io_ptw_pmp_2_addr; 
  assign tlb_io_ptw_pmp_2_mask=io_ptw_pmp_2_mask; 
  assign tlb_io_ptw_pmp_3_cfg_l=io_ptw_pmp_3_cfg_l; 
  assign tlb_io_ptw_pmp_3_cfg_a=io_ptw_pmp_3_cfg_a; 
  assign tlb_io_ptw_pmp_3_cfg_x=io_ptw_pmp_3_cfg_x; 
  assign tlb_io_ptw_pmp_3_cfg_w=io_ptw_pmp_3_cfg_w; 
  assign tlb_io_ptw_pmp_3_cfg_r=io_ptw_pmp_3_cfg_r; 
  assign tlb_io_ptw_pmp_3_addr=io_ptw_pmp_3_addr; 
  assign tlb_io_ptw_pmp_3_mask=io_ptw_pmp_3_mask; 
  assign tlb_io_ptw_pmp_4_cfg_l=io_ptw_pmp_4_cfg_l; 
  assign tlb_io_ptw_pmp_4_cfg_a=io_ptw_pmp_4_cfg_a; 
  assign tlb_io_ptw_pmp_4_cfg_x=io_ptw_pmp_4_cfg_x; 
  assign tlb_io_ptw_pmp_4_cfg_w=io_ptw_pmp_4_cfg_w; 
  assign tlb_io_ptw_pmp_4_cfg_r=io_ptw_pmp_4_cfg_r; 
  assign tlb_io_ptw_pmp_4_addr=io_ptw_pmp_4_addr; 
  assign tlb_io_ptw_pmp_4_mask=io_ptw_pmp_4_mask; 
  assign tlb_io_ptw_pmp_5_cfg_l=io_ptw_pmp_5_cfg_l; 
  assign tlb_io_ptw_pmp_5_cfg_a=io_ptw_pmp_5_cfg_a; 
  assign tlb_io_ptw_pmp_5_cfg_x=io_ptw_pmp_5_cfg_x; 
  assign tlb_io_ptw_pmp_5_cfg_w=io_ptw_pmp_5_cfg_w; 
  assign tlb_io_ptw_pmp_5_cfg_r=io_ptw_pmp_5_cfg_r; 
  assign tlb_io_ptw_pmp_5_addr=io_ptw_pmp_5_addr; 
  assign tlb_io_ptw_pmp_5_mask=io_ptw_pmp_5_mask; 
  assign tlb_io_ptw_pmp_6_cfg_l=io_ptw_pmp_6_cfg_l; 
  assign tlb_io_ptw_pmp_6_cfg_a=io_ptw_pmp_6_cfg_a; 
  assign tlb_io_ptw_pmp_6_cfg_x=io_ptw_pmp_6_cfg_x; 
  assign tlb_io_ptw_pmp_6_cfg_w=io_ptw_pmp_6_cfg_w; 
  assign tlb_io_ptw_pmp_6_cfg_r=io_ptw_pmp_6_cfg_r; 
  assign tlb_io_ptw_pmp_6_addr=io_ptw_pmp_6_addr; 
  assign tlb_io_ptw_pmp_6_mask=io_ptw_pmp_6_mask; 
  assign tlb_io_ptw_pmp_7_cfg_l=io_ptw_pmp_7_cfg_l; 
  assign tlb_io_ptw_pmp_7_cfg_a=io_ptw_pmp_7_cfg_a; 
  assign tlb_io_ptw_pmp_7_cfg_x=io_ptw_pmp_7_cfg_x; 
  assign tlb_io_ptw_pmp_7_cfg_w=io_ptw_pmp_7_cfg_w; 
  assign tlb_io_ptw_pmp_7_cfg_r=io_ptw_pmp_7_cfg_r; 
  assign tlb_io_ptw_pmp_7_addr=io_ptw_pmp_7_addr; 
  assign tlb_io_ptw_pmp_7_mask=io_ptw_pmp_7_mask; 
  assign tlb_io_kill=~s2_valid; 
  assign btb_clock=gated_clock; 
  assign btb_reset=reset; 
  assign btb_io_req_bits_addr=s1_pc[38:0]; 
  assign btb_io_btb_update_valid=io_cpu_btb_update_valid ? io_cpu_btb_update_valid:_btb_io_btb_update_valid_T_4; 
  assign btb_io_btb_update_bits_prediction_entry=io_cpu_btb_update_valid ? io_cpu_btb_update_bits_prediction_entry:5'h1c; 
  assign btb_io_btb_update_bits_pc=_GEN_37[38:0]; 
  assign btb_io_btb_update_bits_isValid=~io_cpu_btb_update_valid|io_cpu_btb_update_bits_isValid; 
  assign btb_io_btb_update_bits_br_pc=_GEN_36[38:0]; 
  assign btb_io_btb_update_bits_cfiType=io_cpu_btb_update_valid ? io_cpu_btb_update_bits_cfiType:btb_io_ras_update_bits_cfiType; 
  assign btb_io_bht_update_valid=io_cpu_bht_update_valid; 
  assign btb_io_bht_update_bits_prediction_history=io_cpu_bht_update_bits_prediction_history; 
  assign btb_io_bht_update_bits_pc=io_cpu_bht_update_bits_pc; 
  assign btb_io_bht_update_bits_branch=io_cpu_bht_update_bits_branch; 
  assign btb_io_bht_update_bits_taken=io_cpu_bht_update_bits_taken; 
  assign btb_io_bht_update_bits_mispredict=io_cpu_bht_update_bits_mispredict; 
  assign btb_io_bht_advance_valid=taken_idx ? _GEN_83:_GEN_47; 
  assign btb_io_bht_advance_bits_bht_value=s2_btb_resp_bits_bht_value; 
  assign btb_io_ras_update_valid=taken_idx ? _taken_btb_io_ras_update_valid_T_17:_taken_btb_io_ras_update_valid_T_8; 
  assign btb_io_ras_update_bits_cfiType=taken_idx ? _taken_btb_io_ras_update_bits_cfiType_T_15:_taken_btb_io_ras_update_bits_cfiType_T_7; 
  assign btb_io_ras_update_bits_returnAddr=_btb_io_ras_update_bits_returnAddr_T_2[38:0]; 
  assign btb_io_flush=_taken_T_34|_taken_T_5; 
  assign Frontend_cov_read_addr=Frontend_state; 
  assign Frontend_cov_read_data=Frontend_cov[Frontend_cov_read_addr]; 
  assign Frontend_cov_write_data=1'h1; 
  assign Frontend_cov_write_addr=Frontend_state; 
  assign Frontend_cov_write_mask=1'h1; 
  assign Frontend_cov_write_en=1'h1; 
  assign s2_partial_insn_valid_shl=s2_partial_insn_valid; 
  assign s2_partial_insn_valid_pad={5'h0,s2_partial_insn_valid_shl}; 
  assign s2_btb_resp_valid_shl={s2_btb_resp_valid,1'h0}; 
  assign s2_btb_resp_valid_pad={4'h0,s2_btb_resp_valid_shl}; 
  assign s2_replay_REG_shl={s2_replay_REG,2'h0}; 
  assign s2_replay_REG_pad={3'h0,s2_replay_REG_shl}; 
  assign s2_btb_resp_bits_bht_value_shl={s2_btb_resp_bits_bht_value,3'h0}; 
  assign s2_btb_resp_bits_bht_value_pad={2'h0,s2_btb_resp_bits_bht_value_shl}; 
  assign s2_valid_shl={s2_valid,4'h0}; 
  assign s2_valid_pad={1'h0,s2_valid_shl}; 
  assign s2_btb_resp_bits_taken_shl={s2_btb_resp_bits_taken,5'h0}; 
  assign s2_btb_resp_bits_taken_pad=s2_btb_resp_bits_taken_shl; 
  assign Frontend_xor4=s2_btb_resp_valid_pad^s2_replay_REG_pad; 
  assign Frontend_xor1=s2_partial_insn_valid_pad^Frontend_xor4; 
  assign Frontend_xor6=s2_valid_pad^s2_btb_resp_bits_taken_pad; 
  assign Frontend_xor2=s2_btb_resp_bits_bht_value_pad^Frontend_xor6; 
  assign Frontend_xor0=Frontend_xor1^Frontend_xor2; 
  assign icache_sum=Frontend_covSum+icache_io_covSum; 
  assign fq_sum=icache_sum+fq_io_covSum; 
  assign tlb_sum=fq_sum+tlb_io_covSum; 
  assign btb_sum=tlb_sum+btb_io_covSum; 
  assign io_covSum=btb_sum; 
  assign stopEn0=~_T_9; 
  assign stopEn1=~_T_18; 
  assign stopEn2=~_T_33; 
  assign icache_metaAssert_wire=icache_metaAssert; 
  assign fq_metaAssert_wire=fq_metaAssert; 
  assign tlb_metaAssert_wire=tlb_metaAssert; 
  assign btb_metaAssert_wire=btb_metaAssert; 
  assign Frontend_or4=stopEn1|stopEn2; 
  assign Frontend_or1=stopEn0|Frontend_or4; 
  assign Frontend_or5=icache_metaAssert_wire|fq_metaAssert_wire; 
  assign Frontend_or6=tlb_metaAssert_wire|btb_metaAssert_wire; 
  assign Frontend_or2=Frontend_or5|Frontend_or6; 
  assign Frontend_or0=Frontend_or1|Frontend_or2; 
  assign metaAssert=Frontend_or0; 
  assign icache_metaReset=metaReset|icache_halt; 
  assign fq_metaReset=metaReset|fq_halt; 
  assign tlb_metaReset=metaReset|tlb_halt; 
  assign btb_metaReset=metaReset|btb_halt; initial
    begin 
    end  
  always @( posedge gated_clock)
       begin 
         if (metaReset)
            begin 
              s1_valid <=1'h0;
            end 
          else 
            begin 
              s1_valid <=io_cpu_req_valid|s0_fq_has_space;
            end 
         if (metaReset)
            begin 
              s2_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s2_valid <=1'h0;
               end 
             else 
               begin 
                 s2_valid <=_GEN_0;
               end 
         if (metaReset)
            begin 
              s1_pc <=40'h0;
            end 
          else 
            begin 
              s1_pc <=io_cpu_npc;
            end 
         if (metaReset)
            begin 
              s1_speculative <=1'h0;
            end 
          else 
            if (io_cpu_req_valid)
               begin 
                 s1_speculative <=io_cpu_req_bits_speculative;
               end 
             else 
               if (s2_replay)
                  begin 
                    s1_speculative <=s2_speculative;
                  end 
                else 
                  begin 
                    s1_speculative <=s0_speculative;
                  end 
         if (metaReset)
            begin 
              s2_pc <=40'h0;
            end 
          else 
            if (reset)
               begin 
                 s2_pc <={8'b0,~_s2_pc_T_1};
               end 
             else 
               if (~s2_replay)
                  begin 
                    s2_pc <=s1_pc;
                  end 
         if (metaReset)
            begin 
              s2_btb_resp_valid <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_btb_resp_valid <=btb_io_resp_valid;
               end 
         if (metaReset)
            begin 
              s2_btb_resp_bits_taken <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_btb_resp_bits_taken <=btb_io_resp_bits_taken;
               end 
         if (metaReset)
            begin 
              s2_btb_resp_bits_bridx <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_btb_resp_bits_bridx <=btb_io_resp_bits_bridx;
               end 
         if (metaReset)
            begin 
              s2_btb_resp_bits_entry <=5'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_btb_resp_bits_entry <=btb_io_resp_bits_entry;
               end 
         if (metaReset)
            begin 
              s2_btb_resp_bits_bht_history <=8'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_btb_resp_bits_bht_history <=btb_io_resp_bits_bht_history;
               end 
         if (metaReset)
            begin 
              s2_btb_resp_bits_bht_value <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_btb_resp_bits_bht_value <=btb_io_resp_bits_bht_value;
               end 
         if (metaReset)
            begin 
              s2_tlb_resp_miss <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_tlb_resp_miss <=tlb_io_resp_miss;
               end 
         if (metaReset)
            begin 
              s2_tlb_resp_pf_inst <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_tlb_resp_pf_inst <=tlb_io_resp_pf_inst;
               end 
         if (metaReset)
            begin 
              s2_tlb_resp_ae_inst <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_tlb_resp_ae_inst <=tlb_io_resp_ae_inst;
               end 
         if (metaReset)
            begin 
              s2_tlb_resp_cacheable <=1'h0;
            end 
          else 
            if (~s2_replay)
               begin 
                 s2_tlb_resp_cacheable <=tlb_io_resp_cacheable;
               end 
         if (metaReset)
            begin 
              s2_speculative <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s2_speculative <=1'h0;
               end 
             else 
               if (~s2_replay)
                  begin 
                    s2_speculative <=s1_speculative;
                  end 
         if (metaReset)
            begin 
              s2_partial_insn_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s2_partial_insn_valid <=1'h0;
               end 
             else 
               if (s2_redirect)
                  begin 
                    s2_partial_insn_valid <=1'h0;
                  end 
                else 
                  if (_T_26)
                     begin 
                       s2_partial_insn_valid <=1'h0;
                     end 
                   else 
                     if (_s2_replay_T)
                        begin 
                          s2_partial_insn_valid <=_taken_T_61;
                        end 
         if (metaReset)
            begin 
              s2_partial_insn <=16'h0;
            end 
          else 
            if (_s2_replay_T)
               begin 
                 if (_taken_T_61)
                    begin 
                      s2_partial_insn <=_taken_lo_T;
                    end 
               end 
         if (metaReset)
            begin 
              wrong_path <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 wrong_path <=1'h0;
               end 
             else 
               if (io_cpu_req_valid)
                  begin 
                    wrong_path <=1'h0;
                  end 
                else 
                  if (taken_idx)
                     begin 
                       if (~s2_btb_taken)
                          begin 
                            wrong_path <=_GEN_77;
                          end 
                        else 
                          begin 
                            wrong_path <=_GEN_76;
                          end 
                     end 
                   else 
                     begin 
                       wrong_path <=_GEN_76;
                     end 
         if (metaReset)
            begin 
              s2_replay_REG <=1'h0;
            end 
          else 
            begin 
              s2_replay_REG <=reset|_s2_replay_T_4;
            end 
         if (metaReset)
            begin 
              fq_io_enq_valid_REG <=1'h0;
            end 
          else 
            begin 
              fq_io_enq_valid_REG <=s1_valid;
            end 
         if (~_T_9)
            begin $display("Assertion failed\n    at Frontend.scala:89 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n");
            end 
         if (~_T_9)
            begin $display("fatal");
            end 
         if (~_T_18)
            begin $display("Assertion failed\n    at Frontend.scala:175 assert(!(s2_speculative && io.ptw.customCSRs.asInstanceOf[RocketCustomCSRs].disableSpeculativeICacheRefill && !icache.io.s2_kill))\n");
            end 
         if (~_T_18)
            begin $display("fatal");
            end 
         if (~_T_33)
            begin $display("Assertion failed\n    at Frontend.scala:320 assert(!s2_partial_insn_valid || fq.io.enq.bits.mask(0))\n");
            end 
         if (~_T_33)
            begin $display("fatal");
            end 
         Frontend_state <=Frontend_xor0;
         if (!(Frontend_cov_read_data))
            begin 
              Frontend_covSum <=Frontend_covSum+1'h1;
            end 
       end
  
  always @( posedge gated_clock)
       begin 
         if (Frontend_cov_write_en&Frontend_cov_write_mask)
            begin 
              Frontend_cov [Frontend_cov_write_addr]<=Frontend_cov_write_data;
            end 
       end
  
endmodule
 
module FPU (
  input clock,
  input reset,
  input [31:0] io_inst,
  input [63:0] io_fromint_data,
  input [2:0] io_fcsr_rm,
  output io_fcsr_flags_valid,
  output [4:0] io_fcsr_flags_bits,
  output [63:0] io_store_data,
  output [63:0] io_toint_data,
  input io_dmem_resp_val,
  input [2:0] io_dmem_resp_type,
  input [4:0] io_dmem_resp_tag,
  input [63:0] io_dmem_resp_data,
  input io_valid,
  output io_fcsr_rdy,
  output io_nack_mem,
  output io_illegal_rm,
  input io_killx,
  input io_killm,
  output io_dec_wen,
  output io_dec_ren1,
  output io_dec_ren2,
  output io_dec_ren3,
  output io_sboard_set,
  output io_sboard_clr,
  output [4:0] io_sboard_clra,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input fpiu_halt,
  input ifpu_halt,
  input sfma_halt,
  input fpmu_halt,
  input divSqrt_1_halt,
  input dfma_halt,
  input divSqrt_halt) ; 
   wire [31:0] fp_decoder_io_inst ;  
   wire fp_decoder_io_sigs_wen ;  
   wire fp_decoder_io_sigs_ren1 ;  
   wire fp_decoder_io_sigs_ren2 ;  
   wire fp_decoder_io_sigs_ren3 ;  
   wire fp_decoder_io_sigs_swap12 ;  
   wire fp_decoder_io_sigs_swap23 ;  
   wire [1:0] fp_decoder_io_sigs_typeTagIn ;  
   wire [1:0] fp_decoder_io_sigs_typeTagOut ;  
   wire fp_decoder_io_sigs_fromint ;  
   wire fp_decoder_io_sigs_toint ;  
   wire fp_decoder_io_sigs_fastpipe ;  
   wire fp_decoder_io_sigs_fma ;  
   wire fp_decoder_io_sigs_div ;  
   wire fp_decoder_io_sigs_sqrt ;  
   wire fp_decoder_io_sigs_wflags ;  
   wire [29:0] fp_decoder_io_covSum ;  
   wire fp_decoder_metaAssert ;  
   reg [64:0] regfile[0:31] ;  
   reg [95:0] _RAND_0 ;  
   wire [64:0] regfile_ex_rs_0_data ;  
   wire [4:0] regfile_ex_rs_0_addr ;  
   wire [64:0] regfile_ex_rs_1_data ;  
   wire [4:0] regfile_ex_rs_1_addr ;  
   wire [64:0] regfile_ex_rs_2_data ;  
   wire [4:0] regfile_ex_rs_2_addr ;  
   wire [64:0] regfile_MPORT_data ;  
   wire [4:0] regfile_MPORT_addr ;  
   wire regfile_MPORT_mask ;  
   wire regfile_MPORT_en ;  
   wire [64:0] regfile_MPORT_1_data ;  
   wire [4:0] regfile_MPORT_1_addr ;  
   wire regfile_MPORT_1_mask ;  
   wire regfile_MPORT_1_en ;  
   wire sfma_clock ;  
   wire sfma_reset ;  
   wire sfma_io_in_valid ;  
   wire sfma_io_in_bits_ren3 ;  
   wire sfma_io_in_bits_swap23 ;  
   wire [2:0] sfma_io_in_bits_rm ;  
   wire [1:0] sfma_io_in_bits_fmaCmd ;  
   wire [64:0] sfma_io_in_bits_in1 ;  
   wire [64:0] sfma_io_in_bits_in2 ;  
   wire [64:0] sfma_io_in_bits_in3 ;  
   wire [64:0] sfma_io_out_bits_data ;  
   wire [4:0] sfma_io_out_bits_exc ;  
   wire [29:0] sfma_io_covSum ;  
   wire sfma_metaAssert ;  
   wire sfma_metaReset ;  
   wire sfma_fma_halt ;  
   wire fpiu_clock ;  
   wire fpiu_io_in_valid ;  
   wire fpiu_io_in_bits_ren2 ;  
   wire [1:0] fpiu_io_in_bits_typeTagIn ;  
   wire [1:0] fpiu_io_in_bits_typeTagOut ;  
   wire fpiu_io_in_bits_wflags ;  
   wire [2:0] fpiu_io_in_bits_rm ;  
   wire [1:0] fpiu_io_in_bits_typ ;  
   wire [1:0] fpiu_io_in_bits_fmt ;  
   wire [64:0] fpiu_io_in_bits_in1 ;  
   wire [64:0] fpiu_io_in_bits_in2 ;  
   wire [2:0] fpiu_io_out_bits_in_rm ;  
   wire [64:0] fpiu_io_out_bits_in_in1 ;  
   wire [64:0] fpiu_io_out_bits_in_in2 ;  
   wire fpiu_io_out_bits_lt ;  
   wire [63:0] fpiu_io_out_bits_store ;  
   wire [63:0] fpiu_io_out_bits_toint ;  
   wire [4:0] fpiu_io_out_bits_exc ;  
   wire [29:0] fpiu_io_covSum ;  
   wire fpiu_metaAssert ;  
   wire fpiu_metaReset ;  
   wire ifpu_clock ;  
   wire ifpu_reset ;  
   wire ifpu_io_in_valid ;  
   wire [1:0] ifpu_io_in_bits_typeTagIn ;  
   wire ifpu_io_in_bits_wflags ;  
   wire [2:0] ifpu_io_in_bits_rm ;  
   wire [1:0] ifpu_io_in_bits_typ ;  
   wire [63:0] ifpu_io_in_bits_in1 ;  
   wire [64:0] ifpu_io_out_bits_data ;  
   wire [4:0] ifpu_io_out_bits_exc ;  
   wire [29:0] ifpu_io_covSum ;  
   wire ifpu_metaAssert ;  
   wire ifpu_metaReset ;  
   wire fpmu_clock ;  
   wire fpmu_reset ;  
   wire fpmu_io_in_valid ;  
   wire fpmu_io_in_bits_ren2 ;  
   wire [1:0] fpmu_io_in_bits_typeTagOut ;  
   wire fpmu_io_in_bits_wflags ;  
   wire [2:0] fpmu_io_in_bits_rm ;  
   wire [64:0] fpmu_io_in_bits_in1 ;  
   wire [64:0] fpmu_io_in_bits_in2 ;  
   wire [64:0] fpmu_io_out_bits_data ;  
   wire [4:0] fpmu_io_out_bits_exc ;  
   wire fpmu_io_lt ;  
   wire [29:0] fpmu_io_covSum ;  
   wire fpmu_metaAssert ;  
   wire fpmu_metaReset ;  
   wire dfma_clock ;  
   wire dfma_reset ;  
   wire dfma_io_in_valid ;  
   wire dfma_io_in_bits_ren3 ;  
   wire dfma_io_in_bits_swap23 ;  
   wire [2:0] dfma_io_in_bits_rm ;  
   wire [1:0] dfma_io_in_bits_fmaCmd ;  
   wire [64:0] dfma_io_in_bits_in1 ;  
   wire [64:0] dfma_io_in_bits_in2 ;  
   wire [64:0] dfma_io_in_bits_in3 ;  
   wire [64:0] dfma_io_out_bits_data ;  
   wire [4:0] dfma_io_out_bits_exc ;  
   wire [29:0] dfma_io_covSum ;  
   wire dfma_metaAssert ;  
   wire dfma_metaReset ;  
   wire dfma_fma_halt ;  
   wire divSqrt_clock ;  
   wire divSqrt_reset ;  
   wire divSqrt_io_inReady ;  
   wire divSqrt_io_inValid ;  
   wire divSqrt_io_sqrtOp ;  
   wire [32:0] divSqrt_io_a ;  
   wire [32:0] divSqrt_io_b ;  
   wire [2:0] divSqrt_io_roundingMode ;  
   wire divSqrt_io_outValid_div ;  
   wire divSqrt_io_outValid_sqrt ;  
   wire [32:0] divSqrt_io_out ;  
   wire [4:0] divSqrt_io_exceptionFlags ;  
   wire [29:0] divSqrt_io_covSum ;  
   wire divSqrt_metaAssert ;  
   wire divSqrt_metaReset ;  
   wire divSqrt_divSqrtRecFNToRaw_halt ;  
   wire divSqrt_1_clock ;  
   wire divSqrt_1_reset ;  
   wire divSqrt_1_io_inReady ;  
   wire divSqrt_1_io_inValid ;  
   wire divSqrt_1_io_sqrtOp ;  
   wire [64:0] divSqrt_1_io_a ;  
   wire [64:0] divSqrt_1_io_b ;  
   wire [2:0] divSqrt_1_io_roundingMode ;  
   wire divSqrt_1_io_outValid_div ;  
   wire divSqrt_1_io_outValid_sqrt ;  
   wire [64:0] divSqrt_1_io_out ;  
   wire [4:0] divSqrt_1_io_exceptionFlags ;  
   wire [29:0] divSqrt_1_io_covSum ;  
   wire divSqrt_1_metaAssert ;  
   wire divSqrt_1_metaReset ;  
   wire divSqrt_1_divSqrtRecFNToRaw_halt ;  
   reg ex_reg_valid ;  
   reg [31:0] _RAND_1 ;  
   reg [31:0] ex_reg_inst ;  
   reg [31:0] _RAND_2 ;  
   reg ex_reg_ctrl_ren2 ;  
   reg [31:0] _RAND_3 ;  
   reg ex_reg_ctrl_ren3 ;  
   reg [31:0] _RAND_4 ;  
   reg ex_reg_ctrl_swap23 ;  
   reg [31:0] _RAND_5 ;  
   reg [1:0] ex_reg_ctrl_typeTagIn ;  
   reg [31:0] _RAND_6 ;  
   reg [1:0] ex_reg_ctrl_typeTagOut ;  
   reg [31:0] _RAND_7 ;  
   reg ex_reg_ctrl_fromint ;  
   reg [31:0] _RAND_8 ;  
   reg ex_reg_ctrl_toint ;  
   reg [31:0] _RAND_9 ;  
   reg ex_reg_ctrl_fastpipe ;  
   reg [31:0] _RAND_10 ;  
   reg ex_reg_ctrl_fma ;  
   reg [31:0] _RAND_11 ;  
   reg ex_reg_ctrl_div ;  
   reg [31:0] _RAND_12 ;  
   reg ex_reg_ctrl_sqrt ;  
   reg [31:0] _RAND_13 ;  
   reg ex_reg_ctrl_wflags ;  
   reg [31:0] _RAND_14 ;  
   reg [4:0] ex_ra_0 ;  
   reg [31:0] _RAND_15 ;  
   reg [4:0] ex_ra_1 ;  
   reg [31:0] _RAND_16 ;  
   reg [4:0] ex_ra_2 ;  
   reg [31:0] _RAND_17 ;  
   reg load_wb ;  
   reg [31:0] _RAND_18 ;  
   wire [1:0] _load_wb_typeTag_T_2 ;  
   reg [1:0] load_wb_typeTag ;  
   reg [31:0] _RAND_19 ;  
   reg [63:0] load_wb_data ;  
   reg [63:0] _RAND_20 ;  
   reg [4:0] load_wb_tag ;  
   reg [31:0] _RAND_21 ;  
   reg mem_reg_valid ;  
   reg [31:0] _RAND_22 ;  
   wire killm ;  
   wire _killx_T ;  
   wire killx ;  
   wire _mem_reg_valid_T_1 ;  
   reg [31:0] mem_reg_inst ;  
   reg [31:0] _RAND_23 ;  
   wire wb_reg_valid_x7 ;  
   reg wb_reg_valid ;  
   reg [31:0] _RAND_24 ;  
   reg [1:0] mem_ctrl_typeTagOut ;  
   reg [31:0] _RAND_25 ;  
   reg mem_ctrl_fromint ;  
   reg [31:0] _RAND_26 ;  
   reg mem_ctrl_toint ;  
   reg [31:0] _RAND_27 ;  
   reg mem_ctrl_fastpipe ;  
   reg [31:0] _RAND_28 ;  
   reg mem_ctrl_fma ;  
   reg [31:0] _RAND_29 ;  
   reg mem_ctrl_div ;  
   reg [31:0] _RAND_30 ;  
   reg mem_ctrl_sqrt ;  
   reg [31:0] _RAND_31 ;  
   reg mem_ctrl_wflags ;  
   reg [31:0] _RAND_32 ;  
   reg wb_ctrl_toint ;  
   reg [31:0] _RAND_33 ;  
   wire wdata_truncIdx ;  
   wire [63:0] _wdata_T_1 ;  
   wire [63:0] _wdata_T_2 ;  
   wire wdata_rawIn_sign ;  
   wire [10:0] wdata_rawIn_expIn ;  
   wire [51:0] wdata_rawIn_fractIn ;  
   wire wdata_rawIn_isZeroExpIn ;  
   wire wdata_rawIn_isZeroFractIn ;  
   wire [5:0] _wdata_rawIn_normDist_T_52 ;  
   wire [5:0] _wdata_rawIn_normDist_T_53 ;  
   wire [5:0] _wdata_rawIn_normDist_T_54 ;  
   wire [5:0] _wdata_rawIn_normDist_T_55 ;  
   wire [5:0] _wdata_rawIn_normDist_T_56 ;  
   wire [5:0] _wdata_rawIn_normDist_T_57 ;  
   wire [5:0] _wdata_rawIn_normDist_T_58 ;  
   wire [5:0] _wdata_rawIn_normDist_T_59 ;  
   wire [5:0] _wdata_rawIn_normDist_T_60 ;  
   wire [5:0] _wdata_rawIn_normDist_T_61 ;  
   wire [5:0] _wdata_rawIn_normDist_T_62 ;  
   wire [5:0] _wdata_rawIn_normDist_T_63 ;  
   wire [5:0] _wdata_rawIn_normDist_T_64 ;  
   wire [5:0] _wdata_rawIn_normDist_T_65 ;  
   wire [5:0] _wdata_rawIn_normDist_T_66 ;  
   wire [5:0] _wdata_rawIn_normDist_T_67 ;  
   wire [5:0] _wdata_rawIn_normDist_T_68 ;  
   wire [5:0] _wdata_rawIn_normDist_T_69 ;  
   wire [5:0] _wdata_rawIn_normDist_T_70 ;  
   wire [5:0] _wdata_rawIn_normDist_T_71 ;  
   wire [5:0] _wdata_rawIn_normDist_T_72 ;  
   wire [5:0] _wdata_rawIn_normDist_T_73 ;  
   wire [5:0] _wdata_rawIn_normDist_T_74 ;  
   wire [5:0] _wdata_rawIn_normDist_T_75 ;  
   wire [5:0] _wdata_rawIn_normDist_T_76 ;  
   wire [5:0] _wdata_rawIn_normDist_T_77 ;  
   wire [5:0] _wdata_rawIn_normDist_T_78 ;  
   wire [5:0] _wdata_rawIn_normDist_T_79 ;  
   wire [5:0] _wdata_rawIn_normDist_T_80 ;  
   wire [5:0] _wdata_rawIn_normDist_T_81 ;  
   wire [5:0] _wdata_rawIn_normDist_T_82 ;  
   wire [5:0] _wdata_rawIn_normDist_T_83 ;  
   wire [5:0] _wdata_rawIn_normDist_T_84 ;  
   wire [5:0] _wdata_rawIn_normDist_T_85 ;  
   wire [5:0] _wdata_rawIn_normDist_T_86 ;  
   wire [5:0] _wdata_rawIn_normDist_T_87 ;  
   wire [5:0] _wdata_rawIn_normDist_T_88 ;  
   wire [5:0] _wdata_rawIn_normDist_T_89 ;  
   wire [5:0] _wdata_rawIn_normDist_T_90 ;  
   wire [5:0] _wdata_rawIn_normDist_T_91 ;  
   wire [5:0] _wdata_rawIn_normDist_T_92 ;  
   wire [5:0] _wdata_rawIn_normDist_T_93 ;  
   wire [5:0] _wdata_rawIn_normDist_T_94 ;  
   wire [5:0] _wdata_rawIn_normDist_T_95 ;  
   wire [5:0] _wdata_rawIn_normDist_T_96 ;  
   wire [5:0] _wdata_rawIn_normDist_T_97 ;  
   wire [5:0] _wdata_rawIn_normDist_T_98 ;  
   wire [5:0] _wdata_rawIn_normDist_T_99 ;  
   wire [5:0] _wdata_rawIn_normDist_T_100 ;  
   wire [5:0] _wdata_rawIn_normDist_T_101 ;  
   wire [5:0] wdata_rawIn_normDist ;  
   wire [114:0] _GEN_168 ;  
   wire [114:0] _wdata_rawIn_subnormFract_T ;  
   wire [51:0] wdata_rawIn_subnormFract ;  
   wire [11:0] _GEN_169 ;  
   wire [11:0] _wdata_rawIn_adjustedExp_T ;  
   wire [11:0] _wdata_rawIn_adjustedExp_T_1 ;  
   wire [1:0] _wdata_rawIn_adjustedExp_T_2 ;  
   wire [10:0] _GEN_170 ;  
   wire [10:0] _wdata_rawIn_adjustedExp_T_3 ;  
   wire [11:0] _GEN_171 ;  
   wire [11:0] wdata_rawIn_adjustedExp ;  
   wire wdata_rawIn_isZero ;  
   wire wdata_rawIn_isSpecial ;  
   wire wdata_rawIn__isNaN ;  
   wire [12:0] wdata_rawIn__sExp ;  
   wire wdata_rawIn_out_sig_hi_lo ;  
   wire [51:0] wdata_rawIn_out_sig_lo ;  
   wire [53:0] wdata_rawIn__sig ;  
   wire [2:0] _wdata_T_4 ;  
   wire [2:0] _GEN_172 ;  
   wire [2:0] wdata_hi_lo ;  
   wire [8:0] wdata_lo_hi ;  
   wire [51:0] wdata_lo_lo ;  
   wire [64:0] _wdata_T_6 ;  
   wire wdata_rawIn_sign_1 ;  
   wire [7:0] wdata_rawIn_expIn_1 ;  
   wire [22:0] wdata_rawIn_fractIn_1 ;  
   wire wdata_rawIn_isZeroExpIn_1 ;  
   wire wdata_rawIn_isZeroFractIn_1 ;  
   wire [4:0] _wdata_rawIn_normDist_T_125 ;  
   wire [4:0] _wdata_rawIn_normDist_T_126 ;  
   wire [4:0] _wdata_rawIn_normDist_T_127 ;  
   wire [4:0] _wdata_rawIn_normDist_T_128 ;  
   wire [4:0] _wdata_rawIn_normDist_T_129 ;  
   wire [4:0] _wdata_rawIn_normDist_T_130 ;  
   wire [4:0] _wdata_rawIn_normDist_T_131 ;  
   wire [4:0] _wdata_rawIn_normDist_T_132 ;  
   wire [4:0] _wdata_rawIn_normDist_T_133 ;  
   wire [4:0] _wdata_rawIn_normDist_T_134 ;  
   wire [4:0] _wdata_rawIn_normDist_T_135 ;  
   wire [4:0] _wdata_rawIn_normDist_T_136 ;  
   wire [4:0] _wdata_rawIn_normDist_T_137 ;  
   wire [4:0] _wdata_rawIn_normDist_T_138 ;  
   wire [4:0] _wdata_rawIn_normDist_T_139 ;  
   wire [4:0] _wdata_rawIn_normDist_T_140 ;  
   wire [4:0] _wdata_rawIn_normDist_T_141 ;  
   wire [4:0] _wdata_rawIn_normDist_T_142 ;  
   wire [4:0] _wdata_rawIn_normDist_T_143 ;  
   wire [4:0] _wdata_rawIn_normDist_T_144 ;  
   wire [4:0] _wdata_rawIn_normDist_T_145 ;  
   wire [4:0] wdata_rawIn_normDist_1 ;  
   wire [53:0] _GEN_173 ;  
   wire [53:0] _wdata_rawIn_subnormFract_T_2 ;  
   wire [22:0] wdata_rawIn_subnormFract_1 ;  
   wire [8:0] _GEN_174 ;  
   wire [8:0] _wdata_rawIn_adjustedExp_T_5 ;  
   wire [8:0] _wdata_rawIn_adjustedExp_T_6 ;  
   wire [1:0] _wdata_rawIn_adjustedExp_T_7 ;  
   wire [7:0] _GEN_175 ;  
   wire [7:0] _wdata_rawIn_adjustedExp_T_8 ;  
   wire [8:0] _GEN_176 ;  
   wire [8:0] wdata_rawIn_adjustedExp_1 ;  
   wire wdata_rawIn_isZero_1 ;  
   wire wdata_rawIn_isSpecial_1 ;  
   wire wdata_rawIn_1_isNaN ;  
   wire [9:0] wdata_rawIn_1_sExp ;  
   wire wdata_rawIn_out_sig_hi_lo_1 ;  
   wire [22:0] wdata_rawIn_out_sig_lo_1 ;  
   wire [24:0] wdata_rawIn_1_sig ;  
   wire [2:0] _wdata_T_8 ;  
   wire [2:0] _GEN_177 ;  
   wire [2:0] wdata_hi_lo_1 ;  
   wire [5:0] wdata_lo_hi_1 ;  
   wire [22:0] wdata_lo_lo_1 ;  
   wire [32:0] _wdata_T_10 ;  
   wire [3:0] wdata_swizzledNaN_hi_hi_hi ;  
   wire wdata_swizzledNaN_hi_hi_lo ;  
   wire [6:0] wdata_swizzledNaN_hi_lo_hi ;  
   wire wdata_swizzledNaN_hi_lo_lo ;  
   wire wdata_swizzledNaN_lo_hi_lo ;  
   wire [30:0] wdata_swizzledNaN_lo_lo ;  
   wire [64:0] wdata_swizzledNaN ;  
   wire _wdata_T_12 ;  
   wire [64:0] wdata ;  
   wire _curOK_T_1 ;  
   wire _curOK_T_5 ;  
   wire _curOK_T_6 ;  
   wire curOK ;  
   wire _T_2 ;  
   wire [5:0] _GEN_178 ;  
   wire [5:0] _T_5 ;  
   wire _T_11 ;  
   wire _ex_rm_T_1 ;  
   wire _sfma_io_in_valid_T ;  
   wire _sfma_io_in_valid_T_1 ;  
   wire sfma_io_in_bits_req_in1_unswizzled_hi_hi ;  
   wire sfma_io_in_bits_req_in1_unswizzled_hi_lo ;  
   wire [30:0] sfma_io_in_bits_req_in1_unswizzled_lo ;  
   wire [32:0] sfma_io_in_bits_req_in1_floats_0 ;  
   wire sfma_io_in_bits_req_in1_isbox ;  
   wire [32:0] _sfma_io_in_bits_req_in1_T ;  
   wire [32:0] _sfma_io_in_bits_req_in1_T_1 ;  
   wire sfma_io_in_bits_req_in2_unswizzled_hi_hi ;  
   wire sfma_io_in_bits_req_in2_unswizzled_hi_lo ;  
   wire [30:0] sfma_io_in_bits_req_in2_unswizzled_lo ;  
   wire [32:0] sfma_io_in_bits_req_in2_floats_0 ;  
   wire sfma_io_in_bits_req_in2_isbox ;  
   wire [32:0] _sfma_io_in_bits_req_in2_T ;  
   wire [32:0] _sfma_io_in_bits_req_in2_T_1 ;  
   wire sfma_io_in_bits_req_in3_unswizzled_hi_hi ;  
   wire sfma_io_in_bits_req_in3_unswizzled_hi_lo ;  
   wire [30:0] sfma_io_in_bits_req_in3_unswizzled_lo ;  
   wire [32:0] sfma_io_in_bits_req_in3_floats_0 ;  
   wire sfma_io_in_bits_req_in3_isbox ;  
   wire [32:0] _sfma_io_in_bits_req_in3_T ;  
   wire [32:0] _sfma_io_in_bits_req_in3_T_1 ;  
   wire _sfma_io_in_bits_req_fmaCmd_T_3 ;  
   wire [1:0] _GEN_179 ;  
   wire _fpiu_io_in_valid_T ;  
   wire _fpiu_io_in_valid_T_1 ;  
   wire _fpiu_io_in_valid_T_2 ;  
   wire _fpiu_io_in_valid_T_3 ;  
   wire fpiu_io_in_bits_req_in1_hi_hi ;  
   wire [22:0] fpiu_io_in_bits_req_in1_fractIn ;  
   wire [8:0] fpiu_io_in_bits_req_in1_expIn ;  
   wire [75:0] _fpiu_io_in_bits_req_in1_fractOut_T ;  
   wire [51:0] fpiu_io_in_bits_req_in1_lo ;  
   wire [2:0] fpiu_io_in_bits_req_in1_expOut_hi ;  
   wire [11:0] _GEN_180 ;  
   wire [11:0] _fpiu_io_in_bits_req_in1_expOut_commonCase_T_1 ;  
   wire [11:0] fpiu_io_in_bits_req_in1_expOut_commonCase ;  
   wire _fpiu_io_in_bits_req_in1_expOut_T ;  
   wire _fpiu_io_in_bits_req_in1_expOut_T_1 ;  
   wire _fpiu_io_in_bits_req_in1_expOut_T_2 ;  
   wire [8:0] fpiu_io_in_bits_req_in1_expOut_lo ;  
   wire [11:0] _fpiu_io_in_bits_req_in1_expOut_T_3 ;  
   wire [11:0] fpiu_io_in_bits_req_in1_hi_lo ;  
   wire [64:0] fpiu_io_in_bits_req_in1_floats_0 ;  
   wire fpiu_io_in_bits_req_in1_truncIdx ;  
   wire _fpiu_io_in_bits_req_in1_T_1 ;  
   wire [64:0] _fpiu_io_in_bits_req_in1_T_3 ;  
   wire fpiu_io_in_bits_req_in2_hi_hi ;  
   wire [22:0] fpiu_io_in_bits_req_in2_fractIn ;  
   wire [8:0] fpiu_io_in_bits_req_in2_expIn ;  
   wire [75:0] _fpiu_io_in_bits_req_in2_fractOut_T ;  
   wire [51:0] fpiu_io_in_bits_req_in2_lo ;  
   wire [2:0] fpiu_io_in_bits_req_in2_expOut_hi ;  
   wire [11:0] _GEN_181 ;  
   wire [11:0] _fpiu_io_in_bits_req_in2_expOut_commonCase_T_1 ;  
   wire [11:0] fpiu_io_in_bits_req_in2_expOut_commonCase ;  
   wire _fpiu_io_in_bits_req_in2_expOut_T ;  
   wire _fpiu_io_in_bits_req_in2_expOut_T_1 ;  
   wire _fpiu_io_in_bits_req_in2_expOut_T_2 ;  
   wire [8:0] fpiu_io_in_bits_req_in2_expOut_lo ;  
   wire [11:0] _fpiu_io_in_bits_req_in2_expOut_T_3 ;  
   wire [11:0] fpiu_io_in_bits_req_in2_hi_lo ;  
   wire [64:0] fpiu_io_in_bits_req_in2_floats_0 ;  
   wire _fpiu_io_in_bits_req_in2_T_1 ;  
   wire [64:0] _fpiu_io_in_bits_req_in2_T_3 ;  
   wire [64:0] _ifpu_io_in_bits_in1_T ;  
   reg [4:0] divSqrt_waddr ;  
   reg [31:0] _RAND_34 ;  
   wire _dfma_io_in_valid_T_1 ;  
   wire _memLatencyMask_T_2 ;  
   wire _memLatencyMask_T_3 ;  
   wire [1:0] _memLatencyMask_T_4 ;  
   wire _memLatencyMask_T_5 ;  
   wire _memLatencyMask_T_6 ;  
   wire [2:0] _memLatencyMask_T_7 ;  
   wire _memLatencyMask_T_8 ;  
   wire [1:0] _GEN_188 ;  
   wire [1:0] _memLatencyMask_T_9 ;  
   wire [2:0] _GEN_189 ;  
   wire [2:0] memLatencyMask ;  
   reg [2:0] wen ;  
   reg [31:0] _RAND_35 ;  
   reg [4:0] wbInfo_0_rd ;  
   reg [31:0] _RAND_36 ;  
   reg wbInfo_0_typeTag ;  
   reg [31:0] _RAND_37 ;  
   reg [1:0] wbInfo_0_pipeid ;  
   reg [31:0] _RAND_38 ;  
   reg [4:0] wbInfo_1_rd ;  
   reg [31:0] _RAND_39 ;  
   reg wbInfo_1_typeTag ;  
   reg [31:0] _RAND_40 ;  
   reg [1:0] wbInfo_1_pipeid ;  
   reg [31:0] _RAND_41 ;  
   reg [4:0] wbInfo_2_rd ;  
   reg [31:0] _RAND_42 ;  
   reg wbInfo_2_typeTag ;  
   reg [31:0] _RAND_43 ;  
   reg [1:0] wbInfo_2_pipeid ;  
   reg [31:0] _RAND_44 ;  
   wire _mem_wen_T ;  
   wire _mem_wen_T_1 ;  
   wire mem_wen ;  
   wire [1:0] _write_port_busy_T ;  
   wire [1:0] _write_port_busy_T_1 ;  
   wire _write_port_busy_T_3 ;  
   wire [2:0] _write_port_busy_T_4 ;  
   wire _write_port_busy_T_6 ;  
   wire [3:0] _write_port_busy_T_7 ;  
   wire [1:0] _write_port_busy_T_8 ;  
   wire [2:0] _GEN_190 ;  
   wire [2:0] _write_port_busy_T_9 ;  
   wire [3:0] _GEN_191 ;  
   wire [3:0] _write_port_busy_T_10 ;  
   wire [3:0] _GEN_192 ;  
   wire [3:0] _write_port_busy_T_11 ;  
   wire _write_port_busy_T_12 ;  
   wire _write_port_busy_T_13 ;  
   wire [2:0] _write_port_busy_T_14 ;  
   wire [2:0] _write_port_busy_T_15 ;  
   wire [3:0] _write_port_busy_T_18 ;  
   wire [4:0] _write_port_busy_T_21 ;  
   wire [2:0] _write_port_busy_T_22 ;  
   wire [3:0] _GEN_193 ;  
   wire [3:0] _write_port_busy_T_23 ;  
   wire [4:0] _GEN_194 ;  
   wire [4:0] _write_port_busy_T_24 ;  
   wire [4:0] _GEN_195 ;  
   wire [4:0] _write_port_busy_T_25 ;  
   wire _write_port_busy_T_26 ;  
   wire _write_port_busy_T_27 ;  
   reg write_port_busy ;  
   reg [31:0] _RAND_45 ;  
   wire _GEN_114 ;  
   wire _GEN_118 ;  
   wire [2:0] _GEN_196 ;  
   wire [2:0] _wen_T_2 ;  
   wire _T_20 ;  
   wire [1:0] _wbInfo_0_pipeid_T_7 ;  
   wire [1:0] _GEN_197 ;  
   wire [1:0] _wbInfo_0_pipeid_T_9 ;  
   wire [1:0] _wbInfo_0_pipeid_T_10 ;  
   wire [1:0] _GEN_123 ;  
   wire _T_23 ;  
   wire [1:0] _GEN_127 ;  
   wire _T_26 ;  
   wire [1:0] _GEN_131 ;  
   wire [1:0] _GEN_136 ;  
   wire [1:0] _GEN_140 ;  
   wire [1:0] _GEN_144 ;  
   wire divSqrt_typeTag ;  
   reg divSqrt_killed ;  
   reg [31:0] _RAND_46 ;  
   wire _T_52 ;  
   wire _GEN_158 ;  
   wire divSqrt_wen ;  
   wire [4:0] waddr ;  
   wire wtypeTag ;  
   wire _wdata_T_13 ;  
   wire [64:0] _wdata_T_14 ;  
   wire _wdata_T_15 ;  
   wire [64:0] _wdata_T_16 ;  
   wire _wdata_T_17 ;  
   wire [64:0] _wdata_T_18 ;  
   wire _divSqrt_wdata_T_1 ;  
   wire [64:0] divSqrt_wdata_maskedNaN ;  
   wire [64:0] _divSqrt_wdata_T_2 ;  
   wire [32:0] _GEN_159 ;  
   wire [64:0] divSqrt_wdata ;  
   wire [64:0] _wdata_T_19 ;  
   wire wdata_opts_bigger_swizzledNaN_hi_hi_lo ;  
   wire wdata_opts_bigger_swizzledNaN_hi_lo_lo ;  
   wire wdata_opts_bigger_swizzledNaN_lo_hi_lo ;  
   wire [30:0] wdata_opts_bigger_swizzledNaN_lo_lo ;  
   wire [64:0] wdata_opts_bigger_swizzledNaN ;  
   wire _wdata_opts_bigger_T ;  
   wire [64:0] wdata_opts_bigger ;  
   wire [64:0] wdata_1 ;  
   wire [4:0] _wexc_T_1 ;  
   wire [4:0] _wexc_T_3 ;  
   wire [4:0] wexc ;  
   wire frfWriteBundle_1_wrenf ;  
   wire unswizzled_hi_hi_1 ;  
   wire unswizzled_hi_lo_1 ;  
   wire [30:0] unswizzled_lo_1 ;  
   wire [32:0] unswizzled_1 ;  
   wire _curOK_T_8 ;  
   wire _curOK_T_12 ;  
   wire _curOK_T_13 ;  
   wire curOK_1 ;  
   wire _T_33 ;  
   wire [5:0] _GEN_200 ;  
   wire [5:0] _T_36 ;  
   wire [11:0] unrecoded_rawIn_exp ;  
   wire unrecoded_rawIn_isZero ;  
   wire unrecoded_rawIn_isSpecial ;  
   wire unrecoded_rawIn__isNaN ;  
   wire unrecoded_rawIn__isInf ;  
   wire unrecoded_rawIn__sign ;  
   wire [12:0] unrecoded_rawIn__sExp ;  
   wire unrecoded_rawIn_out_sig_hi_lo ;  
   wire [51:0] unrecoded_rawIn_out_sig_lo ;  
   wire [53:0] unrecoded_rawIn__sig ;  
   wire unrecoded_isSubnormal ;  
   wire [5:0] unrecoded_denormShiftDist ;  
   wire [52:0] _unrecoded_denormFract_T_1 ;  
   wire [51:0] unrecoded_denormFract ;  
   wire [10:0] _unrecoded_expOut_T_2 ;  
   wire [10:0] _unrecoded_expOut_T_3 ;  
   wire _unrecoded_expOut_T_4 ;  
   wire [10:0] _unrecoded_expOut_T_6 ;  
   wire [10:0] unrecoded_hi_lo ;  
   wire [51:0] _unrecoded_fractOut_T_1 ;  
   wire [51:0] unrecoded_lo ;  
   wire [63:0] unrecoded ;  
   wire [8:0] prevUnrecoded_rawIn_exp ;  
   wire prevUnrecoded_rawIn_isZero ;  
   wire prevUnrecoded_rawIn_isSpecial ;  
   wire prevUnrecoded_rawIn__isNaN ;  
   wire prevUnrecoded_rawIn__isInf ;  
   wire prevUnrecoded_rawIn__sign ;  
   wire [9:0] prevUnrecoded_rawIn__sExp ;  
   wire prevUnrecoded_rawIn_out_sig_hi_lo ;  
   wire [22:0] prevUnrecoded_rawIn_out_sig_lo ;  
   wire [24:0] prevUnrecoded_rawIn__sig ;  
   wire prevUnrecoded_isSubnormal ;  
   wire [4:0] prevUnrecoded_denormShiftDist ;  
   wire [23:0] _prevUnrecoded_denormFract_T_1 ;  
   wire [22:0] prevUnrecoded_denormFract ;  
   wire [7:0] _prevUnrecoded_expOut_T_2 ;  
   wire [7:0] _prevUnrecoded_expOut_T_3 ;  
   wire _prevUnrecoded_expOut_T_4 ;  
   wire [7:0] _prevUnrecoded_expOut_T_6 ;  
   wire [7:0] prevUnrecoded_hi_lo ;  
   wire [22:0] _prevUnrecoded_fractOut_T_1 ;  
   wire [22:0] prevUnrecoded_lo ;  
   wire [31:0] prevUnrecoded ;  
   wire [31:0] hi ;  
   wire [31:0] lo ;  
   wire [63:0] _T_40 ;  
   wire wb_toint_valid ;  
   reg [4:0] wb_toint_exc ;  
   reg [31:0] _RAND_47 ;  
   wire _io_fcsr_flags_valid_T ;  
   wire [4:0] _io_fcsr_flags_bits_T ;  
   wire [4:0] _GEN_160 ;  
   wire [4:0] divSqrt_flags ;  
   wire [4:0] _io_fcsr_flags_bits_T_1 ;  
   wire [4:0] _io_fcsr_flags_bits_T_2 ;  
   wire [4:0] _io_fcsr_flags_bits_T_4 ;  
   wire _divSqrt_write_port_busy_T ;  
   wire _divSqrt_write_port_busy_T_1 ;  
   wire divSqrt_write_port_busy ;  
   wire _io_fcsr_rdy_T ;  
   wire _io_fcsr_rdy_T_1 ;  
   wire _io_fcsr_rdy_T_2 ;  
   wire _io_fcsr_rdy_T_4 ;  
   wire _io_fcsr_rdy_T_6 ;  
   wire _GEN_162 ;  
   wire divSqrt_inFlight ;  
   wire _io_fcsr_rdy_T_7 ;  
   wire _io_nack_mem_T ;  
   wire _io_sboard_set_x27_T_3 ;  
   reg io_sboard_set_REG ;  
   reg [31:0] _RAND_48 ;  
   wire _io_sboard_clr_T_4 ;  
   wire _io_illegal_rm_T_1 ;  
   wire _io_illegal_rm_T_2 ;  
   wire _io_illegal_rm_T_3 ;  
   wire _io_illegal_rm_T_5 ;  
   wire _io_illegal_rm_T_6 ;  
   wire _io_illegal_rm_T_7 ;  
   wire _divSqrt_inValid_T_1 ;  
   wire divSqrt_inValid ;  
   wire _divSqrt_killed_T ;  
   wire divSqrt_io_a_hi_hi ;  
   wire [51:0] divSqrt_io_a_fractIn ;  
   wire [11:0] divSqrt_io_a_expIn ;  
   wire [75:0] _divSqrt_io_a_fractOut_T ;  
   wire [22:0] divSqrt_io_a_lo ;  
   wire [2:0] divSqrt_io_a_expOut_hi ;  
   wire [11:0] _divSqrt_io_a_expOut_commonCase_T_1 ;  
   wire [11:0] divSqrt_io_a_expOut_commonCase ;  
   wire _divSqrt_io_a_expOut_T ;  
   wire _divSqrt_io_a_expOut_T_1 ;  
   wire _divSqrt_io_a_expOut_T_2 ;  
   wire [5:0] divSqrt_io_a_expOut_lo ;  
   wire [8:0] _divSqrt_io_a_expOut_T_3 ;  
   wire [8:0] divSqrt_io_a_hi_lo ;  
   wire [9:0] divSqrt_io_a_hi ;  
   wire divSqrt_io_b_hi_hi ;  
   wire [51:0] divSqrt_io_b_fractIn ;  
   wire [11:0] divSqrt_io_b_expIn ;  
   wire [75:0] _divSqrt_io_b_fractOut_T ;  
   wire [22:0] divSqrt_io_b_lo ;  
   wire [2:0] divSqrt_io_b_expOut_hi ;  
   wire [11:0] _divSqrt_io_b_expOut_commonCase_T_1 ;  
   wire [11:0] divSqrt_io_b_expOut_commonCase ;  
   wire _divSqrt_io_b_expOut_T ;  
   wire _divSqrt_io_b_expOut_T_1 ;  
   wire _divSqrt_io_b_expOut_T_2 ;  
   wire [5:0] divSqrt_io_b_expOut_lo ;  
   wire [8:0] _divSqrt_io_b_expOut_T_3 ;  
   wire [8:0] divSqrt_io_b_hi_lo ;  
   wire [9:0] divSqrt_io_b_hi ;  
   reg [19:0] FPU_state ;  
   reg [31:0] _RAND_49 ;  
   reg FPU_cov[0:1048575] ;  
   reg [31:0] _RAND_50 ;  
   wire FPU_cov_read_data ;  
   wire [19:0] FPU_cov_read_addr ;  
   wire FPU_cov_write_data ;  
   wire [19:0] FPU_cov_write_addr ;  
   wire FPU_cov_write_mask ;  
   wire FPU_cov_write_en ;  
   reg [29:0] FPU_covSum ;  
   reg [31:0] _RAND_51 ;  
   wire [16:0] wbInfo_0_typeTag_shl ;  
   wire [19:0] wbInfo_0_typeTag_pad ;  
   wire [2:0] wb_reg_valid_shl ;  
   wire [19:0] wb_reg_valid_pad ;  
   wire [7:0] mem_ctrl_sqrt_shl ;  
   wire [19:0] mem_ctrl_sqrt_pad ;  
   wire [19:0] divSqrt_killed_shl ;  
   wire [19:0] divSqrt_killed_pad ;  
   wire [8:0] ex_reg_ctrl_typeTagIn_shl ;  
   wire [19:0] ex_reg_ctrl_typeTagIn_pad ;  
   wire [2:0] ex_reg_ctrl_fromint_shl ;  
   wire [19:0] ex_reg_ctrl_fromint_pad ;  
   wire [8:0] mem_ctrl_typeTagOut_shl ;  
   wire [19:0] mem_ctrl_typeTagOut_pad ;  
   wire [7:0] wen_shl ;  
   wire [19:0] wen_pad ;  
   wire [11:0] wb_ctrl_toint_shl ;  
   wire [19:0] wb_ctrl_toint_pad ;  
   wire [18:0] ex_reg_ctrl_fastpipe_shl ;  
   wire [19:0] ex_reg_ctrl_fastpipe_pad ;  
   wire [14:0] write_port_busy_shl ;  
   wire [19:0] write_port_busy_pad ;  
   wire [5:0] mem_ctrl_fastpipe_shl ;  
   wire [19:0] mem_ctrl_fastpipe_pad ;  
   wire [14:0] ex_reg_ctrl_typeTagOut_shl ;  
   wire [19:0] ex_reg_ctrl_typeTagOut_pad ;  
   wire [17:0] mem_reg_valid_shl ;  
   wire [19:0] mem_reg_valid_pad ;  
   wire [13:0] mem_ctrl_div_shl ;  
   wire [19:0] mem_ctrl_div_pad ;  
   wire [11:0] wbInfo_0_pipeid_shl ;  
   wire [19:0] wbInfo_0_pipeid_pad ;  
   wire [1:0] mem_ctrl_toint_shl ;  
   wire [19:0] mem_ctrl_toint_pad ;  
   wire [4:0] ex_reg_ctrl_fma_shl ;  
   wire [19:0] ex_reg_ctrl_fma_pad ;  
   wire [3:0] ex_reg_valid_shl ;  
   wire [19:0] ex_reg_valid_pad ;  
   wire [10:0] mem_ctrl_fromint_shl ;  
   wire [19:0] mem_ctrl_fromint_pad ;  
   wire [2:0] mem_ctrl_fma_shl ;  
   wire [19:0] mem_ctrl_fma_pad ;  
   wire [19:0] FPU_xor7 ;  
   wire [19:0] FPU_xor18 ;  
   wire [19:0] FPU_xor8 ;  
   wire [19:0] FPU_xor3 ;  
   wire [19:0] FPU_xor9 ;  
   wire [19:0] FPU_xor22 ;  
   wire [19:0] FPU_xor10 ;  
   wire [19:0] FPU_xor4 ;  
   wire [19:0] FPU_xor1 ;  
   wire [19:0] FPU_xor11 ;  
   wire [19:0] FPU_xor26 ;  
   wire [19:0] FPU_xor12 ;  
   wire [19:0] FPU_xor5 ;  
   wire [19:0] FPU_xor28 ;  
   wire [19:0] FPU_xor13 ;  
   wire [19:0] FPU_xor30 ;  
   wire [19:0] FPU_xor14 ;  
   wire [19:0] FPU_xor6 ;  
   wire [19:0] FPU_xor2 ;  
   wire [19:0] FPU_xor0 ;  
   wire [29:0] fpiu_sum ;  
   wire [29:0] fp_decoder_sum ;  
   wire [29:0] ifpu_sum ;  
   wire [29:0] sfma_sum ;  
   wire [29:0] fpmu_sum ;  
   wire [29:0] divSqrt_1_sum ;  
   wire [29:0] dfma_sum ;  
   wire [29:0] divSqrt_sum ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire ifpu_metaAssert_wire ;  
   wire fpmu_metaAssert_wire ;  
   wire fp_decoder_metaAssert_wire ;  
   wire fpiu_metaAssert_wire ;  
   wire divSqrt_1_metaAssert_wire ;  
   wire divSqrt_metaAssert_wire ;  
   wire dfma_metaAssert_wire ;  
   wire sfma_metaAssert_wire ;  
   wire FPU_or3 ;  
   wire FPU_or10 ;  
   wire FPU_or4 ;  
   wire FPU_or1 ;  
   wire FPU_or5 ;  
   wire FPU_or14 ;  
   wire FPU_or6 ;  
   wire FPU_or2 ;  
   wire FPU_or0 ;  
   reg FPU_metaAssert ;  
   reg [31:0] _RAND_52 ;  
  FPUDecoder fp_decoder(.io_inst(fp_decoder_io_inst),.io_sigs_wen(fp_decoder_io_sigs_wen),.io_sigs_ren1(fp_decoder_io_sigs_ren1),.io_sigs_ren2(fp_decoder_io_sigs_ren2),.io_sigs_ren3(fp_decoder_io_sigs_ren3),.io_sigs_swap12(fp_decoder_io_sigs_swap12),.io_sigs_swap23(fp_decoder_io_sigs_swap23),.io_sigs_typeTagIn(fp_decoder_io_sigs_typeTagIn),.io_sigs_typeTagOut(fp_decoder_io_sigs_typeTagOut),.io_sigs_fromint(fp_decoder_io_sigs_fromint),.io_sigs_toint(fp_decoder_io_sigs_toint),.io_sigs_fastpipe(fp_decoder_io_sigs_fastpipe),.io_sigs_fma(fp_decoder_io_sigs_fma),.io_sigs_div(fp_decoder_io_sigs_div),.io_sigs_sqrt(fp_decoder_io_sigs_sqrt),.io_sigs_wflags(fp_decoder_io_sigs_wflags),.io_covSum(fp_decoder_io_covSum),.metaAssert(fp_decoder_metaAssert)); 
  FPUFMAPipe sfma(.clock(sfma_clock),.reset(sfma_reset),.io_in_valid(sfma_io_in_valid),.io_in_bits_ren3(sfma_io_in_bits_ren3),.io_in_bits_swap23(sfma_io_in_bits_swap23),.io_in_bits_rm(sfma_io_in_bits_rm),.io_in_bits_fmaCmd(sfma_io_in_bits_fmaCmd),.io_in_bits_in1(sfma_io_in_bits_in1),.io_in_bits_in2(sfma_io_in_bits_in2),.io_in_bits_in3(sfma_io_in_bits_in3),.io_out_bits_data(sfma_io_out_bits_data),.io_out_bits_exc(sfma_io_out_bits_exc),.io_covSum(sfma_io_covSum),.metaAssert(sfma_metaAssert),.metaReset(sfma_metaReset),.fma_halt(sfma_fma_halt)); 
  FPToInt fpiu(.clock(fpiu_clock),.io_in_valid(fpiu_io_in_valid),.io_in_bits_ren2(fpiu_io_in_bits_ren2),.io_in_bits_typeTagIn(fpiu_io_in_bits_typeTagIn),.io_in_bits_typeTagOut(fpiu_io_in_bits_typeTagOut),.io_in_bits_wflags(fpiu_io_in_bits_wflags),.io_in_bits_rm(fpiu_io_in_bits_rm),.io_in_bits_typ(fpiu_io_in_bits_typ),.io_in_bits_fmt(fpiu_io_in_bits_fmt),.io_in_bits_in1(fpiu_io_in_bits_in1),.io_in_bits_in2(fpiu_io_in_bits_in2),.io_out_bits_in_rm(fpiu_io_out_bits_in_rm),.io_out_bits_in_in1(fpiu_io_out_bits_in_in1),.io_out_bits_in_in2(fpiu_io_out_bits_in_in2),.io_out_bits_lt(fpiu_io_out_bits_lt),.io_out_bits_store(fpiu_io_out_bits_store),.io_out_bits_toint(fpiu_io_out_bits_toint),.io_out_bits_exc(fpiu_io_out_bits_exc),.io_covSum(fpiu_io_covSum),.metaAssert(fpiu_metaAssert),.metaReset(fpiu_metaReset)); 
  IntToFP ifpu(.clock(ifpu_clock),.reset(ifpu_reset),.io_in_valid(ifpu_io_in_valid),.io_in_bits_typeTagIn(ifpu_io_in_bits_typeTagIn),.io_in_bits_wflags(ifpu_io_in_bits_wflags),.io_in_bits_rm(ifpu_io_in_bits_rm),.io_in_bits_typ(ifpu_io_in_bits_typ),.io_in_bits_in1(ifpu_io_in_bits_in1),.io_out_bits_data(ifpu_io_out_bits_data),.io_out_bits_exc(ifpu_io_out_bits_exc),.io_covSum(ifpu_io_covSum),.metaAssert(ifpu_metaAssert),.metaReset(ifpu_metaReset)); 
  FPToFP fpmu(.clock(fpmu_clock),.reset(fpmu_reset),.io_in_valid(fpmu_io_in_valid),.io_in_bits_ren2(fpmu_io_in_bits_ren2),.io_in_bits_typeTagOut(fpmu_io_in_bits_typeTagOut),.io_in_bits_wflags(fpmu_io_in_bits_wflags),.io_in_bits_rm(fpmu_io_in_bits_rm),.io_in_bits_in1(fpmu_io_in_bits_in1),.io_in_bits_in2(fpmu_io_in_bits_in2),.io_out_bits_data(fpmu_io_out_bits_data),.io_out_bits_exc(fpmu_io_out_bits_exc),.io_lt(fpmu_io_lt),.io_covSum(fpmu_io_covSum),.metaAssert(fpmu_metaAssert),.metaReset(fpmu_metaReset)); 
  FPUFMAPipe_1 dfma(.clock(dfma_clock),.reset(dfma_reset),.io_in_valid(dfma_io_in_valid),.io_in_bits_ren3(dfma_io_in_bits_ren3),.io_in_bits_swap23(dfma_io_in_bits_swap23),.io_in_bits_rm(dfma_io_in_bits_rm),.io_in_bits_fmaCmd(dfma_io_in_bits_fmaCmd),.io_in_bits_in1(dfma_io_in_bits_in1),.io_in_bits_in2(dfma_io_in_bits_in2),.io_in_bits_in3(dfma_io_in_bits_in3),.io_out_bits_data(dfma_io_out_bits_data),.io_out_bits_exc(dfma_io_out_bits_exc),.io_covSum(dfma_io_covSum),.metaAssert(dfma_metaAssert),.metaReset(dfma_metaReset),.fma_halt(dfma_fma_halt)); 
  DivSqrtRecFN_small divSqrt(.clock(divSqrt_clock),.reset(divSqrt_reset),.io_inReady(divSqrt_io_inReady),.io_inValid(divSqrt_io_inValid),.io_sqrtOp(divSqrt_io_sqrtOp),.io_a(divSqrt_io_a),.io_b(divSqrt_io_b),.io_roundingMode(divSqrt_io_roundingMode),.io_outValid_div(divSqrt_io_outValid_div),.io_outValid_sqrt(divSqrt_io_outValid_sqrt),.io_out(divSqrt_io_out),.io_exceptionFlags(divSqrt_io_exceptionFlags),.io_covSum(divSqrt_io_covSum),.metaAssert(divSqrt_metaAssert),.metaReset(divSqrt_metaReset),.divSqrtRecFNToRaw_halt(divSqrt_divSqrtRecFNToRaw_halt)); 
  DivSqrtRecFN_small_1 divSqrt_1(.clock(divSqrt_1_clock),.reset(divSqrt_1_reset),.io_inReady(divSqrt_1_io_inReady),.io_inValid(divSqrt_1_io_inValid),.io_sqrtOp(divSqrt_1_io_sqrtOp),.io_a(divSqrt_1_io_a),.io_b(divSqrt_1_io_b),.io_roundingMode(divSqrt_1_io_roundingMode),.io_outValid_div(divSqrt_1_io_outValid_div),.io_outValid_sqrt(divSqrt_1_io_outValid_sqrt),.io_out(divSqrt_1_io_out),.io_exceptionFlags(divSqrt_1_io_exceptionFlags),.io_covSum(divSqrt_1_io_covSum),.metaAssert(divSqrt_1_metaAssert),.metaReset(divSqrt_1_metaReset),.divSqrtRecFNToRaw_halt(divSqrt_1_divSqrtRecFNToRaw_halt)); 
  assign regfile_ex_rs_0_addr=ex_ra_0; 
  assign regfile_ex_rs_0_data=regfile[regfile_ex_rs_0_addr]; 
  assign regfile_ex_rs_1_addr=ex_ra_1; 
  assign regfile_ex_rs_1_data=regfile[regfile_ex_rs_1_addr]; 
  assign regfile_ex_rs_2_addr=ex_ra_2; 
  assign regfile_ex_rs_2_data=regfile[regfile_ex_rs_2_addr]; 
  assign regfile_MPORT_data=_wdata_T_12 ? wdata_swizzledNaN:_wdata_T_6; 
  assign regfile_MPORT_addr=load_wb_tag; 
  assign regfile_MPORT_mask=1'h1; 
  assign regfile_MPORT_en=load_wb; 
  assign regfile_MPORT_1_data=wtypeTag ? _wdata_T_19:wdata_opts_bigger; 
  assign regfile_MPORT_1_addr=divSqrt_wen ? divSqrt_waddr:wbInfo_0_rd; 
  assign regfile_MPORT_1_mask=1'h1; 
  assign regfile_MPORT_1_en=wen[0]|divSqrt_wen; 
  assign _load_wb_typeTag_T_2=io_dmem_resp_type[1:0]-2'h2; 
  assign killm=io_killm|io_nack_mem; 
  assign _killx_T=mem_reg_valid&killm; 
  assign killx=io_killx|_killx_T; 
  assign _mem_reg_valid_T_1=ex_reg_valid&~killx; 
  assign wb_reg_valid_x7=mem_reg_valid&~killm; 
  assign wdata_truncIdx=load_wb_typeTag[0]; 
  assign _wdata_T_1=wdata_truncIdx ? 64'h0:64'hffffffff00000000; 
  assign _wdata_T_2=_wdata_T_1|load_wb_data; 
  assign wdata_rawIn_sign=_wdata_T_2[63]; 
  assign wdata_rawIn_expIn=_wdata_T_2[62:52]; 
  assign wdata_rawIn_fractIn=_wdata_T_2[51:0]; 
  assign wdata_rawIn_isZeroExpIn=wdata_rawIn_expIn==11'h0; 
  assign wdata_rawIn_isZeroFractIn=wdata_rawIn_fractIn==52'h0; 
  assign _wdata_rawIn_normDist_T_52=wdata_rawIn_fractIn[1] ? 6'h32:6'h33; 
  assign _wdata_rawIn_normDist_T_53=wdata_rawIn_fractIn[2] ? 6'h31:_wdata_rawIn_normDist_T_52; 
  assign _wdata_rawIn_normDist_T_54=wdata_rawIn_fractIn[3] ? 6'h30:_wdata_rawIn_normDist_T_53; 
  assign _wdata_rawIn_normDist_T_55=wdata_rawIn_fractIn[4] ? 6'h2f:_wdata_rawIn_normDist_T_54; 
  assign _wdata_rawIn_normDist_T_56=wdata_rawIn_fractIn[5] ? 6'h2e:_wdata_rawIn_normDist_T_55; 
  assign _wdata_rawIn_normDist_T_57=wdata_rawIn_fractIn[6] ? 6'h2d:_wdata_rawIn_normDist_T_56; 
  assign _wdata_rawIn_normDist_T_58=wdata_rawIn_fractIn[7] ? 6'h2c:_wdata_rawIn_normDist_T_57; 
  assign _wdata_rawIn_normDist_T_59=wdata_rawIn_fractIn[8] ? 6'h2b:_wdata_rawIn_normDist_T_58; 
  assign _wdata_rawIn_normDist_T_60=wdata_rawIn_fractIn[9] ? 6'h2a:_wdata_rawIn_normDist_T_59; 
  assign _wdata_rawIn_normDist_T_61=wdata_rawIn_fractIn[10] ? 6'h29:_wdata_rawIn_normDist_T_60; 
  assign _wdata_rawIn_normDist_T_62=wdata_rawIn_fractIn[11] ? 6'h28:_wdata_rawIn_normDist_T_61; 
  assign _wdata_rawIn_normDist_T_63=wdata_rawIn_fractIn[12] ? 6'h27:_wdata_rawIn_normDist_T_62; 
  assign _wdata_rawIn_normDist_T_64=wdata_rawIn_fractIn[13] ? 6'h26:_wdata_rawIn_normDist_T_63; 
  assign _wdata_rawIn_normDist_T_65=wdata_rawIn_fractIn[14] ? 6'h25:_wdata_rawIn_normDist_T_64; 
  assign _wdata_rawIn_normDist_T_66=wdata_rawIn_fractIn[15] ? 6'h24:_wdata_rawIn_normDist_T_65; 
  assign _wdata_rawIn_normDist_T_67=wdata_rawIn_fractIn[16] ? 6'h23:_wdata_rawIn_normDist_T_66; 
  assign _wdata_rawIn_normDist_T_68=wdata_rawIn_fractIn[17] ? 6'h22:_wdata_rawIn_normDist_T_67; 
  assign _wdata_rawIn_normDist_T_69=wdata_rawIn_fractIn[18] ? 6'h21:_wdata_rawIn_normDist_T_68; 
  assign _wdata_rawIn_normDist_T_70=wdata_rawIn_fractIn[19] ? 6'h20:_wdata_rawIn_normDist_T_69; 
  assign _wdata_rawIn_normDist_T_71=wdata_rawIn_fractIn[20] ? 6'h1f:_wdata_rawIn_normDist_T_70; 
  assign _wdata_rawIn_normDist_T_72=wdata_rawIn_fractIn[21] ? 6'h1e:_wdata_rawIn_normDist_T_71; 
  assign _wdata_rawIn_normDist_T_73=wdata_rawIn_fractIn[22] ? 6'h1d:_wdata_rawIn_normDist_T_72; 
  assign _wdata_rawIn_normDist_T_74=wdata_rawIn_fractIn[23] ? 6'h1c:_wdata_rawIn_normDist_T_73; 
  assign _wdata_rawIn_normDist_T_75=wdata_rawIn_fractIn[24] ? 6'h1b:_wdata_rawIn_normDist_T_74; 
  assign _wdata_rawIn_normDist_T_76=wdata_rawIn_fractIn[25] ? 6'h1a:_wdata_rawIn_normDist_T_75; 
  assign _wdata_rawIn_normDist_T_77=wdata_rawIn_fractIn[26] ? 6'h19:_wdata_rawIn_normDist_T_76; 
  assign _wdata_rawIn_normDist_T_78=wdata_rawIn_fractIn[27] ? 6'h18:_wdata_rawIn_normDist_T_77; 
  assign _wdata_rawIn_normDist_T_79=wdata_rawIn_fractIn[28] ? 6'h17:_wdata_rawIn_normDist_T_78; 
  assign _wdata_rawIn_normDist_T_80=wdata_rawIn_fractIn[29] ? 6'h16:_wdata_rawIn_normDist_T_79; 
  assign _wdata_rawIn_normDist_T_81=wdata_rawIn_fractIn[30] ? 6'h15:_wdata_rawIn_normDist_T_80; 
  assign _wdata_rawIn_normDist_T_82=wdata_rawIn_fractIn[31] ? 6'h14:_wdata_rawIn_normDist_T_81; 
  assign _wdata_rawIn_normDist_T_83=wdata_rawIn_fractIn[32] ? 6'h13:_wdata_rawIn_normDist_T_82; 
  assign _wdata_rawIn_normDist_T_84=wdata_rawIn_fractIn[33] ? 6'h12:_wdata_rawIn_normDist_T_83; 
  assign _wdata_rawIn_normDist_T_85=wdata_rawIn_fractIn[34] ? 6'h11:_wdata_rawIn_normDist_T_84; 
  assign _wdata_rawIn_normDist_T_86=wdata_rawIn_fractIn[35] ? 6'h10:_wdata_rawIn_normDist_T_85; 
  assign _wdata_rawIn_normDist_T_87=wdata_rawIn_fractIn[36] ? 6'hf:_wdata_rawIn_normDist_T_86; 
  assign _wdata_rawIn_normDist_T_88=wdata_rawIn_fractIn[37] ? 6'he:_wdata_rawIn_normDist_T_87; 
  assign _wdata_rawIn_normDist_T_89=wdata_rawIn_fractIn[38] ? 6'hd:_wdata_rawIn_normDist_T_88; 
  assign _wdata_rawIn_normDist_T_90=wdata_rawIn_fractIn[39] ? 6'hc:_wdata_rawIn_normDist_T_89; 
  assign _wdata_rawIn_normDist_T_91=wdata_rawIn_fractIn[40] ? 6'hb:_wdata_rawIn_normDist_T_90; 
  assign _wdata_rawIn_normDist_T_92=wdata_rawIn_fractIn[41] ? 6'ha:_wdata_rawIn_normDist_T_91; 
  assign _wdata_rawIn_normDist_T_93=wdata_rawIn_fractIn[42] ? 6'h9:_wdata_rawIn_normDist_T_92; 
  assign _wdata_rawIn_normDist_T_94=wdata_rawIn_fractIn[43] ? 6'h8:_wdata_rawIn_normDist_T_93; 
  assign _wdata_rawIn_normDist_T_95=wdata_rawIn_fractIn[44] ? 6'h7:_wdata_rawIn_normDist_T_94; 
  assign _wdata_rawIn_normDist_T_96=wdata_rawIn_fractIn[45] ? 6'h6:_wdata_rawIn_normDist_T_95; 
  assign _wdata_rawIn_normDist_T_97=wdata_rawIn_fractIn[46] ? 6'h5:_wdata_rawIn_normDist_T_96; 
  assign _wdata_rawIn_normDist_T_98=wdata_rawIn_fractIn[47] ? 6'h4:_wdata_rawIn_normDist_T_97; 
  assign _wdata_rawIn_normDist_T_99=wdata_rawIn_fractIn[48] ? 6'h3:_wdata_rawIn_normDist_T_98; 
  assign _wdata_rawIn_normDist_T_100=wdata_rawIn_fractIn[49] ? 6'h2:_wdata_rawIn_normDist_T_99; 
  assign _wdata_rawIn_normDist_T_101=wdata_rawIn_fractIn[50] ? 6'h1:_wdata_rawIn_normDist_T_100; 
  assign wdata_rawIn_normDist=wdata_rawIn_fractIn[51] ? 6'h0:_wdata_rawIn_normDist_T_101; 
  assign _GEN_168={63'b0,wdata_rawIn_fractIn}; 
  assign _wdata_rawIn_subnormFract_T=_GEN_168<<wdata_rawIn_normDist; 
  assign wdata_rawIn_subnormFract={_wdata_rawIn_subnormFract_T[50:0],1'h0}; 
  assign _GEN_169={6'b0,wdata_rawIn_normDist}; 
  assign _wdata_rawIn_adjustedExp_T=_GEN_169^12'hfff; 
  assign _wdata_rawIn_adjustedExp_T_1=wdata_rawIn_isZeroExpIn ? _wdata_rawIn_adjustedExp_T:{1'b0,wdata_rawIn_expIn}; 
  assign _wdata_rawIn_adjustedExp_T_2=wdata_rawIn_isZeroExpIn ? 2'h2:2'h1; 
  assign _GEN_170={9'b0,_wdata_rawIn_adjustedExp_T_2}; 
  assign _wdata_rawIn_adjustedExp_T_3=11'h400|_GEN_170; 
  assign _GEN_171={1'b0,_wdata_rawIn_adjustedExp_T_3}; 
  assign wdata_rawIn_adjustedExp=_wdata_rawIn_adjustedExp_T_1+_GEN_171; 
  assign wdata_rawIn_isZero=wdata_rawIn_isZeroExpIn&wdata_rawIn_isZeroFractIn; 
  assign wdata_rawIn_isSpecial=wdata_rawIn_adjustedExp[11:10]==2'h3; 
  assign wdata_rawIn__isNaN=wdata_rawIn_isSpecial&~wdata_rawIn_isZeroFractIn; 
  assign wdata_rawIn__sExp={1'b0,$signed(wdata_rawIn_adjustedExp)}; 
  assign wdata_rawIn_out_sig_hi_lo=~wdata_rawIn_isZero; 
  assign wdata_rawIn_out_sig_lo=wdata_rawIn_isZeroExpIn ? wdata_rawIn_subnormFract:wdata_rawIn_fractIn; 
  assign wdata_rawIn__sig={1'h0,wdata_rawIn_out_sig_hi_lo,wdata_rawIn_out_sig_lo}; 
  assign _wdata_T_4=wdata_rawIn_isZero ? 3'h0:wdata_rawIn__sExp[11:9]; 
  assign _GEN_172={2'b0,wdata_rawIn__isNaN}; 
  assign wdata_hi_lo=_wdata_T_4|_GEN_172; 
  assign wdata_lo_hi=wdata_rawIn__sExp[8:0]; 
  assign wdata_lo_lo=wdata_rawIn__sig[51:0]; 
  assign _wdata_T_6={wdata_rawIn_sign,wdata_hi_lo,wdata_lo_hi,wdata_lo_lo}; 
  assign wdata_rawIn_sign_1=_wdata_T_2[31]; 
  assign wdata_rawIn_expIn_1=_wdata_T_2[30:23]; 
  assign wdata_rawIn_fractIn_1=_wdata_T_2[22:0]; 
  assign wdata_rawIn_isZeroExpIn_1=wdata_rawIn_expIn_1==8'h0; 
  assign wdata_rawIn_isZeroFractIn_1=wdata_rawIn_fractIn_1==23'h0; 
  assign _wdata_rawIn_normDist_T_125=wdata_rawIn_fractIn_1[1] ? 5'h15:5'h16; 
  assign _wdata_rawIn_normDist_T_126=wdata_rawIn_fractIn_1[2] ? 5'h14:_wdata_rawIn_normDist_T_125; 
  assign _wdata_rawIn_normDist_T_127=wdata_rawIn_fractIn_1[3] ? 5'h13:_wdata_rawIn_normDist_T_126; 
  assign _wdata_rawIn_normDist_T_128=wdata_rawIn_fractIn_1[4] ? 5'h12:_wdata_rawIn_normDist_T_127; 
  assign _wdata_rawIn_normDist_T_129=wdata_rawIn_fractIn_1[5] ? 5'h11:_wdata_rawIn_normDist_T_128; 
  assign _wdata_rawIn_normDist_T_130=wdata_rawIn_fractIn_1[6] ? 5'h10:_wdata_rawIn_normDist_T_129; 
  assign _wdata_rawIn_normDist_T_131=wdata_rawIn_fractIn_1[7] ? 5'hf:_wdata_rawIn_normDist_T_130; 
  assign _wdata_rawIn_normDist_T_132=wdata_rawIn_fractIn_1[8] ? 5'he:_wdata_rawIn_normDist_T_131; 
  assign _wdata_rawIn_normDist_T_133=wdata_rawIn_fractIn_1[9] ? 5'hd:_wdata_rawIn_normDist_T_132; 
  assign _wdata_rawIn_normDist_T_134=wdata_rawIn_fractIn_1[10] ? 5'hc:_wdata_rawIn_normDist_T_133; 
  assign _wdata_rawIn_normDist_T_135=wdata_rawIn_fractIn_1[11] ? 5'hb:_wdata_rawIn_normDist_T_134; 
  assign _wdata_rawIn_normDist_T_136=wdata_rawIn_fractIn_1[12] ? 5'ha:_wdata_rawIn_normDist_T_135; 
  assign _wdata_rawIn_normDist_T_137=wdata_rawIn_fractIn_1[13] ? 5'h9:_wdata_rawIn_normDist_T_136; 
  assign _wdata_rawIn_normDist_T_138=wdata_rawIn_fractIn_1[14] ? 5'h8:_wdata_rawIn_normDist_T_137; 
  assign _wdata_rawIn_normDist_T_139=wdata_rawIn_fractIn_1[15] ? 5'h7:_wdata_rawIn_normDist_T_138; 
  assign _wdata_rawIn_normDist_T_140=wdata_rawIn_fractIn_1[16] ? 5'h6:_wdata_rawIn_normDist_T_139; 
  assign _wdata_rawIn_normDist_T_141=wdata_rawIn_fractIn_1[17] ? 5'h5:_wdata_rawIn_normDist_T_140; 
  assign _wdata_rawIn_normDist_T_142=wdata_rawIn_fractIn_1[18] ? 5'h4:_wdata_rawIn_normDist_T_141; 
  assign _wdata_rawIn_normDist_T_143=wdata_rawIn_fractIn_1[19] ? 5'h3:_wdata_rawIn_normDist_T_142; 
  assign _wdata_rawIn_normDist_T_144=wdata_rawIn_fractIn_1[20] ? 5'h2:_wdata_rawIn_normDist_T_143; 
  assign _wdata_rawIn_normDist_T_145=wdata_rawIn_fractIn_1[21] ? 5'h1:_wdata_rawIn_normDist_T_144; 
  assign wdata_rawIn_normDist_1=wdata_rawIn_fractIn_1[22] ? 5'h0:_wdata_rawIn_normDist_T_145; 
  assign _GEN_173={31'b0,wdata_rawIn_fractIn_1}; 
  assign _wdata_rawIn_subnormFract_T_2=_GEN_173<<wdata_rawIn_normDist_1; 
  assign wdata_rawIn_subnormFract_1={_wdata_rawIn_subnormFract_T_2[21:0],1'h0}; 
  assign _GEN_174={4'b0,wdata_rawIn_normDist_1}; 
  assign _wdata_rawIn_adjustedExp_T_5=_GEN_174^9'h1ff; 
  assign _wdata_rawIn_adjustedExp_T_6=wdata_rawIn_isZeroExpIn_1 ? _wdata_rawIn_adjustedExp_T_5:{1'b0,wdata_rawIn_expIn_1}; 
  assign _wdata_rawIn_adjustedExp_T_7=wdata_rawIn_isZeroExpIn_1 ? 2'h2:2'h1; 
  assign _GEN_175={6'b0,_wdata_rawIn_adjustedExp_T_7}; 
  assign _wdata_rawIn_adjustedExp_T_8=8'h80|_GEN_175; 
  assign _GEN_176={1'b0,_wdata_rawIn_adjustedExp_T_8}; 
  assign wdata_rawIn_adjustedExp_1=_wdata_rawIn_adjustedExp_T_6+_GEN_176; 
  assign wdata_rawIn_isZero_1=wdata_rawIn_isZeroExpIn_1&wdata_rawIn_isZeroFractIn_1; 
  assign wdata_rawIn_isSpecial_1=wdata_rawIn_adjustedExp_1[8:7]==2'h3; 
  assign wdata_rawIn_1_isNaN=wdata_rawIn_isSpecial_1&~wdata_rawIn_isZeroFractIn_1; 
  assign wdata_rawIn_1_sExp={1'b0,$signed(wdata_rawIn_adjustedExp_1)}; 
  assign wdata_rawIn_out_sig_hi_lo_1=~wdata_rawIn_isZero_1; 
  assign wdata_rawIn_out_sig_lo_1=wdata_rawIn_isZeroExpIn_1 ? wdata_rawIn_subnormFract_1:wdata_rawIn_fractIn_1; 
  assign wdata_rawIn_1_sig={1'h0,wdata_rawIn_out_sig_hi_lo_1,wdata_rawIn_out_sig_lo_1}; 
  assign _wdata_T_8=wdata_rawIn_isZero_1 ? 3'h0:wdata_rawIn_1_sExp[8:6]; 
  assign _GEN_177={2'b0,wdata_rawIn_1_isNaN}; 
  assign wdata_hi_lo_1=_wdata_T_8|_GEN_177; 
  assign wdata_lo_hi_1=wdata_rawIn_1_sExp[5:0]; 
  assign wdata_lo_lo_1=wdata_rawIn_1_sig[22:0]; 
  assign _wdata_T_10={wdata_rawIn_sign_1,wdata_hi_lo_1,wdata_lo_hi_1,wdata_lo_lo_1}; 
  assign wdata_swizzledNaN_hi_hi_hi=_wdata_T_6[64:61]; 
  assign wdata_swizzledNaN_hi_hi_lo=&_wdata_T_6[51:32]; 
  assign wdata_swizzledNaN_hi_lo_hi=_wdata_T_6[59:53]; 
  assign wdata_swizzledNaN_hi_lo_lo=_wdata_T_10[31]; 
  assign wdata_swizzledNaN_lo_hi_lo=_wdata_T_10[32]; 
  assign wdata_swizzledNaN_lo_lo=_wdata_T_10[30:0]; 
  assign wdata_swizzledNaN={wdata_swizzledNaN_hi_hi_hi,wdata_swizzledNaN_hi_hi_lo,wdata_swizzledNaN_hi_lo_hi,wdata_swizzledNaN_hi_lo_lo,_wdata_T_6[51:32],wdata_swizzledNaN_lo_hi_lo,wdata_swizzledNaN_lo_lo}; 
  assign _wdata_T_12=&_wdata_T_6[63:61]; 
  assign wdata=_wdata_T_12 ? wdata_swizzledNaN:_wdata_T_6; 
  assign _curOK_T_1=&wdata[63:61]; 
  assign _curOK_T_5=&wdata[51:32]; 
  assign _curOK_T_6=wdata[60]==_curOK_T_5; 
  assign curOK=~_curOK_T_1|_curOK_T_6; 
  assign _T_2=curOK|reset; 
  assign _GEN_178={1'b0,load_wb_tag}; 
  assign _T_5=_GEN_178+6'h20; 
  assign _T_11=~fp_decoder_io_sigs_swap12&~fp_decoder_io_sigs_swap23; 
  assign _ex_rm_T_1=ex_reg_inst[14:12]==3'h7; 
  assign _sfma_io_in_valid_T=ex_reg_valid&ex_reg_ctrl_fma; 
  assign _sfma_io_in_valid_T_1=ex_reg_ctrl_typeTagOut==2'h0; 
  assign sfma_io_in_bits_req_in1_unswizzled_hi_hi=regfile_ex_rs_0_data[31]; 
  assign sfma_io_in_bits_req_in1_unswizzled_hi_lo=regfile_ex_rs_0_data[52]; 
  assign sfma_io_in_bits_req_in1_unswizzled_lo=regfile_ex_rs_0_data[30:0]; 
  assign sfma_io_in_bits_req_in1_floats_0={sfma_io_in_bits_req_in1_unswizzled_hi_hi,sfma_io_in_bits_req_in1_unswizzled_hi_lo,sfma_io_in_bits_req_in1_unswizzled_lo}; 
  assign sfma_io_in_bits_req_in1_isbox=&regfile_ex_rs_0_data[64:60]; 
  assign _sfma_io_in_bits_req_in1_T=sfma_io_in_bits_req_in1_isbox ? 33'h0:33'he0400000; 
  assign _sfma_io_in_bits_req_in1_T_1=sfma_io_in_bits_req_in1_floats_0|_sfma_io_in_bits_req_in1_T; 
  assign sfma_io_in_bits_req_in2_unswizzled_hi_hi=regfile_ex_rs_1_data[31]; 
  assign sfma_io_in_bits_req_in2_unswizzled_hi_lo=regfile_ex_rs_1_data[52]; 
  assign sfma_io_in_bits_req_in2_unswizzled_lo=regfile_ex_rs_1_data[30:0]; 
  assign sfma_io_in_bits_req_in2_floats_0={sfma_io_in_bits_req_in2_unswizzled_hi_hi,sfma_io_in_bits_req_in2_unswizzled_hi_lo,sfma_io_in_bits_req_in2_unswizzled_lo}; 
  assign sfma_io_in_bits_req_in2_isbox=&regfile_ex_rs_1_data[64:60]; 
  assign _sfma_io_in_bits_req_in2_T=sfma_io_in_bits_req_in2_isbox ? 33'h0:33'he0400000; 
  assign _sfma_io_in_bits_req_in2_T_1=sfma_io_in_bits_req_in2_floats_0|_sfma_io_in_bits_req_in2_T; 
  assign sfma_io_in_bits_req_in3_unswizzled_hi_hi=regfile_ex_rs_2_data[31]; 
  assign sfma_io_in_bits_req_in3_unswizzled_hi_lo=regfile_ex_rs_2_data[52]; 
  assign sfma_io_in_bits_req_in3_unswizzled_lo=regfile_ex_rs_2_data[30:0]; 
  assign sfma_io_in_bits_req_in3_floats_0={sfma_io_in_bits_req_in3_unswizzled_hi_hi,sfma_io_in_bits_req_in3_unswizzled_hi_lo,sfma_io_in_bits_req_in3_unswizzled_lo}; 
  assign sfma_io_in_bits_req_in3_isbox=&regfile_ex_rs_2_data[64:60]; 
  assign _sfma_io_in_bits_req_in3_T=sfma_io_in_bits_req_in3_isbox ? 33'h0:33'he0400000; 
  assign _sfma_io_in_bits_req_in3_T_1=sfma_io_in_bits_req_in3_floats_0|_sfma_io_in_bits_req_in3_T; 
  assign _sfma_io_in_bits_req_fmaCmd_T_3=~ex_reg_ctrl_ren3&ex_reg_inst[27]; 
  assign _GEN_179={1'b0,_sfma_io_in_bits_req_fmaCmd_T_3}; 
  assign _fpiu_io_in_valid_T=ex_reg_ctrl_toint|ex_reg_ctrl_div; 
  assign _fpiu_io_in_valid_T_1=_fpiu_io_in_valid_T|ex_reg_ctrl_sqrt; 
  assign _fpiu_io_in_valid_T_2=ex_reg_ctrl_fastpipe&ex_reg_ctrl_wflags; 
  assign _fpiu_io_in_valid_T_3=_fpiu_io_in_valid_T_1|_fpiu_io_in_valid_T_2; 
  assign fpiu_io_in_bits_req_in1_hi_hi=sfma_io_in_bits_req_in1_floats_0[32]; 
  assign fpiu_io_in_bits_req_in1_fractIn=sfma_io_in_bits_req_in1_floats_0[22:0]; 
  assign fpiu_io_in_bits_req_in1_expIn=sfma_io_in_bits_req_in1_floats_0[31:23]; 
  assign _fpiu_io_in_bits_req_in1_fractOut_T={fpiu_io_in_bits_req_in1_fractIn,53'h0}; 
  assign fpiu_io_in_bits_req_in1_lo=_fpiu_io_in_bits_req_in1_fractOut_T[75:24]; 
  assign fpiu_io_in_bits_req_in1_expOut_hi=fpiu_io_in_bits_req_in1_expIn[8:6]; 
  assign _GEN_180={3'b0,fpiu_io_in_bits_req_in1_expIn}; 
  assign _fpiu_io_in_bits_req_in1_expOut_commonCase_T_1=_GEN_180+12'h800; 
  assign fpiu_io_in_bits_req_in1_expOut_commonCase=_fpiu_io_in_bits_req_in1_expOut_commonCase_T_1-12'h100; 
  assign _fpiu_io_in_bits_req_in1_expOut_T=fpiu_io_in_bits_req_in1_expOut_hi==3'h0; 
  assign _fpiu_io_in_bits_req_in1_expOut_T_1=fpiu_io_in_bits_req_in1_expOut_hi>=3'h6; 
  assign _fpiu_io_in_bits_req_in1_expOut_T_2=_fpiu_io_in_bits_req_in1_expOut_T|_fpiu_io_in_bits_req_in1_expOut_T_1; 
  assign fpiu_io_in_bits_req_in1_expOut_lo=fpiu_io_in_bits_req_in1_expOut_commonCase[8:0]; 
  assign _fpiu_io_in_bits_req_in1_expOut_T_3={fpiu_io_in_bits_req_in1_expOut_hi,fpiu_io_in_bits_req_in1_expOut_lo}; 
  assign fpiu_io_in_bits_req_in1_hi_lo=_fpiu_io_in_bits_req_in1_expOut_T_2 ? _fpiu_io_in_bits_req_in1_expOut_T_3:fpiu_io_in_bits_req_in1_expOut_commonCase; 
  assign fpiu_io_in_bits_req_in1_floats_0={fpiu_io_in_bits_req_in1_hi_hi,fpiu_io_in_bits_req_in1_hi_lo,fpiu_io_in_bits_req_in1_lo}; 
  assign fpiu_io_in_bits_req_in1_truncIdx=ex_reg_ctrl_typeTagIn[0]; 
  assign _fpiu_io_in_bits_req_in1_T_1=fpiu_io_in_bits_req_in1_truncIdx|sfma_io_in_bits_req_in1_isbox; 
  assign _fpiu_io_in_bits_req_in1_T_3=fpiu_io_in_bits_req_in1_truncIdx ? regfile_ex_rs_0_data:fpiu_io_in_bits_req_in1_floats_0; 
  assign fpiu_io_in_bits_req_in2_hi_hi=sfma_io_in_bits_req_in2_floats_0[32]; 
  assign fpiu_io_in_bits_req_in2_fractIn=sfma_io_in_bits_req_in2_floats_0[22:0]; 
  assign fpiu_io_in_bits_req_in2_expIn=sfma_io_in_bits_req_in2_floats_0[31:23]; 
  assign _fpiu_io_in_bits_req_in2_fractOut_T={fpiu_io_in_bits_req_in2_fractIn,53'h0}; 
  assign fpiu_io_in_bits_req_in2_lo=_fpiu_io_in_bits_req_in2_fractOut_T[75:24]; 
  assign fpiu_io_in_bits_req_in2_expOut_hi=fpiu_io_in_bits_req_in2_expIn[8:6]; 
  assign _GEN_181={3'b0,fpiu_io_in_bits_req_in2_expIn}; 
  assign _fpiu_io_in_bits_req_in2_expOut_commonCase_T_1=_GEN_181+12'h800; 
  assign fpiu_io_in_bits_req_in2_expOut_commonCase=_fpiu_io_in_bits_req_in2_expOut_commonCase_T_1-12'h100; 
  assign _fpiu_io_in_bits_req_in2_expOut_T=fpiu_io_in_bits_req_in2_expOut_hi==3'h0; 
  assign _fpiu_io_in_bits_req_in2_expOut_T_1=fpiu_io_in_bits_req_in2_expOut_hi>=3'h6; 
  assign _fpiu_io_in_bits_req_in2_expOut_T_2=_fpiu_io_in_bits_req_in2_expOut_T|_fpiu_io_in_bits_req_in2_expOut_T_1; 
  assign fpiu_io_in_bits_req_in2_expOut_lo=fpiu_io_in_bits_req_in2_expOut_commonCase[8:0]; 
  assign _fpiu_io_in_bits_req_in2_expOut_T_3={fpiu_io_in_bits_req_in2_expOut_hi,fpiu_io_in_bits_req_in2_expOut_lo}; 
  assign fpiu_io_in_bits_req_in2_hi_lo=_fpiu_io_in_bits_req_in2_expOut_T_2 ? _fpiu_io_in_bits_req_in2_expOut_T_3:fpiu_io_in_bits_req_in2_expOut_commonCase; 
  assign fpiu_io_in_bits_req_in2_floats_0={fpiu_io_in_bits_req_in2_hi_hi,fpiu_io_in_bits_req_in2_hi_lo,fpiu_io_in_bits_req_in2_lo}; 
  assign _fpiu_io_in_bits_req_in2_T_1=fpiu_io_in_bits_req_in1_truncIdx|sfma_io_in_bits_req_in2_isbox; 
  assign _fpiu_io_in_bits_req_in2_T_3=fpiu_io_in_bits_req_in1_truncIdx ? regfile_ex_rs_1_data:fpiu_io_in_bits_req_in2_floats_0; 
  assign _ifpu_io_in_bits_in1_T={1'b0,io_fromint_data}; 
  assign _dfma_io_in_valid_T_1=ex_reg_ctrl_typeTagOut==2'h1; 
  assign _memLatencyMask_T_2=mem_ctrl_typeTagOut==2'h0; 
  assign _memLatencyMask_T_3=mem_ctrl_fma&_memLatencyMask_T_2; 
  assign _memLatencyMask_T_4=_memLatencyMask_T_3 ? 2'h2:2'h0; 
  assign _memLatencyMask_T_5=mem_ctrl_typeTagOut==2'h1; 
  assign _memLatencyMask_T_6=mem_ctrl_fma&_memLatencyMask_T_5; 
  assign _memLatencyMask_T_7=_memLatencyMask_T_6 ? 3'h4:3'h0; 
  assign _memLatencyMask_T_8=mem_ctrl_fastpipe|mem_ctrl_fromint; 
  assign _GEN_188={1'b0,_memLatencyMask_T_8}; 
  assign _memLatencyMask_T_9=_GEN_188|_memLatencyMask_T_4; 
  assign _GEN_189={1'b0,_memLatencyMask_T_9}; 
  assign memLatencyMask=_GEN_189|_memLatencyMask_T_7; 
  assign _mem_wen_T=mem_ctrl_fma|mem_ctrl_fastpipe; 
  assign _mem_wen_T_1=_mem_wen_T|mem_ctrl_fromint; 
  assign mem_wen=mem_reg_valid&_mem_wen_T_1; 
  assign _write_port_busy_T=ex_reg_ctrl_fastpipe ? 2'h2:2'h0; 
  assign _write_port_busy_T_1=ex_reg_ctrl_fromint ? 2'h2:2'h0; 
  assign _write_port_busy_T_3=ex_reg_ctrl_fma&_sfma_io_in_valid_T_1; 
  assign _write_port_busy_T_4=_write_port_busy_T_3 ? 3'h4:3'h0; 
  assign _write_port_busy_T_6=ex_reg_ctrl_fma&_dfma_io_in_valid_T_1; 
  assign _write_port_busy_T_7=_write_port_busy_T_6 ? 4'h8:4'h0; 
  assign _write_port_busy_T_8=_write_port_busy_T|_write_port_busy_T_1; 
  assign _GEN_190={1'b0,_write_port_busy_T_8}; 
  assign _write_port_busy_T_9=_GEN_190|_write_port_busy_T_4; 
  assign _GEN_191={1'b0,_write_port_busy_T_9}; 
  assign _write_port_busy_T_10=_GEN_191|_write_port_busy_T_7; 
  assign _GEN_192={1'b0,memLatencyMask}; 
  assign _write_port_busy_T_11=_GEN_192&_write_port_busy_T_10; 
  assign _write_port_busy_T_12=|_write_port_busy_T_11; 
  assign _write_port_busy_T_13=mem_wen&_write_port_busy_T_12; 
  assign _write_port_busy_T_14=ex_reg_ctrl_fastpipe ? 3'h4:3'h0; 
  assign _write_port_busy_T_15=ex_reg_ctrl_fromint ? 3'h4:3'h0; 
  assign _write_port_busy_T_18=_write_port_busy_T_3 ? 4'h8:4'h0; 
  assign _write_port_busy_T_21=_write_port_busy_T_6 ? 5'h10:5'h0; 
  assign _write_port_busy_T_22=_write_port_busy_T_14|_write_port_busy_T_15; 
  assign _GEN_193={1'b0,_write_port_busy_T_22}; 
  assign _write_port_busy_T_23=_GEN_193|_write_port_busy_T_18; 
  assign _GEN_194={1'b0,_write_port_busy_T_23}; 
  assign _write_port_busy_T_24=_GEN_194|_write_port_busy_T_21; 
  assign _GEN_195={2'b0,wen}; 
  assign _write_port_busy_T_25=_GEN_195&_write_port_busy_T_24; 
  assign _write_port_busy_T_26=|_write_port_busy_T_25; 
  assign _write_port_busy_T_27=_write_port_busy_T_13|_write_port_busy_T_26; 
  assign _GEN_114=wen[1] ? wbInfo_1_typeTag:wbInfo_0_typeTag; 
  assign _GEN_118=wen[2] ? wbInfo_2_typeTag:wbInfo_1_typeTag; 
  assign _GEN_196={1'b0,wen[2:1]}; 
  assign _wen_T_2=_GEN_196|memLatencyMask; 
  assign _T_20=~write_port_busy&memLatencyMask[0]; 
  assign _wbInfo_0_pipeid_T_7=_memLatencyMask_T_6 ? 2'h3:2'h0; 
  assign _GEN_197={1'b0,mem_ctrl_fromint}; 
  assign _wbInfo_0_pipeid_T_9=_GEN_197|_memLatencyMask_T_4; 
  assign _wbInfo_0_pipeid_T_10=_wbInfo_0_pipeid_T_9|_wbInfo_0_pipeid_T_7; 
  assign _GEN_123=_T_20 ? mem_ctrl_typeTagOut:{1'b0,_GEN_114}; 
  assign _T_23=~write_port_busy&memLatencyMask[1]; 
  assign _GEN_127=_T_23 ? mem_ctrl_typeTagOut:{1'b0,_GEN_118}; 
  assign _T_26=~write_port_busy&memLatencyMask[2]; 
  assign _GEN_131=_T_26 ? mem_ctrl_typeTagOut:{1'b0,wbInfo_2_typeTag}; 
  assign _GEN_136=mem_wen ? _GEN_123:{1'b0,_GEN_114}; 
  assign _GEN_140=mem_wen ? _GEN_127:{1'b0,_GEN_118}; 
  assign _GEN_144=mem_wen ? _GEN_131:{1'b0,wbInfo_2_typeTag}; 
  assign divSqrt_typeTag=divSqrt_1_io_outValid_div|divSqrt_1_io_outValid_sqrt; 
  assign _T_52=divSqrt_io_outValid_div|divSqrt_io_outValid_sqrt; 
  assign _GEN_158=_T_52&~divSqrt_killed; 
  assign divSqrt_wen=divSqrt_typeTag ? ~divSqrt_killed:_GEN_158; 
  assign waddr=divSqrt_wen ? divSqrt_waddr:wbInfo_0_rd; 
  assign wtypeTag=divSqrt_wen ? divSqrt_typeTag:wbInfo_0_typeTag; 
  assign _wdata_T_13=wbInfo_0_pipeid==2'h1; 
  assign _wdata_T_14=_wdata_T_13 ? ifpu_io_out_bits_data:fpmu_io_out_bits_data; 
  assign _wdata_T_15=wbInfo_0_pipeid==2'h2; 
  assign _wdata_T_16=_wdata_T_15 ? sfma_io_out_bits_data:_wdata_T_14; 
  assign _wdata_T_17=wbInfo_0_pipeid==2'h3; 
  assign _wdata_T_18=_wdata_T_17 ? dfma_io_out_bits_data:_wdata_T_16; 
  assign _divSqrt_wdata_T_1=&divSqrt_1_io_out[63:61]; 
  assign divSqrt_wdata_maskedNaN=divSqrt_1_io_out&65'h1efefffffffffffff; 
  assign _divSqrt_wdata_T_2=_divSqrt_wdata_T_1 ? divSqrt_wdata_maskedNaN:divSqrt_1_io_out; 
  assign _GEN_159=divSqrt_io_out; 
  assign divSqrt_wdata=divSqrt_typeTag ? _divSqrt_wdata_T_2:{32'b0,_GEN_159}; 
  assign _wdata_T_19=divSqrt_wen ? divSqrt_wdata:_wdata_T_18; 
  assign wdata_opts_bigger_swizzledNaN_hi_hi_lo=&20'hfffff; 
  assign wdata_opts_bigger_swizzledNaN_hi_lo_lo=_wdata_T_19[31]; 
  assign wdata_opts_bigger_swizzledNaN_lo_hi_lo=_wdata_T_19[32]; 
  assign wdata_opts_bigger_swizzledNaN_lo_lo=_wdata_T_19[30:0]; 
  assign wdata_opts_bigger_swizzledNaN={4'hf,wdata_opts_bigger_swizzledNaN_hi_hi_lo,7'h7f,wdata_opts_bigger_swizzledNaN_hi_lo_lo,20'hfffff,wdata_opts_bigger_swizzledNaN_lo_hi_lo,wdata_opts_bigger_swizzledNaN_lo_lo}; 
  assign _wdata_opts_bigger_T=&3'h7; 
  assign wdata_opts_bigger=_wdata_opts_bigger_T ? wdata_opts_bigger_swizzledNaN:65'h1ffffffffffffffff; 
  assign wdata_1=wtypeTag ? _wdata_T_19:wdata_opts_bigger; 
  assign _wexc_T_1=_wdata_T_13 ? ifpu_io_out_bits_exc:fpmu_io_out_bits_exc; 
  assign _wexc_T_3=_wdata_T_15 ? sfma_io_out_bits_exc:_wexc_T_1; 
  assign wexc=_wdata_T_17 ? dfma_io_out_bits_exc:_wexc_T_3; 
  assign frfWriteBundle_1_wrenf=wen[0]|divSqrt_wen; 
  assign unswizzled_hi_hi_1=wdata_1[31]; 
  assign unswizzled_hi_lo_1=wdata_1[52]; 
  assign unswizzled_lo_1=wdata_1[30:0]; 
  assign unswizzled_1={unswizzled_hi_hi_1,unswizzled_hi_lo_1,unswizzled_lo_1}; 
  assign _curOK_T_8=&wdata_1[63:61]; 
  assign _curOK_T_12=&wdata_1[51:32]; 
  assign _curOK_T_13=wdata_1[60]==_curOK_T_12; 
  assign curOK_1=~_curOK_T_8|_curOK_T_13; 
  assign _T_33=curOK_1|reset; 
  assign _GEN_200={1'b0,waddr}; 
  assign _T_36=_GEN_200+6'h20; 
  assign unrecoded_rawIn_exp=wdata_1[63:52]; 
  assign unrecoded_rawIn_isZero=unrecoded_rawIn_exp[11:9]==3'h0; 
  assign unrecoded_rawIn_isSpecial=unrecoded_rawIn_exp[11:10]==2'h3; 
  assign unrecoded_rawIn__isNaN=unrecoded_rawIn_isSpecial&unrecoded_rawIn_exp[9]; 
  assign unrecoded_rawIn__isInf=unrecoded_rawIn_isSpecial&~unrecoded_rawIn_exp[9]; 
  assign unrecoded_rawIn__sign=wdata_1[64]; 
  assign unrecoded_rawIn__sExp={1'b0,$signed(unrecoded_rawIn_exp)}; 
  assign unrecoded_rawIn_out_sig_hi_lo=~unrecoded_rawIn_isZero; 
  assign unrecoded_rawIn_out_sig_lo=wdata_1[51:0]; 
  assign unrecoded_rawIn__sig={1'h0,unrecoded_rawIn_out_sig_hi_lo,unrecoded_rawIn_out_sig_lo}; 
  assign unrecoded_isSubnormal=$signed(unrecoded_rawIn__sExp)<13'sh402; 
  assign unrecoded_denormShiftDist=6'h1-unrecoded_rawIn__sExp[5:0]; 
  assign _unrecoded_denormFract_T_1=unrecoded_rawIn__sig[53:1]>>unrecoded_denormShiftDist; 
  assign unrecoded_denormFract=_unrecoded_denormFract_T_1[51:0]; 
  assign _unrecoded_expOut_T_2=unrecoded_rawIn__sExp[10:0]-11'h401; 
  assign _unrecoded_expOut_T_3=unrecoded_isSubnormal ? 11'h0:_unrecoded_expOut_T_2; 
  assign _unrecoded_expOut_T_4=unrecoded_rawIn__isNaN|unrecoded_rawIn__isInf; 
  assign _unrecoded_expOut_T_6=_unrecoded_expOut_T_4 ? 11'h7ff:11'h0; 
  assign unrecoded_hi_lo=_unrecoded_expOut_T_3|_unrecoded_expOut_T_6; 
  assign _unrecoded_fractOut_T_1=unrecoded_rawIn__isInf ? 52'h0:unrecoded_rawIn__sig[51:0]; 
  assign unrecoded_lo=unrecoded_isSubnormal ? unrecoded_denormFract:_unrecoded_fractOut_T_1; 
  assign unrecoded={unrecoded_rawIn__sign,unrecoded_hi_lo,unrecoded_lo}; 
  assign prevUnrecoded_rawIn_exp=unswizzled_1[31:23]; 
  assign prevUnrecoded_rawIn_isZero=prevUnrecoded_rawIn_exp[8:6]==3'h0; 
  assign prevUnrecoded_rawIn_isSpecial=prevUnrecoded_rawIn_exp[8:7]==2'h3; 
  assign prevUnrecoded_rawIn__isNaN=prevUnrecoded_rawIn_isSpecial&prevUnrecoded_rawIn_exp[6]; 
  assign prevUnrecoded_rawIn__isInf=prevUnrecoded_rawIn_isSpecial&~prevUnrecoded_rawIn_exp[6]; 
  assign prevUnrecoded_rawIn__sign=unswizzled_1[32]; 
  assign prevUnrecoded_rawIn__sExp={1'b0,$signed(prevUnrecoded_rawIn_exp)}; 
  assign prevUnrecoded_rawIn_out_sig_hi_lo=~prevUnrecoded_rawIn_isZero; 
  assign prevUnrecoded_rawIn_out_sig_lo=unswizzled_1[22:0]; 
  assign prevUnrecoded_rawIn__sig={1'h0,prevUnrecoded_rawIn_out_sig_hi_lo,prevUnrecoded_rawIn_out_sig_lo}; 
  assign prevUnrecoded_isSubnormal=$signed(prevUnrecoded_rawIn__sExp)<10'sh82; 
  assign prevUnrecoded_denormShiftDist=5'h1-prevUnrecoded_rawIn__sExp[4:0]; 
  assign _prevUnrecoded_denormFract_T_1=prevUnrecoded_rawIn__sig[24:1]>>prevUnrecoded_denormShiftDist; 
  assign prevUnrecoded_denormFract=_prevUnrecoded_denormFract_T_1[22:0]; 
  assign _prevUnrecoded_expOut_T_2=prevUnrecoded_rawIn__sExp[7:0]-8'h81; 
  assign _prevUnrecoded_expOut_T_3=prevUnrecoded_isSubnormal ? 8'h0:_prevUnrecoded_expOut_T_2; 
  assign _prevUnrecoded_expOut_T_4=prevUnrecoded_rawIn__isNaN|prevUnrecoded_rawIn__isInf; 
  assign _prevUnrecoded_expOut_T_6=_prevUnrecoded_expOut_T_4 ? 8'hff:8'h0; 
  assign prevUnrecoded_hi_lo=_prevUnrecoded_expOut_T_3|_prevUnrecoded_expOut_T_6; 
  assign _prevUnrecoded_fractOut_T_1=prevUnrecoded_rawIn__isInf ? 23'h0:prevUnrecoded_rawIn__sig[22:0]; 
  assign prevUnrecoded_lo=prevUnrecoded_isSubnormal ? prevUnrecoded_denormFract:_prevUnrecoded_fractOut_T_1; 
  assign prevUnrecoded={prevUnrecoded_rawIn__sign,prevUnrecoded_hi_lo,prevUnrecoded_lo}; 
  assign hi=unrecoded[63:32]; 
  assign lo=_curOK_T_8 ? prevUnrecoded:unrecoded[31:0]; 
  assign _T_40={hi,lo}; 
  assign wb_toint_valid=wb_reg_valid&wb_ctrl_toint; 
  assign _io_fcsr_flags_valid_T=wb_toint_valid|divSqrt_wen; 
  assign _io_fcsr_flags_bits_T=wb_toint_valid ? wb_toint_exc:5'h0; 
  assign _GEN_160=divSqrt_io_exceptionFlags; 
  assign divSqrt_flags=divSqrt_typeTag ? divSqrt_1_io_exceptionFlags:_GEN_160; 
  assign _io_fcsr_flags_bits_T_1=divSqrt_wen ? divSqrt_flags:5'h0; 
  assign _io_fcsr_flags_bits_T_2=_io_fcsr_flags_bits_T|_io_fcsr_flags_bits_T_1; 
  assign _io_fcsr_flags_bits_T_4=wen[0] ? wexc:5'h0; 
  assign _divSqrt_write_port_busy_T=mem_ctrl_div|mem_ctrl_sqrt; 
  assign _divSqrt_write_port_busy_T_1=|wen; 
  assign divSqrt_write_port_busy=_divSqrt_write_port_busy_T&_divSqrt_write_port_busy_T_1; 
  assign _io_fcsr_rdy_T=ex_reg_valid&ex_reg_ctrl_wflags; 
  assign _io_fcsr_rdy_T_1=mem_reg_valid&mem_ctrl_wflags; 
  assign _io_fcsr_rdy_T_2=_io_fcsr_rdy_T|_io_fcsr_rdy_T_1; 
  assign _io_fcsr_rdy_T_4=_io_fcsr_rdy_T_2|wb_toint_valid; 
  assign _io_fcsr_rdy_T_6=_io_fcsr_rdy_T_4|_divSqrt_write_port_busy_T_1; 
  assign _GEN_162=~divSqrt_1_io_inReady|~divSqrt_io_inReady; 
  assign divSqrt_inFlight=divSqrt_killed ? 1'h0:_GEN_162; 
  assign _io_fcsr_rdy_T_7=_io_fcsr_rdy_T_6|divSqrt_inFlight; 
  assign _io_nack_mem_T=write_port_busy|divSqrt_write_port_busy; 
  assign _io_sboard_set_x27_T_3=_memLatencyMask_T_6|mem_ctrl_div; 
  assign _io_sboard_clr_T_4=wen[0]&_wdata_T_17; 
  assign _io_illegal_rm_T_1=io_inst[14:12]==3'h5; 
  assign _io_illegal_rm_T_2=io_inst[14:12]==3'h6; 
  assign _io_illegal_rm_T_3=_io_illegal_rm_T_1|_io_illegal_rm_T_2; 
  assign _io_illegal_rm_T_5=io_inst[14:12]==3'h7; 
  assign _io_illegal_rm_T_6=io_fcsr_rm>=3'h5; 
  assign _io_illegal_rm_T_7=_io_illegal_rm_T_5&_io_illegal_rm_T_6; 
  assign _divSqrt_inValid_T_1=mem_reg_valid&_divSqrt_write_port_busy_T; 
  assign divSqrt_inValid=_divSqrt_inValid_T_1&~divSqrt_inFlight; 
  assign _divSqrt_killed_T=divSqrt_inValid&killm; 
  assign divSqrt_io_a_hi_hi=fpiu_io_out_bits_in_in1[64]; 
  assign divSqrt_io_a_fractIn=fpiu_io_out_bits_in_in1[51:0]; 
  assign divSqrt_io_a_expIn=fpiu_io_out_bits_in_in1[63:52]; 
  assign _divSqrt_io_a_fractOut_T={divSqrt_io_a_fractIn,24'h0}; 
  assign divSqrt_io_a_lo=_divSqrt_io_a_fractOut_T[75:53]; 
  assign divSqrt_io_a_expOut_hi=divSqrt_io_a_expIn[11:9]; 
  assign _divSqrt_io_a_expOut_commonCase_T_1=divSqrt_io_a_expIn+12'h100; 
  assign divSqrt_io_a_expOut_commonCase=_divSqrt_io_a_expOut_commonCase_T_1-12'h800; 
  assign _divSqrt_io_a_expOut_T=divSqrt_io_a_expOut_hi==3'h0; 
  assign _divSqrt_io_a_expOut_T_1=divSqrt_io_a_expOut_hi>=3'h6; 
  assign _divSqrt_io_a_expOut_T_2=_divSqrt_io_a_expOut_T|_divSqrt_io_a_expOut_T_1; 
  assign divSqrt_io_a_expOut_lo=divSqrt_io_a_expOut_commonCase[5:0]; 
  assign _divSqrt_io_a_expOut_T_3={divSqrt_io_a_expOut_hi,divSqrt_io_a_expOut_lo}; 
  assign divSqrt_io_a_hi_lo=_divSqrt_io_a_expOut_T_2 ? _divSqrt_io_a_expOut_T_3:divSqrt_io_a_expOut_commonCase[8:0]; 
  assign divSqrt_io_a_hi={divSqrt_io_a_hi_hi,divSqrt_io_a_hi_lo}; 
  assign divSqrt_io_b_hi_hi=fpiu_io_out_bits_in_in2[64]; 
  assign divSqrt_io_b_fractIn=fpiu_io_out_bits_in_in2[51:0]; 
  assign divSqrt_io_b_expIn=fpiu_io_out_bits_in_in2[63:52]; 
  assign _divSqrt_io_b_fractOut_T={divSqrt_io_b_fractIn,24'h0}; 
  assign divSqrt_io_b_lo=_divSqrt_io_b_fractOut_T[75:53]; 
  assign divSqrt_io_b_expOut_hi=divSqrt_io_b_expIn[11:9]; 
  assign _divSqrt_io_b_expOut_commonCase_T_1=divSqrt_io_b_expIn+12'h100; 
  assign divSqrt_io_b_expOut_commonCase=_divSqrt_io_b_expOut_commonCase_T_1-12'h800; 
  assign _divSqrt_io_b_expOut_T=divSqrt_io_b_expOut_hi==3'h0; 
  assign _divSqrt_io_b_expOut_T_1=divSqrt_io_b_expOut_hi>=3'h6; 
  assign _divSqrt_io_b_expOut_T_2=_divSqrt_io_b_expOut_T|_divSqrt_io_b_expOut_T_1; 
  assign divSqrt_io_b_expOut_lo=divSqrt_io_b_expOut_commonCase[5:0]; 
  assign _divSqrt_io_b_expOut_T_3={divSqrt_io_b_expOut_hi,divSqrt_io_b_expOut_lo}; 
  assign divSqrt_io_b_hi_lo=_divSqrt_io_b_expOut_T_2 ? _divSqrt_io_b_expOut_T_3:divSqrt_io_b_expOut_commonCase[8:0]; 
  assign divSqrt_io_b_hi={divSqrt_io_b_hi_hi,divSqrt_io_b_hi_lo}; 
  assign io_fcsr_flags_valid=_io_fcsr_flags_valid_T|wen[0]; 
  assign io_fcsr_flags_bits=_io_fcsr_flags_bits_T_2|_io_fcsr_flags_bits_T_4; 
  assign io_store_data=fpiu_io_out_bits_store; 
  assign io_toint_data=fpiu_io_out_bits_toint; 
  assign io_fcsr_rdy=~_io_fcsr_rdy_T_7; 
  assign io_nack_mem=_io_nack_mem_T|divSqrt_inFlight; 
  assign io_illegal_rm=_io_illegal_rm_T_3|_io_illegal_rm_T_7; 
  assign io_dec_wen=fp_decoder_io_sigs_wen; 
  assign io_dec_ren1=fp_decoder_io_sigs_ren1; 
  assign io_dec_ren2=fp_decoder_io_sigs_ren2; 
  assign io_dec_ren3=fp_decoder_io_sigs_ren3; 
  assign io_sboard_set=wb_reg_valid&io_sboard_set_REG; 
  assign io_sboard_clr=divSqrt_wen|_io_sboard_clr_T_4; 
  assign io_sboard_clra=divSqrt_wen ? divSqrt_waddr:wbInfo_0_rd; 
  assign fp_decoder_io_inst=io_inst; 
  assign sfma_clock=clock; 
  assign sfma_reset=reset; 
  assign sfma_io_in_valid=_sfma_io_in_valid_T&_sfma_io_in_valid_T_1; 
  assign sfma_io_in_bits_ren3=ex_reg_ctrl_ren3; 
  assign sfma_io_in_bits_swap23=ex_reg_ctrl_swap23; 
  assign sfma_io_in_bits_rm=_ex_rm_T_1 ? io_fcsr_rm:ex_reg_inst[14:12]; 
  assign sfma_io_in_bits_fmaCmd=ex_reg_inst[3:2]|_GEN_179; 
  assign sfma_io_in_bits_in1={32'b0,_sfma_io_in_bits_req_in1_T_1}; 
  assign sfma_io_in_bits_in2={32'b0,_sfma_io_in_bits_req_in2_T_1}; 
  assign sfma_io_in_bits_in3={32'b0,_sfma_io_in_bits_req_in3_T_1}; 
  assign fpiu_clock=clock; 
  assign fpiu_io_in_valid=ex_reg_valid&_fpiu_io_in_valid_T_3; 
  assign fpiu_io_in_bits_ren2=ex_reg_ctrl_ren2; 
  assign fpiu_io_in_bits_typeTagIn=ex_reg_ctrl_typeTagIn; 
  assign fpiu_io_in_bits_typeTagOut=ex_reg_ctrl_typeTagOut; 
  assign fpiu_io_in_bits_wflags=ex_reg_ctrl_wflags; 
  assign fpiu_io_in_bits_rm=_ex_rm_T_1 ? io_fcsr_rm:ex_reg_inst[14:12]; 
  assign fpiu_io_in_bits_typ=ex_reg_inst[21:20]; 
  assign fpiu_io_in_bits_fmt=ex_reg_inst[26:25]; 
  assign fpiu_io_in_bits_in1=_fpiu_io_in_bits_req_in1_T_1 ? _fpiu_io_in_bits_req_in1_T_3:65'he008000000000000; 
  assign fpiu_io_in_bits_in2=_fpiu_io_in_bits_req_in2_T_1 ? _fpiu_io_in_bits_req_in2_T_3:65'he008000000000000; 
  assign ifpu_clock=clock; 
  assign ifpu_reset=reset; 
  assign ifpu_io_in_valid=ex_reg_valid&ex_reg_ctrl_fromint; 
  assign ifpu_io_in_bits_typeTagIn=fpiu_io_in_bits_typeTagIn; 
  assign ifpu_io_in_bits_wflags=fpiu_io_in_bits_wflags; 
  assign ifpu_io_in_bits_rm=fpiu_io_in_bits_rm; 
  assign ifpu_io_in_bits_typ=fpiu_io_in_bits_typ; 
  assign ifpu_io_in_bits_in1=_ifpu_io_in_bits_in1_T[63:0]; 
  assign fpmu_clock=clock; 
  assign fpmu_reset=reset; 
  assign fpmu_io_in_valid=ex_reg_valid&ex_reg_ctrl_fastpipe; 
  assign fpmu_io_in_bits_ren2=fpiu_io_in_bits_ren2; 
  assign fpmu_io_in_bits_typeTagOut=fpiu_io_in_bits_typeTagOut; 
  assign fpmu_io_in_bits_wflags=fpiu_io_in_bits_wflags; 
  assign fpmu_io_in_bits_rm=fpiu_io_in_bits_rm; 
  assign fpmu_io_in_bits_in1=fpiu_io_in_bits_in1; 
  assign fpmu_io_in_bits_in2=fpiu_io_in_bits_in2; 
  assign fpmu_io_lt=fpiu_io_out_bits_lt; 
  assign dfma_clock=clock; 
  assign dfma_reset=reset; 
  assign dfma_io_in_valid=_sfma_io_in_valid_T&_dfma_io_in_valid_T_1; 
  assign dfma_io_in_bits_ren3=ex_reg_ctrl_ren3; 
  assign dfma_io_in_bits_swap23=ex_reg_ctrl_swap23; 
  assign dfma_io_in_bits_rm=_ex_rm_T_1 ? io_fcsr_rm:ex_reg_inst[14:12]; 
  assign dfma_io_in_bits_fmaCmd=ex_reg_inst[3:2]|_GEN_179; 
  assign dfma_io_in_bits_in1=regfile_ex_rs_0_data; 
  assign dfma_io_in_bits_in2=regfile_ex_rs_1_data; 
  assign dfma_io_in_bits_in3=regfile_ex_rs_2_data; 
  assign divSqrt_clock=clock; 
  assign divSqrt_reset=divSqrt_killed; 
  assign divSqrt_io_inValid=divSqrt_inValid&_memLatencyMask_T_2; 
  assign divSqrt_io_sqrtOp=mem_ctrl_sqrt; 
  assign divSqrt_io_a={divSqrt_io_a_hi,divSqrt_io_a_lo}; 
  assign divSqrt_io_b={divSqrt_io_b_hi,divSqrt_io_b_lo}; 
  assign divSqrt_io_roundingMode=fpiu_io_out_bits_in_rm; 
  assign divSqrt_1_clock=clock; 
  assign divSqrt_1_reset=divSqrt_killed; 
  assign divSqrt_1_io_inValid=divSqrt_inValid&_memLatencyMask_T_5; 
  assign divSqrt_1_io_sqrtOp=mem_ctrl_sqrt; 
  assign divSqrt_1_io_a=fpiu_io_out_bits_in_in1; 
  assign divSqrt_1_io_b=fpiu_io_out_bits_in_in2; 
  assign divSqrt_1_io_roundingMode=fpiu_io_out_bits_in_rm; 
  assign FPU_cov_read_addr=FPU_state; 
  assign FPU_cov_read_data=FPU_cov[FPU_cov_read_addr]; 
  assign FPU_cov_write_data=1'h1; 
  assign FPU_cov_write_addr=FPU_state; 
  assign FPU_cov_write_mask=1'h1; 
  assign FPU_cov_write_en=1'h1; 
  assign wbInfo_0_typeTag_shl={wbInfo_0_typeTag,16'h0}; 
  assign wbInfo_0_typeTag_pad={3'h0,wbInfo_0_typeTag_shl}; 
  assign wb_reg_valid_shl={wb_reg_valid,2'h0}; 
  assign wb_reg_valid_pad={17'h0,wb_reg_valid_shl}; 
  assign mem_ctrl_sqrt_shl={mem_ctrl_sqrt,7'h0}; 
  assign mem_ctrl_sqrt_pad={12'h0,mem_ctrl_sqrt_shl}; 
  assign divSqrt_killed_shl={divSqrt_killed,19'h0}; 
  assign divSqrt_killed_pad=divSqrt_killed_shl; 
  assign ex_reg_ctrl_typeTagIn_shl={ex_reg_ctrl_typeTagIn,7'h0}; 
  assign ex_reg_ctrl_typeTagIn_pad={11'h0,ex_reg_ctrl_typeTagIn_shl}; 
  assign ex_reg_ctrl_fromint_shl={ex_reg_ctrl_fromint,2'h0}; 
  assign ex_reg_ctrl_fromint_pad={17'h0,ex_reg_ctrl_fromint_shl}; 
  assign mem_ctrl_typeTagOut_shl={mem_ctrl_typeTagOut,7'h0}; 
  assign mem_ctrl_typeTagOut_pad={11'h0,mem_ctrl_typeTagOut_shl}; 
  assign wen_shl={wen,5'h0}; 
  assign wen_pad={12'h0,wen_shl}; 
  assign wb_ctrl_toint_shl={wb_ctrl_toint,11'h0}; 
  assign wb_ctrl_toint_pad={8'h0,wb_ctrl_toint_shl}; 
  assign ex_reg_ctrl_fastpipe_shl={ex_reg_ctrl_fastpipe,18'h0}; 
  assign ex_reg_ctrl_fastpipe_pad={1'h0,ex_reg_ctrl_fastpipe_shl}; 
  assign write_port_busy_shl={write_port_busy,14'h0}; 
  assign write_port_busy_pad={5'h0,write_port_busy_shl}; 
  assign mem_ctrl_fastpipe_shl={mem_ctrl_fastpipe,5'h0}; 
  assign mem_ctrl_fastpipe_pad={14'h0,mem_ctrl_fastpipe_shl}; 
  assign ex_reg_ctrl_typeTagOut_shl={ex_reg_ctrl_typeTagOut,13'h0}; 
  assign ex_reg_ctrl_typeTagOut_pad={5'h0,ex_reg_ctrl_typeTagOut_shl}; 
  assign mem_reg_valid_shl={mem_reg_valid,17'h0}; 
  assign mem_reg_valid_pad={2'h0,mem_reg_valid_shl}; 
  assign mem_ctrl_div_shl={mem_ctrl_div,13'h0}; 
  assign mem_ctrl_div_pad={6'h0,mem_ctrl_div_shl}; 
  assign wbInfo_0_pipeid_shl={wbInfo_0_pipeid,10'h0}; 
  assign wbInfo_0_pipeid_pad={8'h0,wbInfo_0_pipeid_shl}; 
  assign mem_ctrl_toint_shl={mem_ctrl_toint,1'h0}; 
  assign mem_ctrl_toint_pad={18'h0,mem_ctrl_toint_shl}; 
  assign ex_reg_ctrl_fma_shl={ex_reg_ctrl_fma,4'h0}; 
  assign ex_reg_ctrl_fma_pad={15'h0,ex_reg_ctrl_fma_shl}; 
  assign ex_reg_valid_shl={ex_reg_valid,3'h0}; 
  assign ex_reg_valid_pad={16'h0,ex_reg_valid_shl}; 
  assign mem_ctrl_fromint_shl={mem_ctrl_fromint,10'h0}; 
  assign mem_ctrl_fromint_pad={9'h0,mem_ctrl_fromint_shl}; 
  assign mem_ctrl_fma_shl={mem_ctrl_fma,2'h0}; 
  assign mem_ctrl_fma_pad={17'h0,mem_ctrl_fma_shl}; 
  assign FPU_xor7=wbInfo_0_typeTag_pad^wb_reg_valid_pad; 
  assign FPU_xor18=divSqrt_killed_pad^ex_reg_ctrl_typeTagIn_pad; 
  assign FPU_xor8=mem_ctrl_sqrt_pad^FPU_xor18; 
  assign FPU_xor3=FPU_xor7^FPU_xor8; 
  assign FPU_xor9=ex_reg_ctrl_fromint_pad^mem_ctrl_typeTagOut_pad; 
  assign FPU_xor22=wb_ctrl_toint_pad^ex_reg_ctrl_fastpipe_pad; 
  assign FPU_xor10=wen_pad^FPU_xor22; 
  assign FPU_xor4=FPU_xor9^FPU_xor10; 
  assign FPU_xor1=FPU_xor3^FPU_xor4; 
  assign FPU_xor11=write_port_busy_pad^mem_ctrl_fastpipe_pad; 
  assign FPU_xor26=mem_reg_valid_pad^mem_ctrl_div_pad; 
  assign FPU_xor12=ex_reg_ctrl_typeTagOut_pad^FPU_xor26; 
  assign FPU_xor5=FPU_xor11^FPU_xor12; 
  assign FPU_xor28=mem_ctrl_toint_pad^ex_reg_ctrl_fma_pad; 
  assign FPU_xor13=wbInfo_0_pipeid_pad^FPU_xor28; 
  assign FPU_xor30=mem_ctrl_fromint_pad^mem_ctrl_fma_pad; 
  assign FPU_xor14=ex_reg_valid_pad^FPU_xor30; 
  assign FPU_xor6=FPU_xor13^FPU_xor14; 
  assign FPU_xor2=FPU_xor5^FPU_xor6; 
  assign FPU_xor0=FPU_xor1^FPU_xor2; 
  assign fpiu_sum=FPU_covSum+fpiu_io_covSum; 
  assign fp_decoder_sum=fpiu_sum+fp_decoder_io_covSum; 
  assign ifpu_sum=fp_decoder_sum+ifpu_io_covSum; 
  assign sfma_sum=ifpu_sum+sfma_io_covSum; 
  assign fpmu_sum=sfma_sum+fpmu_io_covSum; 
  assign divSqrt_1_sum=fpmu_sum+divSqrt_1_io_covSum; 
  assign dfma_sum=divSqrt_1_sum+dfma_io_covSum; 
  assign divSqrt_sum=dfma_sum+divSqrt_io_covSum; 
  assign io_covSum=divSqrt_sum; 
  assign stopEn0=load_wb&~_T_2; 
  assign stopEn1=frfWriteBundle_1_wrenf&~_T_33; 
  assign fpiu_metaAssert_wire=fpiu_metaAssert; 
  assign divSqrt_metaAssert_wire=divSqrt_metaAssert; 
  assign fp_decoder_metaAssert_wire=fp_decoder_metaAssert; 
  assign dfma_metaAssert_wire=dfma_metaAssert; 
  assign ifpu_metaAssert_wire=ifpu_metaAssert; 
  assign divSqrt_1_metaAssert_wire=divSqrt_1_metaAssert; 
  assign sfma_metaAssert_wire=sfma_metaAssert; 
  assign fpmu_metaAssert_wire=fpmu_metaAssert; 
  assign FPU_or3=stopEn0|stopEn1; 
  assign FPU_or10=divSqrt_metaAssert_wire|divSqrt_1_metaAssert_wire; 
  assign FPU_or4=fp_decoder_metaAssert_wire|FPU_or10; 
  assign FPU_or1=FPU_or3|FPU_or4; 
  assign FPU_or5=fpiu_metaAssert_wire|dfma_metaAssert_wire; 
  assign FPU_or14=ifpu_metaAssert_wire|sfma_metaAssert_wire; 
  assign FPU_or6=fpmu_metaAssert_wire|FPU_or14; 
  assign FPU_or2=FPU_or5|FPU_or6; 
  assign FPU_or0=FPU_or1|FPU_or2; 
  assign metaAssert=FPU_metaAssert; 
  assign fpiu_metaReset=metaReset|fpiu_halt; 
  assign ifpu_metaReset=metaReset|ifpu_halt; 
  assign sfma_metaReset=metaReset|sfma_halt; 
  assign fpmu_metaReset=metaReset|fpmu_halt; 
  assign divSqrt_1_metaReset=metaReset|divSqrt_1_halt; 
  assign dfma_metaReset=metaReset|dfma_halt; 
  assign divSqrt_metaReset=metaReset|divSqrt_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (regfile_MPORT_en&regfile_MPORT_mask)
            begin 
              regfile [regfile_MPORT_addr]<=regfile_MPORT_data;
            end 
         if (regfile_MPORT_1_en&regfile_MPORT_1_mask)
            begin 
              regfile [regfile_MPORT_1_addr]<=regfile_MPORT_1_data;
            end 
         if (metaReset)
            begin 
              ex_reg_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 ex_reg_valid <=1'h0;
               end 
             else 
               begin 
                 ex_reg_valid <=io_valid;
               end 
         if (metaReset)
            begin 
              ex_reg_inst <=32'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_inst <=io_inst;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_ren2 <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_ren2 <=fp_decoder_io_sigs_ren2;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_ren3 <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_ren3 <=fp_decoder_io_sigs_ren3;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_swap23 <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_swap23 <=fp_decoder_io_sigs_swap23;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_typeTagIn <=2'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_typeTagIn <=fp_decoder_io_sigs_typeTagIn;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_typeTagOut <=2'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_typeTagOut <=fp_decoder_io_sigs_typeTagOut;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_fromint <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_fromint <=fp_decoder_io_sigs_fromint;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_toint <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_toint <=fp_decoder_io_sigs_toint;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_fastpipe <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_fastpipe <=fp_decoder_io_sigs_fastpipe;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_fma <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_fma <=fp_decoder_io_sigs_fma;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_div <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_div <=fp_decoder_io_sigs_div;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_sqrt <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_sqrt <=fp_decoder_io_sigs_sqrt;
               end 
         if (metaReset)
            begin 
              ex_reg_ctrl_wflags <=1'h0;
            end 
          else 
            if (io_valid)
               begin 
                 ex_reg_ctrl_wflags <=fp_decoder_io_sigs_wflags;
               end 
         if (metaReset)
            begin 
              ex_ra_0 <=5'h0;
            end 
          else 
            if (io_valid)
               begin 
                 if (fp_decoder_io_sigs_ren2)
                    begin 
                      if (fp_decoder_io_sigs_swap12)
                         begin 
                           ex_ra_0 <=io_inst[24:20];
                         end 
                       else 
                         if (fp_decoder_io_sigs_ren1)
                            begin 
                              if (~fp_decoder_io_sigs_swap12)
                                 begin 
                                   ex_ra_0 <=io_inst[19:15];
                                 end 
                            end 
                    end 
                  else 
                    if (fp_decoder_io_sigs_ren1)
                       begin 
                         if (~fp_decoder_io_sigs_swap12)
                            begin 
                              ex_ra_0 <=io_inst[19:15];
                            end 
                       end 
               end 
         if (metaReset)
            begin 
              ex_ra_1 <=5'h0;
            end 
          else 
            if (io_valid)
               begin 
                 if (fp_decoder_io_sigs_ren2)
                    begin 
                      if (_T_11)
                         begin 
                           ex_ra_1 <=io_inst[24:20];
                         end 
                       else 
                         if (fp_decoder_io_sigs_ren1)
                            begin 
                              if (fp_decoder_io_sigs_swap12)
                                 begin 
                                   ex_ra_1 <=io_inst[19:15];
                                 end 
                            end 
                    end 
                  else 
                    if (fp_decoder_io_sigs_ren1)
                       begin 
                         if (fp_decoder_io_sigs_swap12)
                            begin 
                              ex_ra_1 <=io_inst[19:15];
                            end 
                       end 
               end 
         if (metaReset)
            begin 
              ex_ra_2 <=5'h0;
            end 
          else 
            if (io_valid)
               begin 
                 if (fp_decoder_io_sigs_ren3)
                    begin 
                      ex_ra_2 <=io_inst[31:27];
                    end 
                  else 
                    if (fp_decoder_io_sigs_ren2)
                       begin 
                         if (fp_decoder_io_sigs_swap23)
                            begin 
                              ex_ra_2 <=io_inst[24:20];
                            end 
                       end 
               end 
         if (metaReset)
            begin 
              load_wb <=1'h0;
            end 
          else 
            begin 
              load_wb <=io_dmem_resp_val;
            end 
         if (metaReset)
            begin 
              load_wb_typeTag <=2'h0;
            end 
          else 
            if (io_dmem_resp_val)
               begin 
                 load_wb_typeTag <=_load_wb_typeTag_T_2;
               end 
         if (metaReset)
            begin 
              load_wb_data <=64'h0;
            end 
          else 
            if (io_dmem_resp_val)
               begin 
                 load_wb_data <=io_dmem_resp_data;
               end 
         if (metaReset)
            begin 
              load_wb_tag <=5'h0;
            end 
          else 
            if (io_dmem_resp_val)
               begin 
                 load_wb_tag <=io_dmem_resp_tag;
               end 
         if (metaReset)
            begin 
              mem_reg_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 mem_reg_valid <=1'h0;
               end 
             else 
               begin 
                 mem_reg_valid <=_mem_reg_valid_T_1;
               end 
         if (metaReset)
            begin 
              mem_reg_inst <=32'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_reg_inst <=ex_reg_inst;
               end 
         if (metaReset)
            begin 
              wb_reg_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 wb_reg_valid <=1'h0;
               end 
             else 
               begin 
                 wb_reg_valid <=wb_reg_valid_x7;
               end 
         if (metaReset)
            begin 
              mem_ctrl_typeTagOut <=2'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_typeTagOut <=ex_reg_ctrl_typeTagOut;
               end 
         if (metaReset)
            begin 
              mem_ctrl_fromint <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_fromint <=ex_reg_ctrl_fromint;
               end 
         if (metaReset)
            begin 
              mem_ctrl_toint <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_toint <=ex_reg_ctrl_toint;
               end 
         if (metaReset)
            begin 
              mem_ctrl_fastpipe <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_fastpipe <=ex_reg_ctrl_fastpipe;
               end 
         if (metaReset)
            begin 
              mem_ctrl_fma <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_fma <=ex_reg_ctrl_fma;
               end 
         if (metaReset)
            begin 
              mem_ctrl_div <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_div <=ex_reg_ctrl_div;
               end 
         if (metaReset)
            begin 
              mem_ctrl_sqrt <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_sqrt <=ex_reg_ctrl_sqrt;
               end 
         if (metaReset)
            begin 
              mem_ctrl_wflags <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 mem_ctrl_wflags <=ex_reg_ctrl_wflags;
               end 
         if (metaReset)
            begin 
              wb_ctrl_toint <=1'h0;
            end 
          else 
            if (mem_reg_valid)
               begin 
                 wb_ctrl_toint <=mem_ctrl_toint;
               end 
         if (metaReset)
            begin 
              divSqrt_waddr <=5'h0;
            end 
          else 
            if (divSqrt_inValid)
               begin 
                 divSqrt_waddr <=mem_reg_inst[11:7];
               end 
         if (metaReset)
            begin 
              wen <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 wen <=3'h0;
               end 
             else 
               if (mem_wen)
                  begin 
                    if (~killm)
                       begin 
                         wen <=_wen_T_2;
                       end 
                     else 
                       begin 
                         wen <={1'b0,wen[2:1]};
                       end 
                  end 
                else 
                  begin 
                    wen <={1'b0,wen[2:1]};
                  end 
         if (metaReset)
            begin 
              wbInfo_0_rd <=5'h0;
            end 
          else 
            if (mem_wen)
               begin 
                 if (_T_20)
                    begin 
                      wbInfo_0_rd <=mem_reg_inst[11:7];
                    end 
                  else 
                    if (wen[1])
                       begin 
                         wbInfo_0_rd <=wbInfo_1_rd;
                       end 
               end 
             else 
               if (wen[1])
                  begin 
                    wbInfo_0_rd <=wbInfo_1_rd;
                  end 
         if (metaReset)
            begin 
              wbInfo_0_typeTag <=1'h0;
            end 
          else 
            begin 
              wbInfo_0_typeTag <=_GEN_136[0];
            end 
         if (metaReset)
            begin 
              wbInfo_0_pipeid <=2'h0;
            end 
          else 
            if (mem_wen)
               begin 
                 if (_T_20)
                    begin 
                      wbInfo_0_pipeid <=_wbInfo_0_pipeid_T_10;
                    end 
                  else 
                    if (wen[1])
                       begin 
                         wbInfo_0_pipeid <=wbInfo_1_pipeid;
                       end 
               end 
             else 
               if (wen[1])
                  begin 
                    wbInfo_0_pipeid <=wbInfo_1_pipeid;
                  end 
         if (metaReset)
            begin 
              wbInfo_1_rd <=5'h0;
            end 
          else 
            if (mem_wen)
               begin 
                 if (_T_23)
                    begin 
                      wbInfo_1_rd <=mem_reg_inst[11:7];
                    end 
                  else 
                    if (wen[2])
                       begin 
                         wbInfo_1_rd <=wbInfo_2_rd;
                       end 
               end 
             else 
               if (wen[2])
                  begin 
                    wbInfo_1_rd <=wbInfo_2_rd;
                  end 
         if (metaReset)
            begin 
              wbInfo_1_typeTag <=1'h0;
            end 
          else 
            begin 
              wbInfo_1_typeTag <=_GEN_140[0];
            end 
         if (metaReset)
            begin 
              wbInfo_1_pipeid <=2'h0;
            end 
          else 
            if (mem_wen)
               begin 
                 if (_T_23)
                    begin 
                      wbInfo_1_pipeid <=_wbInfo_0_pipeid_T_10;
                    end 
                  else 
                    if (wen[2])
                       begin 
                         wbInfo_1_pipeid <=wbInfo_2_pipeid;
                       end 
               end 
             else 
               if (wen[2])
                  begin 
                    wbInfo_1_pipeid <=wbInfo_2_pipeid;
                  end 
         if (metaReset)
            begin 
              wbInfo_2_rd <=5'h0;
            end 
          else 
            if (mem_wen)
               begin 
                 if (_T_26)
                    begin 
                      wbInfo_2_rd <=mem_reg_inst[11:7];
                    end 
               end 
         if (metaReset)
            begin 
              wbInfo_2_typeTag <=1'h0;
            end 
          else 
            begin 
              wbInfo_2_typeTag <=_GEN_144[0];
            end 
         if (metaReset)
            begin 
              wbInfo_2_pipeid <=2'h0;
            end 
          else 
            if (mem_wen)
               begin 
                 if (_T_26)
                    begin 
                      wbInfo_2_pipeid <=_wbInfo_0_pipeid_T_10;
                    end 
               end 
         if (metaReset)
            begin 
              write_port_busy <=1'h0;
            end 
          else 
            if (ex_reg_valid)
               begin 
                 write_port_busy <=_write_port_busy_T_27;
               end 
         if (metaReset)
            begin 
              divSqrt_killed <=1'h0;
            end 
          else 
            begin 
              divSqrt_killed <=reset|_divSqrt_killed_T;
            end 
         if (metaReset)
            begin 
              wb_toint_exc <=5'h0;
            end 
          else 
            if (mem_ctrl_toint)
               begin 
                 wb_toint_exc <=fpiu_io_out_bits_exc;
               end 
         if (metaReset)
            begin 
              io_sboard_set_REG <=1'h0;
            end 
          else 
            begin 
              io_sboard_set_REG <=_io_sboard_set_x27_T_3|mem_ctrl_sqrt;
            end 
         if (load_wb&~_T_2)
            begin $display("Assertion failed\n    at FPU.scala:800 assert(consistent(wdata))\n");
            end 
         if (load_wb&~_T_2)
            begin $display("fatal");
            end 
         if (load_wb&~reset)
            begin $display("f%d p%d 0x%x\n",load_wb_tag,_T_5,load_wb_data);
            end 
         if (frfWriteBundle_1_wrenf&~_T_33)
            begin $display("Assertion failed\n    at FPU.scala:938 assert(consistent(wdata))\n");
            end 
         if (frfWriteBundle_1_wrenf&~_T_33)
            begin $display("fatal");
            end 
         if (frfWriteBundle_1_wrenf&~reset)
            begin $display("f%d p%d 0x%x\n",waddr,_T_36,_T_40);
            end 
         FPU_state <=FPU_xor0;
         if (!(FPU_cov_read_data))
            begin 
              FPU_covSum <=FPU_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              FPU_metaAssert <=1'h0;
            end 
          else 
            begin 
              FPU_metaAssert <=FPU_metaAssert|FPU_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (FPU_cov_write_en&FPU_cov_write_mask)
            begin 
              FPU_cov [FPU_cov_write_addr]<=FPU_cov_write_data;
            end 
       end
  
endmodule
 
module HellaCacheArbiter (
  input clock,
  output io_requestor_0_req_ready,
  input io_requestor_0_req_valid,
  input [39:0] io_requestor_0_req_bits_addr,
  input io_requestor_0_s1_kill,
  output io_requestor_0_s2_nack,
  output io_requestor_0_resp_valid,
  output [63:0] io_requestor_0_resp_bits_data,
  output io_requestor_0_s2_xcpt_ae_ld,
  output io_requestor_1_req_ready,
  input io_requestor_1_req_valid,
  input [39:0] io_requestor_1_req_bits_addr,
  input [6:0] io_requestor_1_req_bits_tag,
  input [4:0] io_requestor_1_req_bits_cmd,
  input [1:0] io_requestor_1_req_bits_size,
  input io_requestor_1_req_bits_signed,
  input io_requestor_1_s1_kill,
  input [63:0] io_requestor_1_s1_data_data,
  output io_requestor_1_s2_nack,
  output io_requestor_1_resp_valid,
  output [6:0] io_requestor_1_resp_bits_tag,
  output [1:0] io_requestor_1_resp_bits_size,
  output [63:0] io_requestor_1_resp_bits_data,
  output io_requestor_1_resp_bits_replay,
  output io_requestor_1_resp_bits_has_data,
  output [63:0] io_requestor_1_resp_bits_data_word_bypass,
  output io_requestor_1_replay_next,
  output io_requestor_1_s2_xcpt_ma_ld,
  output io_requestor_1_s2_xcpt_ma_st,
  output io_requestor_1_s2_xcpt_pf_ld,
  output io_requestor_1_s2_xcpt_pf_st,
  output io_requestor_1_s2_xcpt_ae_ld,
  output io_requestor_1_s2_xcpt_ae_st,
  output io_requestor_1_ordered,
  output io_requestor_1_perf_release,
  output io_requestor_1_perf_grant,
  input io_mem_req_ready,
  output io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [6:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [1:0] io_mem_req_bits_size,
  output io_mem_req_bits_signed,
  output io_mem_req_bits_phys,
  output io_mem_s1_kill,
  output [63:0] io_mem_s1_data_data,
  input io_mem_s2_nack,
  input io_mem_resp_valid,
  input [6:0] io_mem_resp_bits_tag,
  input [1:0] io_mem_resp_bits_size,
  input [63:0] io_mem_resp_bits_data,
  input io_mem_resp_bits_replay,
  input io_mem_resp_bits_has_data,
  input [63:0] io_mem_resp_bits_data_word_bypass,
  input io_mem_replay_next,
  input io_mem_s2_xcpt_ma_ld,
  input io_mem_s2_xcpt_ma_st,
  input io_mem_s2_xcpt_pf_ld,
  input io_mem_s2_xcpt_pf_st,
  input io_mem_s2_xcpt_ae_ld,
  input io_mem_s2_xcpt_ae_st,
  input io_mem_ordered,
  input io_mem_perf_release,
  input io_mem_perf_grant,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg s1_id ;  
   reg [31:0] _RAND_0 ;  
   reg s2_id ;  
   reg [31:0] _RAND_1 ;  
   wire [7:0] _io_mem_req_bits_tag_T ;  
   wire [7:0] _GEN_1 ;  
   wire tag_hit ;  
   reg HellaCacheArbiter_state ;  
   reg [31:0] _RAND_2 ;  
   reg HellaCacheArbiter_cov[0:1] ;  
   reg [31:0] _RAND_3 ;  
   wire HellaCacheArbiter_cov_read_data ;  
   wire HellaCacheArbiter_cov_read_addr ;  
   wire HellaCacheArbiter_cov_write_data ;  
   wire HellaCacheArbiter_cov_write_addr ;  
   wire HellaCacheArbiter_cov_write_mask ;  
   wire HellaCacheArbiter_cov_write_en ;  
   reg [29:0] HellaCacheArbiter_covSum ;  
   reg [31:0] _RAND_4 ;  
   wire s1_id_shl ;  
   wire s1_id_pad ;  
  assign _io_mem_req_bits_tag_T={io_requestor_1_req_bits_tag,1'h1}; 
  assign _GEN_1=io_requestor_0_req_valid ? 8'h0:_io_mem_req_bits_tag_T; 
  assign tag_hit=~io_mem_resp_bits_tag[0]; 
  assign io_requestor_0_req_ready=io_mem_req_ready; 
  assign io_requestor_0_s2_nack=io_mem_s2_nack&~s2_id; 
  assign io_requestor_0_resp_valid=io_mem_resp_valid&tag_hit; 
  assign io_requestor_0_resp_bits_data=io_mem_resp_bits_data; 
  assign io_requestor_0_s2_xcpt_ae_ld=io_mem_s2_xcpt_ae_ld; 
  assign io_requestor_1_req_ready=io_requestor_0_req_ready&~io_requestor_0_req_valid; 
  assign io_requestor_1_s2_nack=io_mem_s2_nack&s2_id; 
  assign io_requestor_1_resp_valid=io_mem_resp_valid&io_mem_resp_bits_tag[0]; 
  assign io_requestor_1_resp_bits_tag={1'b0,io_mem_resp_bits_tag[6:1]}; 
  assign io_requestor_1_resp_bits_size=io_mem_resp_bits_size; 
  assign io_requestor_1_resp_bits_data=io_mem_resp_bits_data; 
  assign io_requestor_1_resp_bits_replay=io_mem_resp_bits_replay; 
  assign io_requestor_1_resp_bits_has_data=io_mem_resp_bits_has_data; 
  assign io_requestor_1_resp_bits_data_word_bypass=io_mem_resp_bits_data_word_bypass; 
  assign io_requestor_1_replay_next=io_mem_replay_next; 
  assign io_requestor_1_s2_xcpt_ma_ld=io_mem_s2_xcpt_ma_ld; 
  assign io_requestor_1_s2_xcpt_ma_st=io_mem_s2_xcpt_ma_st; 
  assign io_requestor_1_s2_xcpt_pf_ld=io_mem_s2_xcpt_pf_ld; 
  assign io_requestor_1_s2_xcpt_pf_st=io_mem_s2_xcpt_pf_st; 
  assign io_requestor_1_s2_xcpt_ae_ld=io_mem_s2_xcpt_ae_ld; 
  assign io_requestor_1_s2_xcpt_ae_st=io_mem_s2_xcpt_ae_st; 
  assign io_requestor_1_ordered=io_mem_ordered; 
  assign io_requestor_1_perf_release=io_mem_perf_release; 
  assign io_requestor_1_perf_grant=io_mem_perf_grant; 
  assign io_mem_req_valid=io_requestor_0_req_valid|io_requestor_1_req_valid; 
  assign io_mem_req_bits_addr=io_requestor_0_req_valid ? io_requestor_0_req_bits_addr:io_requestor_1_req_bits_addr; 
  assign io_mem_req_bits_tag=_GEN_1[6:0]; 
  assign io_mem_req_bits_cmd=io_requestor_0_req_valid ? 5'h0:io_requestor_1_req_bits_cmd; 
  assign io_mem_req_bits_size=io_requestor_0_req_valid ? 2'h3:io_requestor_1_req_bits_size; 
  assign io_mem_req_bits_signed=io_requestor_0_req_valid ? 1'h0:io_requestor_1_req_bits_signed; 
  assign io_mem_req_bits_phys=io_requestor_0_req_valid; 
  assign io_mem_s1_kill=s1_id ? io_requestor_1_s1_kill:io_requestor_0_s1_kill; 
  assign io_mem_s1_data_data=s1_id ? io_requestor_1_s1_data_data:64'h0; 
  assign HellaCacheArbiter_cov_read_addr=HellaCacheArbiter_state; 
  assign HellaCacheArbiter_cov_read_data=HellaCacheArbiter_cov[HellaCacheArbiter_cov_read_addr]; 
  assign HellaCacheArbiter_cov_write_data=1'h1; 
  assign HellaCacheArbiter_cov_write_addr=HellaCacheArbiter_state; 
  assign HellaCacheArbiter_cov_write_mask=1'h1; 
  assign HellaCacheArbiter_cov_write_en=1'h1; 
  assign s1_id_shl=s1_id; 
  assign s1_id_pad=s1_id_shl; 
  assign io_covSum=HellaCacheArbiter_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              s1_id <=1'h0;
            end 
          else 
            if (io_requestor_0_req_valid)
               begin 
                 s1_id <=1'h0;
               end 
             else 
               begin 
                 s1_id <=1'h1;
               end 
         if (metaReset)
            begin 
              s2_id <=1'h0;
            end 
          else 
            begin 
              s2_id <=s1_id;
            end 
         HellaCacheArbiter_state <=s1_id_pad;
         if (!(HellaCacheArbiter_cov_read_data))
            begin 
              HellaCacheArbiter_covSum <=HellaCacheArbiter_covSum+1'h1;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (HellaCacheArbiter_cov_write_en&HellaCacheArbiter_cov_write_mask)
            begin 
              HellaCacheArbiter_cov [HellaCacheArbiter_cov_write_addr]<=HellaCacheArbiter_cov_write_data;
            end 
       end
  
endmodule
 
module PTW (
  input clock,
  input reset,
  output io_requestor_0_req_ready,
  input io_requestor_0_req_valid,
  input [26:0] io_requestor_0_req_bits_bits_addr,
  output io_requestor_0_resp_valid,
  output io_requestor_0_resp_bits_ae,
  output [53:0] io_requestor_0_resp_bits_pte_ppn,
  output io_requestor_0_resp_bits_pte_d,
  output io_requestor_0_resp_bits_pte_a,
  output io_requestor_0_resp_bits_pte_g,
  output io_requestor_0_resp_bits_pte_u,
  output io_requestor_0_resp_bits_pte_x,
  output io_requestor_0_resp_bits_pte_w,
  output io_requestor_0_resp_bits_pte_r,
  output io_requestor_0_resp_bits_pte_v,
  output [1:0] io_requestor_0_resp_bits_level,
  output io_requestor_0_resp_bits_homogeneous,
  output [3:0] io_requestor_0_ptbr_mode,
  output io_requestor_0_status_debug,
  output [1:0] io_requestor_0_status_dprv,
  output io_requestor_0_status_mxr,
  output io_requestor_0_status_sum,
  output io_requestor_0_pmp_0_cfg_l,
  output [1:0] io_requestor_0_pmp_0_cfg_a,
  output io_requestor_0_pmp_0_cfg_x,
  output io_requestor_0_pmp_0_cfg_w,
  output io_requestor_0_pmp_0_cfg_r,
  output [29:0] io_requestor_0_pmp_0_addr,
  output [31:0] io_requestor_0_pmp_0_mask,
  output io_requestor_0_pmp_1_cfg_l,
  output [1:0] io_requestor_0_pmp_1_cfg_a,
  output io_requestor_0_pmp_1_cfg_x,
  output io_requestor_0_pmp_1_cfg_w,
  output io_requestor_0_pmp_1_cfg_r,
  output [29:0] io_requestor_0_pmp_1_addr,
  output [31:0] io_requestor_0_pmp_1_mask,
  output io_requestor_0_pmp_2_cfg_l,
  output [1:0] io_requestor_0_pmp_2_cfg_a,
  output io_requestor_0_pmp_2_cfg_x,
  output io_requestor_0_pmp_2_cfg_w,
  output io_requestor_0_pmp_2_cfg_r,
  output [29:0] io_requestor_0_pmp_2_addr,
  output [31:0] io_requestor_0_pmp_2_mask,
  output io_requestor_0_pmp_3_cfg_l,
  output [1:0] io_requestor_0_pmp_3_cfg_a,
  output io_requestor_0_pmp_3_cfg_x,
  output io_requestor_0_pmp_3_cfg_w,
  output io_requestor_0_pmp_3_cfg_r,
  output [29:0] io_requestor_0_pmp_3_addr,
  output [31:0] io_requestor_0_pmp_3_mask,
  output io_requestor_0_pmp_4_cfg_l,
  output [1:0] io_requestor_0_pmp_4_cfg_a,
  output io_requestor_0_pmp_4_cfg_x,
  output io_requestor_0_pmp_4_cfg_w,
  output io_requestor_0_pmp_4_cfg_r,
  output [29:0] io_requestor_0_pmp_4_addr,
  output [31:0] io_requestor_0_pmp_4_mask,
  output io_requestor_0_pmp_5_cfg_l,
  output [1:0] io_requestor_0_pmp_5_cfg_a,
  output io_requestor_0_pmp_5_cfg_x,
  output io_requestor_0_pmp_5_cfg_w,
  output io_requestor_0_pmp_5_cfg_r,
  output [29:0] io_requestor_0_pmp_5_addr,
  output [31:0] io_requestor_0_pmp_5_mask,
  output io_requestor_0_pmp_6_cfg_l,
  output [1:0] io_requestor_0_pmp_6_cfg_a,
  output io_requestor_0_pmp_6_cfg_x,
  output io_requestor_0_pmp_6_cfg_w,
  output io_requestor_0_pmp_6_cfg_r,
  output [29:0] io_requestor_0_pmp_6_addr,
  output [31:0] io_requestor_0_pmp_6_mask,
  output io_requestor_0_pmp_7_cfg_l,
  output [1:0] io_requestor_0_pmp_7_cfg_a,
  output io_requestor_0_pmp_7_cfg_x,
  output io_requestor_0_pmp_7_cfg_w,
  output io_requestor_0_pmp_7_cfg_r,
  output [29:0] io_requestor_0_pmp_7_addr,
  output [31:0] io_requestor_0_pmp_7_mask,
  output io_requestor_1_req_ready,
  input io_requestor_1_req_valid,
  input io_requestor_1_req_bits_valid,
  input [26:0] io_requestor_1_req_bits_bits_addr,
  output io_requestor_1_resp_valid,
  output io_requestor_1_resp_bits_ae,
  output [53:0] io_requestor_1_resp_bits_pte_ppn,
  output io_requestor_1_resp_bits_pte_d,
  output io_requestor_1_resp_bits_pte_a,
  output io_requestor_1_resp_bits_pte_g,
  output io_requestor_1_resp_bits_pte_u,
  output io_requestor_1_resp_bits_pte_x,
  output io_requestor_1_resp_bits_pte_w,
  output io_requestor_1_resp_bits_pte_r,
  output io_requestor_1_resp_bits_pte_v,
  output [1:0] io_requestor_1_resp_bits_level,
  output io_requestor_1_resp_bits_homogeneous,
  output [3:0] io_requestor_1_ptbr_mode,
  output io_requestor_1_status_debug,
  output [1:0] io_requestor_1_status_prv,
  output io_requestor_1_pmp_0_cfg_l,
  output [1:0] io_requestor_1_pmp_0_cfg_a,
  output io_requestor_1_pmp_0_cfg_x,
  output io_requestor_1_pmp_0_cfg_w,
  output io_requestor_1_pmp_0_cfg_r,
  output [29:0] io_requestor_1_pmp_0_addr,
  output [31:0] io_requestor_1_pmp_0_mask,
  output io_requestor_1_pmp_1_cfg_l,
  output [1:0] io_requestor_1_pmp_1_cfg_a,
  output io_requestor_1_pmp_1_cfg_x,
  output io_requestor_1_pmp_1_cfg_w,
  output io_requestor_1_pmp_1_cfg_r,
  output [29:0] io_requestor_1_pmp_1_addr,
  output [31:0] io_requestor_1_pmp_1_mask,
  output io_requestor_1_pmp_2_cfg_l,
  output [1:0] io_requestor_1_pmp_2_cfg_a,
  output io_requestor_1_pmp_2_cfg_x,
  output io_requestor_1_pmp_2_cfg_w,
  output io_requestor_1_pmp_2_cfg_r,
  output [29:0] io_requestor_1_pmp_2_addr,
  output [31:0] io_requestor_1_pmp_2_mask,
  output io_requestor_1_pmp_3_cfg_l,
  output [1:0] io_requestor_1_pmp_3_cfg_a,
  output io_requestor_1_pmp_3_cfg_x,
  output io_requestor_1_pmp_3_cfg_w,
  output io_requestor_1_pmp_3_cfg_r,
  output [29:0] io_requestor_1_pmp_3_addr,
  output [31:0] io_requestor_1_pmp_3_mask,
  output io_requestor_1_pmp_4_cfg_l,
  output [1:0] io_requestor_1_pmp_4_cfg_a,
  output io_requestor_1_pmp_4_cfg_x,
  output io_requestor_1_pmp_4_cfg_w,
  output io_requestor_1_pmp_4_cfg_r,
  output [29:0] io_requestor_1_pmp_4_addr,
  output [31:0] io_requestor_1_pmp_4_mask,
  output io_requestor_1_pmp_5_cfg_l,
  output [1:0] io_requestor_1_pmp_5_cfg_a,
  output io_requestor_1_pmp_5_cfg_x,
  output io_requestor_1_pmp_5_cfg_w,
  output io_requestor_1_pmp_5_cfg_r,
  output [29:0] io_requestor_1_pmp_5_addr,
  output [31:0] io_requestor_1_pmp_5_mask,
  output io_requestor_1_pmp_6_cfg_l,
  output [1:0] io_requestor_1_pmp_6_cfg_a,
  output io_requestor_1_pmp_6_cfg_x,
  output io_requestor_1_pmp_6_cfg_w,
  output io_requestor_1_pmp_6_cfg_r,
  output [29:0] io_requestor_1_pmp_6_addr,
  output [31:0] io_requestor_1_pmp_6_mask,
  output io_requestor_1_pmp_7_cfg_l,
  output [1:0] io_requestor_1_pmp_7_cfg_a,
  output io_requestor_1_pmp_7_cfg_x,
  output io_requestor_1_pmp_7_cfg_w,
  output io_requestor_1_pmp_7_cfg_r,
  output [29:0] io_requestor_1_pmp_7_addr,
  output [31:0] io_requestor_1_pmp_7_mask,
  output [63:0] io_requestor_1_customCSRs_csrs_0_value,
  input io_mem_req_ready,
  output io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output io_mem_s1_kill,
  input io_mem_s2_nack,
  input io_mem_resp_valid,
  input [63:0] io_mem_resp_bits_data,
  input io_mem_s2_xcpt_ae_ld,
  input [3:0] io_dpath_ptbr_mode,
  input [43:0] io_dpath_ptbr_ppn,
  input io_dpath_sfence_valid,
  input io_dpath_sfence_bits_rs1,
  input io_dpath_status_debug,
  input [1:0] io_dpath_status_dprv,
  input [1:0] io_dpath_status_prv,
  input io_dpath_status_mxr,
  input io_dpath_status_sum,
  input io_dpath_pmp_0_cfg_l,
  input [1:0] io_dpath_pmp_0_cfg_a,
  input io_dpath_pmp_0_cfg_x,
  input io_dpath_pmp_0_cfg_w,
  input io_dpath_pmp_0_cfg_r,
  input [29:0] io_dpath_pmp_0_addr,
  input [31:0] io_dpath_pmp_0_mask,
  input io_dpath_pmp_1_cfg_l,
  input [1:0] io_dpath_pmp_1_cfg_a,
  input io_dpath_pmp_1_cfg_x,
  input io_dpath_pmp_1_cfg_w,
  input io_dpath_pmp_1_cfg_r,
  input [29:0] io_dpath_pmp_1_addr,
  input [31:0] io_dpath_pmp_1_mask,
  input io_dpath_pmp_2_cfg_l,
  input [1:0] io_dpath_pmp_2_cfg_a,
  input io_dpath_pmp_2_cfg_x,
  input io_dpath_pmp_2_cfg_w,
  input io_dpath_pmp_2_cfg_r,
  input [29:0] io_dpath_pmp_2_addr,
  input [31:0] io_dpath_pmp_2_mask,
  input io_dpath_pmp_3_cfg_l,
  input [1:0] io_dpath_pmp_3_cfg_a,
  input io_dpath_pmp_3_cfg_x,
  input io_dpath_pmp_3_cfg_w,
  input io_dpath_pmp_3_cfg_r,
  input [29:0] io_dpath_pmp_3_addr,
  input [31:0] io_dpath_pmp_3_mask,
  input io_dpath_pmp_4_cfg_l,
  input [1:0] io_dpath_pmp_4_cfg_a,
  input io_dpath_pmp_4_cfg_x,
  input io_dpath_pmp_4_cfg_w,
  input io_dpath_pmp_4_cfg_r,
  input [29:0] io_dpath_pmp_4_addr,
  input [31:0] io_dpath_pmp_4_mask,
  input io_dpath_pmp_5_cfg_l,
  input [1:0] io_dpath_pmp_5_cfg_a,
  input io_dpath_pmp_5_cfg_x,
  input io_dpath_pmp_5_cfg_w,
  input io_dpath_pmp_5_cfg_r,
  input [29:0] io_dpath_pmp_5_addr,
  input [31:0] io_dpath_pmp_5_mask,
  input io_dpath_pmp_6_cfg_l,
  input [1:0] io_dpath_pmp_6_cfg_a,
  input io_dpath_pmp_6_cfg_x,
  input io_dpath_pmp_6_cfg_w,
  input io_dpath_pmp_6_cfg_r,
  input [29:0] io_dpath_pmp_6_addr,
  input [31:0] io_dpath_pmp_6_mask,
  input io_dpath_pmp_7_cfg_l,
  input [1:0] io_dpath_pmp_7_cfg_a,
  input io_dpath_pmp_7_cfg_x,
  input io_dpath_pmp_7_cfg_w,
  input io_dpath_pmp_7_cfg_r,
  input [29:0] io_dpath_pmp_7_addr,
  input [31:0] io_dpath_pmp_7_mask,
  output io_dpath_perf_l2hit,
  output io_dpath_perf_pte_miss,
  output io_dpath_perf_pte_hit,
  input [63:0] io_dpath_customCSRs_csrs_0_value,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire arb_io_in_0_ready ;  
   wire arb_io_in_0_valid ;  
   wire [26:0] arb_io_in_0_bits_bits_addr ;  
   wire arb_io_in_1_ready ;  
   wire arb_io_in_1_valid ;  
   wire arb_io_in_1_bits_valid ;  
   wire [26:0] arb_io_in_1_bits_bits_addr ;  
   wire arb_io_out_ready ;  
   wire arb_io_out_valid ;  
   wire arb_io_out_bits_valid ;  
   wire [26:0] arb_io_out_bits_bits_addr ;  
   wire arb_io_chosen ;  
   wire [29:0] arb_io_covSum ;  
   wire arb_metaAssert ;  
   wire [2:0] state_barrier_io_x ;  
   wire [2:0] state_barrier_io_y ;  
   wire [29:0] state_barrier_io_covSum ;  
   wire state_barrier_metaAssert ;  
   wire [53:0] r_pte_barrier_io_x_ppn ;  
   wire r_pte_barrier_io_x_d ;  
   wire r_pte_barrier_io_x_a ;  
   wire r_pte_barrier_io_x_g ;  
   wire r_pte_barrier_io_x_u ;  
   wire r_pte_barrier_io_x_x ;  
   wire r_pte_barrier_io_x_w ;  
   wire r_pte_barrier_io_x_r ;  
   wire r_pte_barrier_io_x_v ;  
   wire [53:0] r_pte_barrier_io_y_ppn ;  
   wire r_pte_barrier_io_y_d ;  
   wire r_pte_barrier_io_y_a ;  
   wire r_pte_barrier_io_y_g ;  
   wire r_pte_barrier_io_y_u ;  
   wire r_pte_barrier_io_y_x ;  
   wire r_pte_barrier_io_y_w ;  
   wire r_pte_barrier_io_y_r ;  
   wire r_pte_barrier_io_y_v ;  
   wire [29:0] r_pte_barrier_io_covSum ;  
   wire r_pte_barrier_metaAssert ;  
   reg [2:0] state ;  
   reg [31:0] _RAND_0 ;  
   wire _arb_io_out_ready_T ;  
   reg l2_refill ;  
   reg [31:0] _RAND_1 ;  
   reg resp_valid_0 ;  
   reg [31:0] _RAND_2 ;  
   reg resp_valid_1 ;  
   reg [31:0] _RAND_3 ;  
   wire _clock_en_T ;  
   reg invalidated ;  
   reg [31:0] _RAND_4 ;  
   reg [1:0] count ;  
   reg [31:0] _RAND_5 ;  
   reg resp_ae ;  
   reg [31:0] _RAND_6 ;  
   reg [26:0] r_req_addr ;  
   reg [31:0] _RAND_7 ;  
   reg r_req_dest ;  
   reg [31:0] _RAND_8 ;  
   reg [53:0] r_pte_ppn ;  
   reg [63:0] _RAND_9 ;  
   reg r_pte_d ;  
   reg [31:0] _RAND_10 ;  
   reg r_pte_a ;  
   reg [31:0] _RAND_11 ;  
   reg r_pte_g ;  
   reg [31:0] _RAND_12 ;  
   reg r_pte_u ;  
   reg [31:0] _RAND_13 ;  
   reg r_pte_x ;  
   reg [31:0] _RAND_14 ;  
   reg r_pte_w ;  
   reg [31:0] _RAND_15 ;  
   reg r_pte_r ;  
   reg [31:0] _RAND_16 ;  
   reg r_pte_v ;  
   reg [31:0] _RAND_17 ;  
   reg mem_resp_valid ;  
   reg [31:0] _RAND_18 ;  
   reg [63:0] mem_resp_data ;  
   reg [63:0] _RAND_19 ;  
   wire tmp_v ;  
   wire tmp_r ;  
   wire tmp_w ;  
   wire tmp_x ;  
   wire tmp_u ;  
   wire tmp_g ;  
   wire tmp_a ;  
   wire tmp_d ;  
   wire [53:0] tmp_ppn ;  
   wire _T_11 ;  
   wire _T_12 ;  
   wire _T_13 ;  
   wire _T_15 ;  
   wire _T_16 ;  
   wire _GEN_0 ;  
   wire _T_17 ;  
   wire _T_19 ;  
   wire _T_20 ;  
   wire _GEN_1 ;  
   wire res_v ;  
   wire invalid_paddr ;  
   wire _traverse_T_1 ;  
   wire _traverse_T_3 ;  
   wire _traverse_T_5 ;  
   wire _traverse_T_7 ;  
   wire _traverse_T_8 ;  
   wire traverse ;  
   wire [8:0] vpn_idxs_0 ;  
   wire [8:0] vpn_idxs_1 ;  
   wire [8:0] vpn_idxs_2 ;  
   wire _pte_addr_vpn_idx_T ;  
   wire [8:0] _pte_addr_vpn_idx_T_1 ;  
   wire _pte_addr_vpn_idx_T_2 ;  
   wire [8:0] _pte_addr_vpn_idx_T_3 ;  
   wire _pte_addr_vpn_idx_T_4 ;  
   wire [8:0] vpn_idx ;  
   wire [62:0] _pte_addr_T ;  
   wire [65:0] pte_addr ;  
   wire [35:0] fragmented_superpage_ppn_choices_hi ;  
   wire [17:0] fragmented_superpage_ppn_choices_lo ;  
   wire [53:0] choices_0 ;  
   wire [44:0] fragmented_superpage_ppn_choices_hi_1 ;  
   wire [53:0] choices_1 ;  
   wire fragmented_superpage_ppn_truncIdx ;  
   wire [53:0] fragmented_superpage_ppn ;  
   wire _T_22 ;  
   reg [6:0] state_reg ;  
   reg [31:0] _RAND_20 ;  
   reg [7:0] valid ;  
   reg [31:0] _RAND_21 ;  
   reg [31:0] tags_0 ;  
   reg [31:0] _RAND_22 ;  
   reg [31:0] tags_1 ;  
   reg [31:0] _RAND_23 ;  
   reg [31:0] tags_2 ;  
   reg [31:0] _RAND_24 ;  
   reg [31:0] tags_3 ;  
   reg [31:0] _RAND_25 ;  
   reg [31:0] tags_4 ;  
   reg [31:0] _RAND_26 ;  
   reg [31:0] tags_5 ;  
   reg [31:0] _RAND_27 ;  
   reg [31:0] tags_6 ;  
   reg [31:0] _RAND_28 ;  
   reg [31:0] tags_7 ;  
   reg [31:0] _RAND_29 ;  
   reg [19:0] data_0 ;  
   reg [31:0] _RAND_30 ;  
   reg [19:0] data_1 ;  
   reg [31:0] _RAND_31 ;  
   reg [19:0] data_2 ;  
   reg [31:0] _RAND_32 ;  
   reg [19:0] data_3 ;  
   reg [31:0] _RAND_33 ;  
   reg [19:0] data_4 ;  
   reg [31:0] _RAND_34 ;  
   reg [19:0] data_5 ;  
   reg [31:0] _RAND_35 ;  
   reg [19:0] data_6 ;  
   reg [31:0] _RAND_36 ;  
   reg [19:0] data_7 ;  
   reg [31:0] _RAND_37 ;  
   wire [65:0] _GEN_115 ;  
   wire lo_lo_lo ;  
   wire [65:0] _GEN_116 ;  
   wire lo_lo_hi ;  
   wire [65:0] _GEN_117 ;  
   wire lo_hi_lo ;  
   wire [65:0] _GEN_118 ;  
   wire lo_hi_hi ;  
   wire [65:0] _GEN_119 ;  
   wire hi_lo_lo ;  
   wire [65:0] _GEN_120 ;  
   wire hi_lo_hi ;  
   wire [65:0] _GEN_121 ;  
   wire hi_hi_lo ;  
   wire [65:0] _GEN_122 ;  
   wire hi_hi_hi ;  
   wire [7:0] _T_23 ;  
   wire [7:0] hits ;  
   wire hit ;  
   wire _T_24 ;  
   wire _T_26 ;  
   wire _T_28 ;  
   wire _T_29 ;  
   wire hi_1 ;  
   wire [2:0] left_subtree_state ;  
   wire [2:0] right_subtree_state ;  
   wire hi_2 ;  
   wire left_subtree_state_1 ;  
   wire right_subtree_state_1 ;  
   wire lo_1 ;  
   wire [1:0] _T_32 ;  
   wire hi_3 ;  
   wire left_subtree_state_2 ;  
   wire right_subtree_state_2 ;  
   wire lo_2 ;  
   wire [1:0] _T_35 ;  
   wire [1:0] lo_3 ;  
   wire [2:0] _T_36 ;  
   wire _T_38 ;  
   wire _T_39 ;  
   wire _T_40 ;  
   wire _T_41 ;  
   wire _T_42 ;  
   wire _T_43 ;  
   wire _T_44 ;  
   wire [2:0] _T_46 ;  
   wire [2:0] _T_47 ;  
   wire [2:0] _T_48 ;  
   wire [2:0] _T_49 ;  
   wire [2:0] _T_50 ;  
   wire [2:0] _T_51 ;  
   wire [2:0] _T_52 ;  
   wire [2:0] r ;  
   wire [7:0] _T_53 ;  
   wire [7:0] _T_54 ;  
   wire [53:0] res_ppn ;  
   wire _T_55 ;  
   wire _T_56 ;  
   wire [3:0] hi_4 ;  
   wire [3:0] lo_4 ;  
   wire hi_5 ;  
   wire [3:0] _T_57 ;  
   wire [1:0] hi_6 ;  
   wire [1:0] lo_5 ;  
   wire hi_7 ;  
   wire [1:0] _T_58 ;  
   wire lo_6 ;  
   wire [2:0] state_reg_touch_way_sized ;  
   wire state_reg_hi_hi ;  
   wire state_reg_hi_hi_1 ;  
   wire state_reg_hi_lo ;  
   wire state_reg_lo ;  
   wire [2:0] _state_reg_T_7 ;  
   wire [2:0] state_reg_hi_lo_1 ;  
   wire state_reg_hi_lo_2 ;  
   wire state_reg_lo_1 ;  
   wire [2:0] _state_reg_T_15 ;  
   wire [2:0] state_reg_lo_2 ;  
   wire [6:0] _state_reg_T_16 ;  
   wire _T_61 ;  
   wire pte_cache_hit ;  
   wire [19:0] _T_79 ;  
   wire [19:0] _T_80 ;  
   wire [19:0] _T_81 ;  
   wire [19:0] _T_82 ;  
   wire [19:0] _T_83 ;  
   wire [19:0] _T_84 ;  
   wire [19:0] _T_85 ;  
   wire [19:0] _T_86 ;  
   wire [19:0] _T_87 ;  
   wire [19:0] _T_88 ;  
   wire [19:0] _T_89 ;  
   wire [19:0] _T_90 ;  
   wire [19:0] _T_91 ;  
   wire [19:0] _T_92 ;  
   wire [19:0] pte_cache_data ;  
   reg pte_hit ;  
   reg [31:0] _RAND_38 ;  
   wire _io_dpath_perf_pte_hit_T_1 ;  
   wire _T_94 ;  
   wire _T_95 ;  
   wire _T_98 ;  
   wire _invalidated_T_1 ;  
   wire _io_mem_req_valid_T_1 ;  
   wire [65:0] _pmaPgLevelHomogeneous_T_6 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_7 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_9 ;  
   wire _pmaPgLevelHomogeneous_T_10 ;  
   wire [65:0] _pmaPgLevelHomogeneous_T_11 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_12 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_14 ;  
   wire _pmaPgLevelHomogeneous_T_15 ;  
   wire [65:0] _pmaPgLevelHomogeneous_T_16 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_17 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_19 ;  
   wire _pmaPgLevelHomogeneous_T_20 ;  
   wire _pmaPgLevelHomogeneous_T_22 ;  
   wire pmaPgLevelHomogeneous_1 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_26 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_53 ;  
   wire _pmaPgLevelHomogeneous_T_54 ;  
   wire [65:0] _pmaPgLevelHomogeneous_T_55 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_56 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_58 ;  
   wire _pmaPgLevelHomogeneous_T_59 ;  
   wire [65:0] _pmaPgLevelHomogeneous_T_60 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_61 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_63 ;  
   wire _pmaPgLevelHomogeneous_T_64 ;  
   wire [65:0] _pmaPgLevelHomogeneous_T_65 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_66 ;  
   wire [66:0] _pmaPgLevelHomogeneous_T_68 ;  
   wire _pmaPgLevelHomogeneous_T_69 ;  
   wire _pmaPgLevelHomogeneous_T_86 ;  
   wire _pmaPgLevelHomogeneous_T_87 ;  
   wire _pmaPgLevelHomogeneous_T_88 ;  
   wire _pmaPgLevelHomogeneous_T_89 ;  
   wire _pmaPgLevelHomogeneous_T_90 ;  
   wire pmaPgLevelHomogeneous_2 ;  
   wire _pmaHomogeneous_T_1 ;  
   wire _pmaHomogeneous_T_3 ;  
   wire pmaHomogeneous ;  
   wire [65:0] _pmpHomogeneous_T_1 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_4 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_6 ;  
   wire pmpHomogeneous_maskHomogeneous ;  
   wire [31:0] _pmpHomogeneous_T_3 ;  
   wire [31:0] _pmpHomogeneous_T_5 ;  
   wire [65:0] _GEN_123 ;  
   wire [65:0] _pmpHomogeneous_T_7 ;  
   wire _pmpHomogeneous_T_9 ;  
   wire _pmpHomogeneous_T_16 ;  
   wire _pmpHomogeneous_T_23 ;  
   wire _pmpHomogeneous_T_25 ;  
   wire _pmpHomogeneous_T_27 ;  
   wire _pmpHomogeneous_T_29 ;  
   wire _pmpHomogeneous_T_30 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_4 ;  
   wire pmpHomogeneous_beginsAfterUpper ;  
   wire [31:0] _pmpHomogeneous_pgMask_T_1 ;  
   wire [31:0] _pmpHomogeneous_pgMask_T_3 ;  
   wire [31:0] pmpHomogeneous_pgMask ;  
   wire [65:0] _GEN_127 ;  
   wire [65:0] _pmpHomogeneous_endsBeforeLower_T ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_5 ;  
   wire [65:0] _GEN_129 ;  
   wire pmpHomogeneous_endsBeforeUpper ;  
   wire _pmpHomogeneous_T_35 ;  
   wire _pmpHomogeneous_T_36 ;  
   wire _pmpHomogeneous_T_37 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_12 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_14 ;  
   wire pmpHomogeneous_maskHomogeneous_1 ;  
   wire [31:0] _pmpHomogeneous_T_40 ;  
   wire [31:0] _pmpHomogeneous_T_42 ;  
   wire [65:0] _GEN_130 ;  
   wire [65:0] _pmpHomogeneous_T_44 ;  
   wire _pmpHomogeneous_T_46 ;  
   wire _pmpHomogeneous_T_53 ;  
   wire _pmpHomogeneous_T_60 ;  
   wire _pmpHomogeneous_T_62 ;  
   wire _pmpHomogeneous_T_64 ;  
   wire _pmpHomogeneous_T_66 ;  
   wire _pmpHomogeneous_T_67 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_9 ;  
   wire pmpHomogeneous_beginsAfterUpper_1 ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_11 ;  
   wire [65:0] _GEN_138 ;  
   wire pmpHomogeneous_endsBeforeUpper_1 ;  
   wire _pmpHomogeneous_T_70 ;  
   wire _pmpHomogeneous_T_71 ;  
   wire _pmpHomogeneous_T_72 ;  
   wire _pmpHomogeneous_T_73 ;  
   wire _pmpHomogeneous_T_74 ;  
   wire _pmpHomogeneous_T_75 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_20 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_22 ;  
   wire pmpHomogeneous_maskHomogeneous_2 ;  
   wire [31:0] _pmpHomogeneous_T_77 ;  
   wire [31:0] _pmpHomogeneous_T_79 ;  
   wire [65:0] _GEN_139 ;  
   wire [65:0] _pmpHomogeneous_T_81 ;  
   wire _pmpHomogeneous_T_83 ;  
   wire _pmpHomogeneous_T_90 ;  
   wire _pmpHomogeneous_T_97 ;  
   wire _pmpHomogeneous_T_99 ;  
   wire _pmpHomogeneous_T_101 ;  
   wire _pmpHomogeneous_T_103 ;  
   wire _pmpHomogeneous_T_104 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_14 ;  
   wire pmpHomogeneous_beginsAfterUpper_2 ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_17 ;  
   wire [65:0] _GEN_147 ;  
   wire pmpHomogeneous_endsBeforeUpper_2 ;  
   wire _pmpHomogeneous_T_107 ;  
   wire _pmpHomogeneous_T_108 ;  
   wire _pmpHomogeneous_T_109 ;  
   wire _pmpHomogeneous_T_110 ;  
   wire _pmpHomogeneous_T_111 ;  
   wire _pmpHomogeneous_T_112 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_28 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_30 ;  
   wire pmpHomogeneous_maskHomogeneous_3 ;  
   wire [31:0] _pmpHomogeneous_T_114 ;  
   wire [31:0] _pmpHomogeneous_T_116 ;  
   wire [65:0] _GEN_148 ;  
   wire [65:0] _pmpHomogeneous_T_118 ;  
   wire _pmpHomogeneous_T_120 ;  
   wire _pmpHomogeneous_T_127 ;  
   wire _pmpHomogeneous_T_134 ;  
   wire _pmpHomogeneous_T_136 ;  
   wire _pmpHomogeneous_T_138 ;  
   wire _pmpHomogeneous_T_140 ;  
   wire _pmpHomogeneous_T_141 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_19 ;  
   wire pmpHomogeneous_beginsAfterUpper_3 ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_23 ;  
   wire [65:0] _GEN_156 ;  
   wire pmpHomogeneous_endsBeforeUpper_3 ;  
   wire _pmpHomogeneous_T_144 ;  
   wire _pmpHomogeneous_T_145 ;  
   wire _pmpHomogeneous_T_146 ;  
   wire _pmpHomogeneous_T_147 ;  
   wire _pmpHomogeneous_T_148 ;  
   wire _pmpHomogeneous_T_149 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_36 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_38 ;  
   wire pmpHomogeneous_maskHomogeneous_4 ;  
   wire [31:0] _pmpHomogeneous_T_151 ;  
   wire [31:0] _pmpHomogeneous_T_153 ;  
   wire [65:0] _GEN_157 ;  
   wire [65:0] _pmpHomogeneous_T_155 ;  
   wire _pmpHomogeneous_T_157 ;  
   wire _pmpHomogeneous_T_164 ;  
   wire _pmpHomogeneous_T_171 ;  
   wire _pmpHomogeneous_T_173 ;  
   wire _pmpHomogeneous_T_175 ;  
   wire _pmpHomogeneous_T_177 ;  
   wire _pmpHomogeneous_T_178 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_24 ;  
   wire pmpHomogeneous_beginsAfterUpper_4 ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_29 ;  
   wire [65:0] _GEN_165 ;  
   wire pmpHomogeneous_endsBeforeUpper_4 ;  
   wire _pmpHomogeneous_T_181 ;  
   wire _pmpHomogeneous_T_182 ;  
   wire _pmpHomogeneous_T_183 ;  
   wire _pmpHomogeneous_T_184 ;  
   wire _pmpHomogeneous_T_185 ;  
   wire _pmpHomogeneous_T_186 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_44 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_46 ;  
   wire pmpHomogeneous_maskHomogeneous_5 ;  
   wire [31:0] _pmpHomogeneous_T_188 ;  
   wire [31:0] _pmpHomogeneous_T_190 ;  
   wire [65:0] _GEN_166 ;  
   wire [65:0] _pmpHomogeneous_T_192 ;  
   wire _pmpHomogeneous_T_194 ;  
   wire _pmpHomogeneous_T_201 ;  
   wire _pmpHomogeneous_T_208 ;  
   wire _pmpHomogeneous_T_210 ;  
   wire _pmpHomogeneous_T_212 ;  
   wire _pmpHomogeneous_T_214 ;  
   wire _pmpHomogeneous_T_215 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_29 ;  
   wire pmpHomogeneous_beginsAfterUpper_5 ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_35 ;  
   wire [65:0] _GEN_174 ;  
   wire pmpHomogeneous_endsBeforeUpper_5 ;  
   wire _pmpHomogeneous_T_218 ;  
   wire _pmpHomogeneous_T_219 ;  
   wire _pmpHomogeneous_T_220 ;  
   wire _pmpHomogeneous_T_221 ;  
   wire _pmpHomogeneous_T_222 ;  
   wire _pmpHomogeneous_T_223 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_52 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_54 ;  
   wire pmpHomogeneous_maskHomogeneous_6 ;  
   wire [31:0] _pmpHomogeneous_T_225 ;  
   wire [31:0] _pmpHomogeneous_T_227 ;  
   wire [65:0] _GEN_175 ;  
   wire [65:0] _pmpHomogeneous_T_229 ;  
   wire _pmpHomogeneous_T_231 ;  
   wire _pmpHomogeneous_T_238 ;  
   wire _pmpHomogeneous_T_245 ;  
   wire _pmpHomogeneous_T_247 ;  
   wire _pmpHomogeneous_T_249 ;  
   wire _pmpHomogeneous_T_251 ;  
   wire _pmpHomogeneous_T_252 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_34 ;  
   wire pmpHomogeneous_beginsAfterUpper_6 ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_41 ;  
   wire [65:0] _GEN_183 ;  
   wire pmpHomogeneous_endsBeforeUpper_6 ;  
   wire _pmpHomogeneous_T_255 ;  
   wire _pmpHomogeneous_T_256 ;  
   wire _pmpHomogeneous_T_257 ;  
   wire _pmpHomogeneous_T_258 ;  
   wire _pmpHomogeneous_T_259 ;  
   wire _pmpHomogeneous_T_260 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_60 ;  
   wire _pmpHomogeneous_maskHomogeneous_T_62 ;  
   wire pmpHomogeneous_maskHomogeneous_7 ;  
   wire [31:0] _pmpHomogeneous_T_262 ;  
   wire [31:0] _pmpHomogeneous_T_264 ;  
   wire [65:0] _GEN_184 ;  
   wire [65:0] _pmpHomogeneous_T_266 ;  
   wire _pmpHomogeneous_T_268 ;  
   wire _pmpHomogeneous_T_275 ;  
   wire _pmpHomogeneous_T_282 ;  
   wire _pmpHomogeneous_T_284 ;  
   wire _pmpHomogeneous_T_286 ;  
   wire _pmpHomogeneous_T_288 ;  
   wire _pmpHomogeneous_T_289 ;  
   wire _pmpHomogeneous_beginsAfterUpper_T_39 ;  
   wire pmpHomogeneous_beginsAfterUpper_7 ;  
   wire [31:0] _pmpHomogeneous_endsBeforeUpper_T_47 ;  
   wire [65:0] _GEN_192 ;  
   wire pmpHomogeneous_endsBeforeUpper_7 ;  
   wire _pmpHomogeneous_T_292 ;  
   wire _pmpHomogeneous_T_293 ;  
   wire _pmpHomogeneous_T_294 ;  
   wire _pmpHomogeneous_T_295 ;  
   wire _pmpHomogeneous_T_296 ;  
   wire pmpHomogeneous ;  
   wire homogeneous ;  
   wire _T_100 ;  
   wire [2:0] _next_state_T ;  
   wire [2:0] _GEN_40 ;  
   wire _count_T_1 ;  
   wire _T_102 ;  
   wire [1:0] _count_T_3 ;  
   wire [2:0] _next_state_T_1 ;  
   wire [2:0] _GEN_43 ;  
   wire _T_103 ;  
   wire _T_104 ;  
   wire [2:0] _GEN_47 ;  
   wire _GEN_48 ;  
   wire _GEN_49 ;  
   wire _T_107 ;  
   wire [2:0] _GEN_54 ;  
   wire _GEN_55 ;  
   wire _GEN_56 ;  
   wire [2:0] _GEN_60 ;  
   wire _GEN_61 ;  
   wire _GEN_62 ;  
   wire _GEN_63 ;  
   wire _GEN_64 ;  
   wire [2:0] _GEN_67 ;  
   wire _GEN_68 ;  
   wire _GEN_70 ;  
   wire _GEN_71 ;  
   wire _GEN_75 ;  
   wire [2:0] _GEN_76 ;  
   wire _GEN_77 ;  
   wire _GEN_79 ;  
   wire _GEN_80 ;  
   wire [2:0] _GEN_82 ;  
   wire _GEN_87 ;  
   wire _GEN_88 ;  
   wire _r_pte_T_2 ;  
   wire _r_pte_T_4 ;  
   wire _r_pte_T_6 ;  
   wire [53:0] pte_2_ppn ;  
   wire [53:0] _r_pte_T_8_ppn ;  
   wire [53:0] pte_1_ppn ;  
   wire [53:0] _r_pte_T_9_ppn ;  
   wire _r_pte_T_9_d ;  
   wire _r_pte_T_9_a ;  
   wire _r_pte_T_9_g ;  
   wire _r_pte_T_9_u ;  
   wire _r_pte_T_9_x ;  
   wire _r_pte_T_9_w ;  
   wire _r_pte_T_9_r ;  
   wire _r_pte_T_9_v ;  
   wire [53:0] _r_pte_T_10_ppn ;  
   wire _r_pte_T_10_d ;  
   wire _r_pte_T_10_a ;  
   wire _r_pte_T_10_g ;  
   wire _r_pte_T_10_u ;  
   wire _r_pte_T_10_x ;  
   wire _r_pte_T_10_w ;  
   wire _r_pte_T_10_r ;  
   wire _r_pte_T_10_v ;  
   wire _GEN_90 ;  
   wire _GEN_91 ;  
   wire _T_121 ;  
   wire _T_123 ;  
   wire _l2_refill_T_1 ;  
   wire _l2_refill_T_3 ;  
   wire ae ;  
   wire [2:0] _GEN_102 ;  
   wire _GEN_104 ;  
   wire [2:0] _GEN_108 ;  
   wire _T_131 ;  
   wire _T_133 ;  
   reg [19:0] PTW_state ;  
   reg [31:0] _RAND_39 ;  
   reg PTW_cov[0:1048575] ;  
   reg [31:0] _RAND_40 ;  
   wire PTW_cov_read_data ;  
   wire [19:0] PTW_cov_read_addr ;  
   wire PTW_cov_write_data ;  
   wire [19:0] PTW_cov_write_addr ;  
   wire PTW_cov_write_mask ;  
   wire PTW_cov_write_en ;  
   reg [29:0] PTW_covSum ;  
   reg [31:0] _RAND_41 ;  
   wire [10:0] valid_shl ;  
   wire [19:0] valid_pad ;  
   wire [17:0] count_shl ;  
   wire [19:0] count_pad ;  
   wire [8:0] state_reg_shl ;  
   wire [19:0] state_reg_pad ;  
   wire [6:0] mem_resp_valid_shl ;  
   wire [19:0] mem_resp_valid_pad ;  
   wire [9:0] state_shl ;  
   wire [19:0] state_pad ;  
   wire [13:0] invalidated_shl ;  
   wire [19:0] invalidated_pad ;  
   wire [19:0] PTW_xor4 ;  
   wire [19:0] PTW_xor1 ;  
   wire [19:0] PTW_xor6 ;  
   wire [19:0] PTW_xor2 ;  
   wire [19:0] PTW_xor0 ;  
   wire [29:0] arb_sum ;  
   wire [29:0] state_barrier_sum ;  
   wire [29:0] r_pte_barrier_sum ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire stopEn2 ;  
   wire arb_metaAssert_wire ;  
   wire state_barrier_metaAssert_wire ;  
   wire r_pte_barrier_metaAssert_wire ;  
   wire PTW_or4 ;  
   wire PTW_or1 ;  
   wire PTW_or6 ;  
   wire PTW_or2 ;  
   wire PTW_or0 ;  
   reg PTW_metaAssert ;  
   reg [31:0] _RAND_42 ;  
  Arbiter arb(.io_in_0_ready(arb_io_in_0_ready),.io_in_0_valid(arb_io_in_0_valid),.io_in_0_bits_bits_addr(arb_io_in_0_bits_bits_addr),.io_in_1_ready(arb_io_in_1_ready),.io_in_1_valid(arb_io_in_1_valid),.io_in_1_bits_valid(arb_io_in_1_bits_valid),.io_in_1_bits_bits_addr(arb_io_in_1_bits_bits_addr),.io_out_ready(arb_io_out_ready),.io_out_valid(arb_io_out_valid),.io_out_bits_valid(arb_io_out_bits_valid),.io_out_bits_bits_addr(arb_io_out_bits_bits_addr),.io_chosen(arb_io_chosen),.io_covSum(arb_io_covSum),.metaAssert(arb_metaAssert)); 
  OptimizationBarrier_42 state_barrier(.io_x(state_barrier_io_x),.io_y(state_barrier_io_y),.io_covSum(state_barrier_io_covSum),.metaAssert(state_barrier_metaAssert)); 
  OptimizationBarrier_43 r_pte_barrier(.io_x_ppn(r_pte_barrier_io_x_ppn),.io_x_d(r_pte_barrier_io_x_d),.io_x_a(r_pte_barrier_io_x_a),.io_x_g(r_pte_barrier_io_x_g),.io_x_u(r_pte_barrier_io_x_u),.io_x_x(r_pte_barrier_io_x_x),.io_x_w(r_pte_barrier_io_x_w),.io_x_r(r_pte_barrier_io_x_r),.io_x_v(r_pte_barrier_io_x_v),.io_y_ppn(r_pte_barrier_io_y_ppn),.io_y_d(r_pte_barrier_io_y_d),.io_y_a(r_pte_barrier_io_y_a),.io_y_g(r_pte_barrier_io_y_g),.io_y_u(r_pte_barrier_io_y_u),.io_y_x(r_pte_barrier_io_y_x),.io_y_w(r_pte_barrier_io_y_w),.io_y_r(r_pte_barrier_io_y_r),.io_y_v(r_pte_barrier_io_y_v),.io_covSum(r_pte_barrier_io_covSum),.metaAssert(r_pte_barrier_metaAssert)); 
  assign _arb_io_out_ready_T=state==3'h0; 
  assign _clock_en_T=state!=3'h0; 
  assign tmp_v=mem_resp_data[0]; 
  assign tmp_r=mem_resp_data[1]; 
  assign tmp_w=mem_resp_data[2]; 
  assign tmp_x=mem_resp_data[3]; 
  assign tmp_u=mem_resp_data[4]; 
  assign tmp_g=mem_resp_data[5]; 
  assign tmp_a=mem_resp_data[6]; 
  assign tmp_d=mem_resp_data[7]; 
  assign tmp_ppn=mem_resp_data[63:10]; 
  assign _T_11=tmp_r|tmp_w; 
  assign _T_12=_T_11|tmp_x; 
  assign _T_13=count<=2'h0; 
  assign _T_15=tmp_ppn[17:9]!=9'h0; 
  assign _T_16=_T_13&_T_15; 
  assign _GEN_0=_T_16 ? 1'h0:tmp_v; 
  assign _T_17=count<=2'h1; 
  assign _T_19=tmp_ppn[8:0]!=9'h0; 
  assign _T_20=_T_17&_T_19; 
  assign _GEN_1=_T_20 ? 1'h0:_GEN_0; 
  assign res_v=_T_12 ? _GEN_1:tmp_v; 
  assign invalid_paddr=tmp_ppn[53:20]!=34'h0; 
  assign _traverse_T_1=res_v&~tmp_r; 
  assign _traverse_T_3=_traverse_T_1&~tmp_w; 
  assign _traverse_T_5=_traverse_T_3&~tmp_x; 
  assign _traverse_T_7=_traverse_T_5&~invalid_paddr; 
  assign _traverse_T_8=count<2'h2; 
  assign traverse=_traverse_T_7&_traverse_T_8; 
  assign vpn_idxs_0=r_req_addr[26:18]; 
  assign vpn_idxs_1=r_req_addr[17:9]; 
  assign vpn_idxs_2=r_req_addr[8:0]; 
  assign _pte_addr_vpn_idx_T=count==2'h1; 
  assign _pte_addr_vpn_idx_T_1=_pte_addr_vpn_idx_T ? vpn_idxs_1:vpn_idxs_0; 
  assign _pte_addr_vpn_idx_T_2=count==2'h2; 
  assign _pte_addr_vpn_idx_T_3=_pte_addr_vpn_idx_T_2 ? vpn_idxs_2:_pte_addr_vpn_idx_T_1; 
  assign _pte_addr_vpn_idx_T_4=count==2'h3; 
  assign vpn_idx=_pte_addr_vpn_idx_T_4 ? vpn_idxs_2:_pte_addr_vpn_idx_T_3; 
  assign _pte_addr_T={r_pte_ppn,vpn_idx}; 
  assign pte_addr={_pte_addr_T,3'h0}; 
  assign fragmented_superpage_ppn_choices_hi=r_pte_ppn[53:18]; 
  assign fragmented_superpage_ppn_choices_lo=r_req_addr[17:0]; 
  assign choices_0={fragmented_superpage_ppn_choices_hi,fragmented_superpage_ppn_choices_lo}; 
  assign fragmented_superpage_ppn_choices_hi_1=r_pte_ppn[53:9]; 
  assign choices_1={fragmented_superpage_ppn_choices_hi_1,vpn_idxs_2}; 
  assign fragmented_superpage_ppn_truncIdx=count[0]; 
  assign fragmented_superpage_ppn=fragmented_superpage_ppn_truncIdx ? choices_1:choices_0; 
  assign _T_22=arb_io_out_ready&arb_io_out_valid; 
  assign _GEN_115={34'b0,tags_0}; 
  assign lo_lo_lo=_GEN_115==pte_addr; 
  assign _GEN_116={34'b0,tags_1}; 
  assign lo_lo_hi=_GEN_116==pte_addr; 
  assign _GEN_117={34'b0,tags_2}; 
  assign lo_hi_lo=_GEN_117==pte_addr; 
  assign _GEN_118={34'b0,tags_3}; 
  assign lo_hi_hi=_GEN_118==pte_addr; 
  assign _GEN_119={34'b0,tags_4}; 
  assign hi_lo_lo=_GEN_119==pte_addr; 
  assign _GEN_120={34'b0,tags_5}; 
  assign hi_lo_hi=_GEN_120==pte_addr; 
  assign _GEN_121={34'b0,tags_6}; 
  assign hi_hi_lo=_GEN_121==pte_addr; 
  assign _GEN_122={34'b0,tags_7}; 
  assign hi_hi_hi=_GEN_122==pte_addr; 
  assign _T_23={hi_hi_hi,hi_hi_lo,hi_lo_hi,hi_lo_lo,lo_hi_hi,lo_hi_lo,lo_lo_hi,lo_lo_lo}; 
  assign hits=_T_23&valid; 
  assign hit=|hits; 
  assign _T_24=mem_resp_valid&traverse; 
  assign _T_26=_T_24&~hit; 
  assign _T_28=_T_26&~invalidated; 
  assign _T_29=&valid; 
  assign hi_1=state_reg[6]; 
  assign left_subtree_state=state_reg[5:3]; 
  assign right_subtree_state=state_reg[2:0]; 
  assign hi_2=left_subtree_state[2]; 
  assign left_subtree_state_1=left_subtree_state[1]; 
  assign right_subtree_state_1=left_subtree_state[0]; 
  assign lo_1=hi_2 ? left_subtree_state_1:right_subtree_state_1; 
  assign _T_32={hi_2,lo_1}; 
  assign hi_3=right_subtree_state[2]; 
  assign left_subtree_state_2=right_subtree_state[1]; 
  assign right_subtree_state_2=right_subtree_state[0]; 
  assign lo_2=hi_3 ? left_subtree_state_2:right_subtree_state_2; 
  assign _T_35={hi_3,lo_2}; 
  assign lo_3=hi_1 ? _T_32:_T_35; 
  assign _T_36={hi_1,lo_3}; 
  assign _T_38=~valid[0]; 
  assign _T_39=~valid[1]; 
  assign _T_40=~valid[2]; 
  assign _T_41=~valid[3]; 
  assign _T_42=~valid[4]; 
  assign _T_43=~valid[5]; 
  assign _T_44=~valid[6]; 
  assign _T_46=_T_44 ? 3'h6:3'h7; 
  assign _T_47=_T_43 ? 3'h5:_T_46; 
  assign _T_48=_T_42 ? 3'h4:_T_47; 
  assign _T_49=_T_41 ? 3'h3:_T_48; 
  assign _T_50=_T_40 ? 3'h2:_T_49; 
  assign _T_51=_T_39 ? 3'h1:_T_50; 
  assign _T_52=_T_38 ? 3'h0:_T_51; 
  assign r=_T_29 ? _T_36:_T_52; 
  assign _T_53=8'h1<<r; 
  assign _T_54=valid|_T_53; 
  assign res_ppn={34'b0,tmp_ppn[19:0]}; 
  assign _T_55=state==3'h1; 
  assign _T_56=hit&_T_55; 
  assign hi_4=hits[7:4]; 
  assign lo_4=hits[3:0]; 
  assign hi_5=|hi_4; 
  assign _T_57=hi_4|lo_4; 
  assign hi_6=_T_57[3:2]; 
  assign lo_5=_T_57[1:0]; 
  assign hi_7=|hi_6; 
  assign _T_58=hi_6|lo_5; 
  assign lo_6=_T_58[1]; 
  assign state_reg_touch_way_sized={hi_5,hi_7,lo_6}; 
  assign state_reg_hi_hi=~state_reg_touch_way_sized[2]; 
  assign state_reg_hi_hi_1=~state_reg_touch_way_sized[1]; 
  assign state_reg_hi_lo=state_reg_hi_hi_1 ? left_subtree_state_1:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo=state_reg_hi_hi_1 ? ~state_reg_touch_way_sized[0]:right_subtree_state_1; 
  assign _state_reg_T_7={state_reg_hi_hi_1,state_reg_hi_lo,state_reg_lo}; 
  assign state_reg_hi_lo_1=state_reg_hi_hi ? left_subtree_state:_state_reg_T_7; 
  assign state_reg_hi_lo_2=state_reg_hi_hi_1 ? left_subtree_state_2:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo_1=state_reg_hi_hi_1 ? ~state_reg_touch_way_sized[0]:right_subtree_state_2; 
  assign _state_reg_T_15={state_reg_hi_hi_1,state_reg_hi_lo_2,state_reg_lo_1}; 
  assign state_reg_lo_2=state_reg_hi_hi ? _state_reg_T_15:right_subtree_state; 
  assign _state_reg_T_16={state_reg_hi_hi,state_reg_hi_lo_1,state_reg_lo_2}; 
  assign _T_61=io_dpath_sfence_valid&~io_dpath_sfence_bits_rs1; 
  assign pte_cache_hit=hit&_traverse_T_8; 
  assign _T_79=hits[0] ? data_0:20'h0; 
  assign _T_80=hits[1] ? data_1:20'h0; 
  assign _T_81=hits[2] ? data_2:20'h0; 
  assign _T_82=hits[3] ? data_3:20'h0; 
  assign _T_83=hits[4] ? data_4:20'h0; 
  assign _T_84=hits[5] ? data_5:20'h0; 
  assign _T_85=hits[6] ? data_6:20'h0; 
  assign _T_86=hits[7] ? data_7:20'h0; 
  assign _T_87=_T_79|_T_80; 
  assign _T_88=_T_87|_T_81; 
  assign _T_89=_T_88|_T_82; 
  assign _T_90=_T_89|_T_83; 
  assign _T_91=_T_90|_T_84; 
  assign _T_92=_T_91|_T_85; 
  assign pte_cache_data=_T_92|_T_86; 
  assign _io_dpath_perf_pte_hit_T_1=pte_hit&_T_55; 
  assign _T_94=io_dpath_perf_pte_miss|io_dpath_perf_pte_hit; 
  assign _T_95=io_dpath_perf_l2hit&_T_94; 
  assign _T_98=~_T_95|reset; 
  assign _invalidated_T_1=invalidated&_clock_en_T; 
  assign _io_mem_req_valid_T_1=state==3'h3; 
  assign _pmaPgLevelHomogeneous_T_6=pte_addr^66'hc000000; 
  assign _pmaPgLevelHomogeneous_T_7={1'b0,$signed(_pmaPgLevelHomogeneous_T_6)}; 
  assign _pmaPgLevelHomogeneous_T_9=$signed(_pmaPgLevelHomogeneous_T_7)&-67'sh4000000; 
  assign _pmaPgLevelHomogeneous_T_10=$signed(_pmaPgLevelHomogeneous_T_9)==67'sh0; 
  assign _pmaPgLevelHomogeneous_T_11=pte_addr^66'h60000000; 
  assign _pmaPgLevelHomogeneous_T_12={1'b0,$signed(_pmaPgLevelHomogeneous_T_11)}; 
  assign _pmaPgLevelHomogeneous_T_14=$signed(_pmaPgLevelHomogeneous_T_12)&-67'sh20000000; 
  assign _pmaPgLevelHomogeneous_T_15=$signed(_pmaPgLevelHomogeneous_T_14)==67'sh0; 
  assign _pmaPgLevelHomogeneous_T_16=pte_addr^66'h80000000; 
  assign _pmaPgLevelHomogeneous_T_17={1'b0,$signed(_pmaPgLevelHomogeneous_T_16)}; 
  assign _pmaPgLevelHomogeneous_T_19=$signed(_pmaPgLevelHomogeneous_T_17)&-67'sh10000000; 
  assign _pmaPgLevelHomogeneous_T_20=$signed(_pmaPgLevelHomogeneous_T_19)==67'sh0; 
  assign _pmaPgLevelHomogeneous_T_22=_pmaPgLevelHomogeneous_T_10|_pmaPgLevelHomogeneous_T_15; 
  assign pmaPgLevelHomogeneous_1=_pmaPgLevelHomogeneous_T_22|_pmaPgLevelHomogeneous_T_20; 
  assign _pmaPgLevelHomogeneous_T_26={1'b0,$signed(pte_addr)}; 
  assign _pmaPgLevelHomogeneous_T_53=$signed(_pmaPgLevelHomogeneous_T_26)&-67'sh1000; 
  assign _pmaPgLevelHomogeneous_T_54=$signed(_pmaPgLevelHomogeneous_T_53)==67'sh0; 
  assign _pmaPgLevelHomogeneous_T_55=pte_addr^66'h3000; 
  assign _pmaPgLevelHomogeneous_T_56={1'b0,$signed(_pmaPgLevelHomogeneous_T_55)}; 
  assign _pmaPgLevelHomogeneous_T_58=$signed(_pmaPgLevelHomogeneous_T_56)&-67'sh1000; 
  assign _pmaPgLevelHomogeneous_T_59=$signed(_pmaPgLevelHomogeneous_T_58)==67'sh0; 
  assign _pmaPgLevelHomogeneous_T_60=pte_addr^66'h10000; 
  assign _pmaPgLevelHomogeneous_T_61={1'b0,$signed(_pmaPgLevelHomogeneous_T_60)}; 
  assign _pmaPgLevelHomogeneous_T_63=$signed(_pmaPgLevelHomogeneous_T_61)&-67'sh10000; 
  assign _pmaPgLevelHomogeneous_T_64=$signed(_pmaPgLevelHomogeneous_T_63)==67'sh0; 
  assign _pmaPgLevelHomogeneous_T_65=pte_addr^66'h2000000; 
  assign _pmaPgLevelHomogeneous_T_66={1'b0,$signed(_pmaPgLevelHomogeneous_T_65)}; 
  assign _pmaPgLevelHomogeneous_T_68=$signed(_pmaPgLevelHomogeneous_T_66)&-67'sh10000; 
  assign _pmaPgLevelHomogeneous_T_69=$signed(_pmaPgLevelHomogeneous_T_68)==67'sh0; 
  assign _pmaPgLevelHomogeneous_T_86=_pmaPgLevelHomogeneous_T_54|_pmaPgLevelHomogeneous_T_59; 
  assign _pmaPgLevelHomogeneous_T_87=_pmaPgLevelHomogeneous_T_86|_pmaPgLevelHomogeneous_T_64; 
  assign _pmaPgLevelHomogeneous_T_88=_pmaPgLevelHomogeneous_T_87|_pmaPgLevelHomogeneous_T_69; 
  assign _pmaPgLevelHomogeneous_T_89=_pmaPgLevelHomogeneous_T_88|_pmaPgLevelHomogeneous_T_10; 
  assign _pmaPgLevelHomogeneous_T_90=_pmaPgLevelHomogeneous_T_89|_pmaPgLevelHomogeneous_T_15; 
  assign pmaPgLevelHomogeneous_2=_pmaPgLevelHomogeneous_T_90|_pmaPgLevelHomogeneous_T_20; 
  assign _pmaHomogeneous_T_1=_pte_addr_vpn_idx_T&pmaPgLevelHomogeneous_1; 
  assign _pmaHomogeneous_T_3=_pte_addr_vpn_idx_T_2 ? pmaPgLevelHomogeneous_2:_pmaHomogeneous_T_1; 
  assign pmaHomogeneous=_pte_addr_vpn_idx_T_4 ? pmaPgLevelHomogeneous_2:_pmaHomogeneous_T_3; 
  assign _pmpHomogeneous_T_1={pte_addr[65:12],12'h0}; 
  assign _pmpHomogeneous_maskHomogeneous_T_4=_pte_addr_vpn_idx_T ? io_dpath_pmp_0_mask[20]:io_dpath_pmp_0_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_6=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_0_mask[11]:_pmpHomogeneous_maskHomogeneous_T_4; 
  assign pmpHomogeneous_maskHomogeneous=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_0_mask[11]:_pmpHomogeneous_maskHomogeneous_T_6; 
  assign _pmpHomogeneous_T_3={io_dpath_pmp_0_addr,2'h0}; 
  assign _pmpHomogeneous_T_5=~_pmpHomogeneous_T_3|32'h3; 
  assign _GEN_123={34'b0,~_pmpHomogeneous_T_5}; 
  assign _pmpHomogeneous_T_7=_pmpHomogeneous_T_1^_GEN_123; 
  assign _pmpHomogeneous_T_9=_pmpHomogeneous_T_7[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_16=_pmpHomogeneous_T_7[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_23=_pmpHomogeneous_T_7[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_25=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_16:_pmpHomogeneous_T_9; 
  assign _pmpHomogeneous_T_27=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_23:_pmpHomogeneous_T_25; 
  assign _pmpHomogeneous_T_29=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_23:_pmpHomogeneous_T_27; 
  assign _pmpHomogeneous_T_30=pmpHomogeneous_maskHomogeneous|_pmpHomogeneous_T_29; 
  assign _pmpHomogeneous_beginsAfterUpper_T_4=_pmpHomogeneous_T_1<_GEN_123; 
  assign pmpHomogeneous_beginsAfterUpper=~_pmpHomogeneous_beginsAfterUpper_T_4; 
  assign _pmpHomogeneous_pgMask_T_1=_pte_addr_vpn_idx_T ? 32'hffe00000:32'hc0000000; 
  assign _pmpHomogeneous_pgMask_T_3=_pte_addr_vpn_idx_T_2 ? 32'hfffff000:_pmpHomogeneous_pgMask_T_1; 
  assign pmpHomogeneous_pgMask=_pte_addr_vpn_idx_T_4 ? 32'hfffff000:_pmpHomogeneous_pgMask_T_3; 
  assign _GEN_127={34'b0,pmpHomogeneous_pgMask}; 
  assign _pmpHomogeneous_endsBeforeLower_T=_pmpHomogeneous_T_1&_GEN_127; 
  assign _pmpHomogeneous_endsBeforeUpper_T_5=~_pmpHomogeneous_T_5&pmpHomogeneous_pgMask; 
  assign _GEN_129={34'b0,_pmpHomogeneous_endsBeforeUpper_T_5}; 
  assign pmpHomogeneous_endsBeforeUpper=_pmpHomogeneous_endsBeforeLower_T<_GEN_129; 
  assign _pmpHomogeneous_T_35=pmpHomogeneous_beginsAfterUpper|pmpHomogeneous_endsBeforeUpper; 
  assign _pmpHomogeneous_T_36=~io_dpath_pmp_0_cfg_a[0]|_pmpHomogeneous_T_35; 
  assign _pmpHomogeneous_T_37=io_dpath_pmp_0_cfg_a[1] ? _pmpHomogeneous_T_30:_pmpHomogeneous_T_36; 
  assign _pmpHomogeneous_maskHomogeneous_T_12=_pte_addr_vpn_idx_T ? io_dpath_pmp_1_mask[20]:io_dpath_pmp_1_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_14=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_1_mask[11]:_pmpHomogeneous_maskHomogeneous_T_12; 
  assign pmpHomogeneous_maskHomogeneous_1=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_1_mask[11]:_pmpHomogeneous_maskHomogeneous_T_14; 
  assign _pmpHomogeneous_T_40={io_dpath_pmp_1_addr,2'h0}; 
  assign _pmpHomogeneous_T_42=~_pmpHomogeneous_T_40|32'h3; 
  assign _GEN_130={34'b0,~_pmpHomogeneous_T_42}; 
  assign _pmpHomogeneous_T_44=_pmpHomogeneous_T_1^_GEN_130; 
  assign _pmpHomogeneous_T_46=_pmpHomogeneous_T_44[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_53=_pmpHomogeneous_T_44[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_60=_pmpHomogeneous_T_44[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_62=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_53:_pmpHomogeneous_T_46; 
  assign _pmpHomogeneous_T_64=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_60:_pmpHomogeneous_T_62; 
  assign _pmpHomogeneous_T_66=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_60:_pmpHomogeneous_T_64; 
  assign _pmpHomogeneous_T_67=pmpHomogeneous_maskHomogeneous_1|_pmpHomogeneous_T_66; 
  assign _pmpHomogeneous_beginsAfterUpper_T_9=_pmpHomogeneous_T_1<_GEN_130; 
  assign pmpHomogeneous_beginsAfterUpper_1=~_pmpHomogeneous_beginsAfterUpper_T_9; 
  assign _pmpHomogeneous_endsBeforeUpper_T_11=~_pmpHomogeneous_T_42&pmpHomogeneous_pgMask; 
  assign _GEN_138={34'b0,_pmpHomogeneous_endsBeforeUpper_T_11}; 
  assign pmpHomogeneous_endsBeforeUpper_1=_pmpHomogeneous_endsBeforeLower_T<_GEN_138; 
  assign _pmpHomogeneous_T_70=pmpHomogeneous_endsBeforeUpper|pmpHomogeneous_beginsAfterUpper_1; 
  assign _pmpHomogeneous_T_71=pmpHomogeneous_beginsAfterUpper&pmpHomogeneous_endsBeforeUpper_1; 
  assign _pmpHomogeneous_T_72=_pmpHomogeneous_T_70|_pmpHomogeneous_T_71; 
  assign _pmpHomogeneous_T_73=~io_dpath_pmp_1_cfg_a[0]|_pmpHomogeneous_T_72; 
  assign _pmpHomogeneous_T_74=io_dpath_pmp_1_cfg_a[1] ? _pmpHomogeneous_T_67:_pmpHomogeneous_T_73; 
  assign _pmpHomogeneous_T_75=_pmpHomogeneous_T_37&_pmpHomogeneous_T_74; 
  assign _pmpHomogeneous_maskHomogeneous_T_20=_pte_addr_vpn_idx_T ? io_dpath_pmp_2_mask[20]:io_dpath_pmp_2_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_22=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_2_mask[11]:_pmpHomogeneous_maskHomogeneous_T_20; 
  assign pmpHomogeneous_maskHomogeneous_2=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_2_mask[11]:_pmpHomogeneous_maskHomogeneous_T_22; 
  assign _pmpHomogeneous_T_77={io_dpath_pmp_2_addr,2'h0}; 
  assign _pmpHomogeneous_T_79=~_pmpHomogeneous_T_77|32'h3; 
  assign _GEN_139={34'b0,~_pmpHomogeneous_T_79}; 
  assign _pmpHomogeneous_T_81=_pmpHomogeneous_T_1^_GEN_139; 
  assign _pmpHomogeneous_T_83=_pmpHomogeneous_T_81[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_90=_pmpHomogeneous_T_81[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_97=_pmpHomogeneous_T_81[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_99=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_90:_pmpHomogeneous_T_83; 
  assign _pmpHomogeneous_T_101=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_97:_pmpHomogeneous_T_99; 
  assign _pmpHomogeneous_T_103=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_97:_pmpHomogeneous_T_101; 
  assign _pmpHomogeneous_T_104=pmpHomogeneous_maskHomogeneous_2|_pmpHomogeneous_T_103; 
  assign _pmpHomogeneous_beginsAfterUpper_T_14=_pmpHomogeneous_T_1<_GEN_139; 
  assign pmpHomogeneous_beginsAfterUpper_2=~_pmpHomogeneous_beginsAfterUpper_T_14; 
  assign _pmpHomogeneous_endsBeforeUpper_T_17=~_pmpHomogeneous_T_79&pmpHomogeneous_pgMask; 
  assign _GEN_147={34'b0,_pmpHomogeneous_endsBeforeUpper_T_17}; 
  assign pmpHomogeneous_endsBeforeUpper_2=_pmpHomogeneous_endsBeforeLower_T<_GEN_147; 
  assign _pmpHomogeneous_T_107=pmpHomogeneous_endsBeforeUpper_1|pmpHomogeneous_beginsAfterUpper_2; 
  assign _pmpHomogeneous_T_108=pmpHomogeneous_beginsAfterUpper_1&pmpHomogeneous_endsBeforeUpper_2; 
  assign _pmpHomogeneous_T_109=_pmpHomogeneous_T_107|_pmpHomogeneous_T_108; 
  assign _pmpHomogeneous_T_110=~io_dpath_pmp_2_cfg_a[0]|_pmpHomogeneous_T_109; 
  assign _pmpHomogeneous_T_111=io_dpath_pmp_2_cfg_a[1] ? _pmpHomogeneous_T_104:_pmpHomogeneous_T_110; 
  assign _pmpHomogeneous_T_112=_pmpHomogeneous_T_75&_pmpHomogeneous_T_111; 
  assign _pmpHomogeneous_maskHomogeneous_T_28=_pte_addr_vpn_idx_T ? io_dpath_pmp_3_mask[20]:io_dpath_pmp_3_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_30=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_3_mask[11]:_pmpHomogeneous_maskHomogeneous_T_28; 
  assign pmpHomogeneous_maskHomogeneous_3=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_3_mask[11]:_pmpHomogeneous_maskHomogeneous_T_30; 
  assign _pmpHomogeneous_T_114={io_dpath_pmp_3_addr,2'h0}; 
  assign _pmpHomogeneous_T_116=~_pmpHomogeneous_T_114|32'h3; 
  assign _GEN_148={34'b0,~_pmpHomogeneous_T_116}; 
  assign _pmpHomogeneous_T_118=_pmpHomogeneous_T_1^_GEN_148; 
  assign _pmpHomogeneous_T_120=_pmpHomogeneous_T_118[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_127=_pmpHomogeneous_T_118[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_134=_pmpHomogeneous_T_118[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_136=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_127:_pmpHomogeneous_T_120; 
  assign _pmpHomogeneous_T_138=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_134:_pmpHomogeneous_T_136; 
  assign _pmpHomogeneous_T_140=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_134:_pmpHomogeneous_T_138; 
  assign _pmpHomogeneous_T_141=pmpHomogeneous_maskHomogeneous_3|_pmpHomogeneous_T_140; 
  assign _pmpHomogeneous_beginsAfterUpper_T_19=_pmpHomogeneous_T_1<_GEN_148; 
  assign pmpHomogeneous_beginsAfterUpper_3=~_pmpHomogeneous_beginsAfterUpper_T_19; 
  assign _pmpHomogeneous_endsBeforeUpper_T_23=~_pmpHomogeneous_T_116&pmpHomogeneous_pgMask; 
  assign _GEN_156={34'b0,_pmpHomogeneous_endsBeforeUpper_T_23}; 
  assign pmpHomogeneous_endsBeforeUpper_3=_pmpHomogeneous_endsBeforeLower_T<_GEN_156; 
  assign _pmpHomogeneous_T_144=pmpHomogeneous_endsBeforeUpper_2|pmpHomogeneous_beginsAfterUpper_3; 
  assign _pmpHomogeneous_T_145=pmpHomogeneous_beginsAfterUpper_2&pmpHomogeneous_endsBeforeUpper_3; 
  assign _pmpHomogeneous_T_146=_pmpHomogeneous_T_144|_pmpHomogeneous_T_145; 
  assign _pmpHomogeneous_T_147=~io_dpath_pmp_3_cfg_a[0]|_pmpHomogeneous_T_146; 
  assign _pmpHomogeneous_T_148=io_dpath_pmp_3_cfg_a[1] ? _pmpHomogeneous_T_141:_pmpHomogeneous_T_147; 
  assign _pmpHomogeneous_T_149=_pmpHomogeneous_T_112&_pmpHomogeneous_T_148; 
  assign _pmpHomogeneous_maskHomogeneous_T_36=_pte_addr_vpn_idx_T ? io_dpath_pmp_4_mask[20]:io_dpath_pmp_4_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_38=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_4_mask[11]:_pmpHomogeneous_maskHomogeneous_T_36; 
  assign pmpHomogeneous_maskHomogeneous_4=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_4_mask[11]:_pmpHomogeneous_maskHomogeneous_T_38; 
  assign _pmpHomogeneous_T_151={io_dpath_pmp_4_addr,2'h0}; 
  assign _pmpHomogeneous_T_153=~_pmpHomogeneous_T_151|32'h3; 
  assign _GEN_157={34'b0,~_pmpHomogeneous_T_153}; 
  assign _pmpHomogeneous_T_155=_pmpHomogeneous_T_1^_GEN_157; 
  assign _pmpHomogeneous_T_157=_pmpHomogeneous_T_155[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_164=_pmpHomogeneous_T_155[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_171=_pmpHomogeneous_T_155[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_173=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_164:_pmpHomogeneous_T_157; 
  assign _pmpHomogeneous_T_175=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_171:_pmpHomogeneous_T_173; 
  assign _pmpHomogeneous_T_177=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_171:_pmpHomogeneous_T_175; 
  assign _pmpHomogeneous_T_178=pmpHomogeneous_maskHomogeneous_4|_pmpHomogeneous_T_177; 
  assign _pmpHomogeneous_beginsAfterUpper_T_24=_pmpHomogeneous_T_1<_GEN_157; 
  assign pmpHomogeneous_beginsAfterUpper_4=~_pmpHomogeneous_beginsAfterUpper_T_24; 
  assign _pmpHomogeneous_endsBeforeUpper_T_29=~_pmpHomogeneous_T_153&pmpHomogeneous_pgMask; 
  assign _GEN_165={34'b0,_pmpHomogeneous_endsBeforeUpper_T_29}; 
  assign pmpHomogeneous_endsBeforeUpper_4=_pmpHomogeneous_endsBeforeLower_T<_GEN_165; 
  assign _pmpHomogeneous_T_181=pmpHomogeneous_endsBeforeUpper_3|pmpHomogeneous_beginsAfterUpper_4; 
  assign _pmpHomogeneous_T_182=pmpHomogeneous_beginsAfterUpper_3&pmpHomogeneous_endsBeforeUpper_4; 
  assign _pmpHomogeneous_T_183=_pmpHomogeneous_T_181|_pmpHomogeneous_T_182; 
  assign _pmpHomogeneous_T_184=~io_dpath_pmp_4_cfg_a[0]|_pmpHomogeneous_T_183; 
  assign _pmpHomogeneous_T_185=io_dpath_pmp_4_cfg_a[1] ? _pmpHomogeneous_T_178:_pmpHomogeneous_T_184; 
  assign _pmpHomogeneous_T_186=_pmpHomogeneous_T_149&_pmpHomogeneous_T_185; 
  assign _pmpHomogeneous_maskHomogeneous_T_44=_pte_addr_vpn_idx_T ? io_dpath_pmp_5_mask[20]:io_dpath_pmp_5_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_46=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_5_mask[11]:_pmpHomogeneous_maskHomogeneous_T_44; 
  assign pmpHomogeneous_maskHomogeneous_5=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_5_mask[11]:_pmpHomogeneous_maskHomogeneous_T_46; 
  assign _pmpHomogeneous_T_188={io_dpath_pmp_5_addr,2'h0}; 
  assign _pmpHomogeneous_T_190=~_pmpHomogeneous_T_188|32'h3; 
  assign _GEN_166={34'b0,~_pmpHomogeneous_T_190}; 
  assign _pmpHomogeneous_T_192=_pmpHomogeneous_T_1^_GEN_166; 
  assign _pmpHomogeneous_T_194=_pmpHomogeneous_T_192[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_201=_pmpHomogeneous_T_192[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_208=_pmpHomogeneous_T_192[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_210=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_201:_pmpHomogeneous_T_194; 
  assign _pmpHomogeneous_T_212=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_208:_pmpHomogeneous_T_210; 
  assign _pmpHomogeneous_T_214=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_208:_pmpHomogeneous_T_212; 
  assign _pmpHomogeneous_T_215=pmpHomogeneous_maskHomogeneous_5|_pmpHomogeneous_T_214; 
  assign _pmpHomogeneous_beginsAfterUpper_T_29=_pmpHomogeneous_T_1<_GEN_166; 
  assign pmpHomogeneous_beginsAfterUpper_5=~_pmpHomogeneous_beginsAfterUpper_T_29; 
  assign _pmpHomogeneous_endsBeforeUpper_T_35=~_pmpHomogeneous_T_190&pmpHomogeneous_pgMask; 
  assign _GEN_174={34'b0,_pmpHomogeneous_endsBeforeUpper_T_35}; 
  assign pmpHomogeneous_endsBeforeUpper_5=_pmpHomogeneous_endsBeforeLower_T<_GEN_174; 
  assign _pmpHomogeneous_T_218=pmpHomogeneous_endsBeforeUpper_4|pmpHomogeneous_beginsAfterUpper_5; 
  assign _pmpHomogeneous_T_219=pmpHomogeneous_beginsAfterUpper_4&pmpHomogeneous_endsBeforeUpper_5; 
  assign _pmpHomogeneous_T_220=_pmpHomogeneous_T_218|_pmpHomogeneous_T_219; 
  assign _pmpHomogeneous_T_221=~io_dpath_pmp_5_cfg_a[0]|_pmpHomogeneous_T_220; 
  assign _pmpHomogeneous_T_222=io_dpath_pmp_5_cfg_a[1] ? _pmpHomogeneous_T_215:_pmpHomogeneous_T_221; 
  assign _pmpHomogeneous_T_223=_pmpHomogeneous_T_186&_pmpHomogeneous_T_222; 
  assign _pmpHomogeneous_maskHomogeneous_T_52=_pte_addr_vpn_idx_T ? io_dpath_pmp_6_mask[20]:io_dpath_pmp_6_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_54=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_6_mask[11]:_pmpHomogeneous_maskHomogeneous_T_52; 
  assign pmpHomogeneous_maskHomogeneous_6=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_6_mask[11]:_pmpHomogeneous_maskHomogeneous_T_54; 
  assign _pmpHomogeneous_T_225={io_dpath_pmp_6_addr,2'h0}; 
  assign _pmpHomogeneous_T_227=~_pmpHomogeneous_T_225|32'h3; 
  assign _GEN_175={34'b0,~_pmpHomogeneous_T_227}; 
  assign _pmpHomogeneous_T_229=_pmpHomogeneous_T_1^_GEN_175; 
  assign _pmpHomogeneous_T_231=_pmpHomogeneous_T_229[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_238=_pmpHomogeneous_T_229[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_245=_pmpHomogeneous_T_229[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_247=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_238:_pmpHomogeneous_T_231; 
  assign _pmpHomogeneous_T_249=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_245:_pmpHomogeneous_T_247; 
  assign _pmpHomogeneous_T_251=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_245:_pmpHomogeneous_T_249; 
  assign _pmpHomogeneous_T_252=pmpHomogeneous_maskHomogeneous_6|_pmpHomogeneous_T_251; 
  assign _pmpHomogeneous_beginsAfterUpper_T_34=_pmpHomogeneous_T_1<_GEN_175; 
  assign pmpHomogeneous_beginsAfterUpper_6=~_pmpHomogeneous_beginsAfterUpper_T_34; 
  assign _pmpHomogeneous_endsBeforeUpper_T_41=~_pmpHomogeneous_T_227&pmpHomogeneous_pgMask; 
  assign _GEN_183={34'b0,_pmpHomogeneous_endsBeforeUpper_T_41}; 
  assign pmpHomogeneous_endsBeforeUpper_6=_pmpHomogeneous_endsBeforeLower_T<_GEN_183; 
  assign _pmpHomogeneous_T_255=pmpHomogeneous_endsBeforeUpper_5|pmpHomogeneous_beginsAfterUpper_6; 
  assign _pmpHomogeneous_T_256=pmpHomogeneous_beginsAfterUpper_5&pmpHomogeneous_endsBeforeUpper_6; 
  assign _pmpHomogeneous_T_257=_pmpHomogeneous_T_255|_pmpHomogeneous_T_256; 
  assign _pmpHomogeneous_T_258=~io_dpath_pmp_6_cfg_a[0]|_pmpHomogeneous_T_257; 
  assign _pmpHomogeneous_T_259=io_dpath_pmp_6_cfg_a[1] ? _pmpHomogeneous_T_252:_pmpHomogeneous_T_258; 
  assign _pmpHomogeneous_T_260=_pmpHomogeneous_T_223&_pmpHomogeneous_T_259; 
  assign _pmpHomogeneous_maskHomogeneous_T_60=_pte_addr_vpn_idx_T ? io_dpath_pmp_7_mask[20]:io_dpath_pmp_7_mask[29]; 
  assign _pmpHomogeneous_maskHomogeneous_T_62=_pte_addr_vpn_idx_T_2 ? io_dpath_pmp_7_mask[11]:_pmpHomogeneous_maskHomogeneous_T_60; 
  assign pmpHomogeneous_maskHomogeneous_7=_pte_addr_vpn_idx_T_4 ? io_dpath_pmp_7_mask[11]:_pmpHomogeneous_maskHomogeneous_T_62; 
  assign _pmpHomogeneous_T_262={io_dpath_pmp_7_addr,2'h0}; 
  assign _pmpHomogeneous_T_264=~_pmpHomogeneous_T_262|32'h3; 
  assign _GEN_184={34'b0,~_pmpHomogeneous_T_264}; 
  assign _pmpHomogeneous_T_266=_pmpHomogeneous_T_1^_GEN_184; 
  assign _pmpHomogeneous_T_268=_pmpHomogeneous_T_266[65:30]!=36'h0; 
  assign _pmpHomogeneous_T_275=_pmpHomogeneous_T_266[65:21]!=45'h0; 
  assign _pmpHomogeneous_T_282=_pmpHomogeneous_T_266[65:12]!=54'h0; 
  assign _pmpHomogeneous_T_284=_pte_addr_vpn_idx_T ? _pmpHomogeneous_T_275:_pmpHomogeneous_T_268; 
  assign _pmpHomogeneous_T_286=_pte_addr_vpn_idx_T_2 ? _pmpHomogeneous_T_282:_pmpHomogeneous_T_284; 
  assign _pmpHomogeneous_T_288=_pte_addr_vpn_idx_T_4 ? _pmpHomogeneous_T_282:_pmpHomogeneous_T_286; 
  assign _pmpHomogeneous_T_289=pmpHomogeneous_maskHomogeneous_7|_pmpHomogeneous_T_288; 
  assign _pmpHomogeneous_beginsAfterUpper_T_39=_pmpHomogeneous_T_1<_GEN_184; 
  assign pmpHomogeneous_beginsAfterUpper_7=~_pmpHomogeneous_beginsAfterUpper_T_39; 
  assign _pmpHomogeneous_endsBeforeUpper_T_47=~_pmpHomogeneous_T_264&pmpHomogeneous_pgMask; 
  assign _GEN_192={34'b0,_pmpHomogeneous_endsBeforeUpper_T_47}; 
  assign pmpHomogeneous_endsBeforeUpper_7=_pmpHomogeneous_endsBeforeLower_T<_GEN_192; 
  assign _pmpHomogeneous_T_292=pmpHomogeneous_endsBeforeUpper_6|pmpHomogeneous_beginsAfterUpper_7; 
  assign _pmpHomogeneous_T_293=pmpHomogeneous_beginsAfterUpper_6&pmpHomogeneous_endsBeforeUpper_7; 
  assign _pmpHomogeneous_T_294=_pmpHomogeneous_T_292|_pmpHomogeneous_T_293; 
  assign _pmpHomogeneous_T_295=~io_dpath_pmp_7_cfg_a[0]|_pmpHomogeneous_T_294; 
  assign _pmpHomogeneous_T_296=io_dpath_pmp_7_cfg_a[1] ? _pmpHomogeneous_T_289:_pmpHomogeneous_T_295; 
  assign pmpHomogeneous=_pmpHomogeneous_T_260&_pmpHomogeneous_T_296; 
  assign homogeneous=pmaHomogeneous&pmpHomogeneous; 
  assign _T_100=3'h0==state; 
  assign _next_state_T=arb_io_out_bits_valid ? 3'h1:3'h0; 
  assign _GEN_40=_T_22 ? _next_state_T:state; 
  assign _count_T_1=1'h0-1'h0; 
  assign _T_102=3'h1==state; 
  assign _count_T_3=count+2'h1; 
  assign _next_state_T_1=io_mem_req_ready ? 3'h2:3'h1; 
  assign _GEN_43=pte_cache_hit ? state:_next_state_T_1; 
  assign _T_103=3'h2==state; 
  assign _T_104=3'h4==state; 
  assign _GEN_47=io_mem_s2_xcpt_ae_ld ? 3'h0:3'h5; 
  assign _GEN_48=io_mem_s2_xcpt_ae_ld&~r_req_dest; 
  assign _GEN_49=io_mem_s2_xcpt_ae_ld&r_req_dest; 
  assign _T_107=3'h7==state; 
  assign _GEN_54=_T_107 ? 3'h0:state; 
  assign _GEN_55=_T_107&~r_req_dest; 
  assign _GEN_56=_T_107&r_req_dest; 
  assign _GEN_60=_T_104 ? _GEN_47:_GEN_54; 
  assign _GEN_61=_T_104&_traverse_T_8; 
  assign _GEN_62=_T_104&io_mem_s2_xcpt_ae_ld; 
  assign _GEN_63=_T_104 ? _GEN_48:_GEN_55; 
  assign _GEN_64=_T_104 ? _GEN_49:_GEN_56; 
  assign _GEN_67=_T_103 ? 3'h4:_GEN_60; 
  assign _GEN_68=_T_103 ? 1'h0:_GEN_61; 
  assign _GEN_70=_T_103 ? 1'h0:_GEN_63; 
  assign _GEN_71=_T_103 ? 1'h0:_GEN_64; 
  assign _GEN_75=_T_102&pte_cache_hit; 
  assign _GEN_76=_T_102 ? _GEN_43:_GEN_67; 
  assign _GEN_77=_T_102 ? 1'h0:_GEN_68; 
  assign _GEN_79=_T_102 ? 1'h0:_GEN_70; 
  assign _GEN_80=_T_102 ? 1'h0:_GEN_71; 
  assign _GEN_82=_T_100 ? _GEN_40:_GEN_76; 
  assign _GEN_87=_T_100 ? 1'h0:_GEN_79; 
  assign _GEN_88=_T_100 ? 1'h0:_GEN_80; 
  assign _r_pte_T_2=state==3'h7; 
  assign _r_pte_T_4=_r_pte_T_2&~homogeneous; 
  assign _r_pte_T_6=_T_55&pte_cache_hit; 
  assign pte_2_ppn={10'b0,io_dpath_ptbr_ppn}; 
  assign _r_pte_T_8_ppn=_T_22 ? pte_2_ppn:r_pte_ppn; 
  assign pte_1_ppn={34'b0,pte_cache_data}; 
  assign _r_pte_T_9_ppn=_r_pte_T_6 ? pte_1_ppn:_r_pte_T_8_ppn; 
  assign _r_pte_T_9_d=_r_pte_T_6 ? 1'h0:r_pte_d; 
  assign _r_pte_T_9_a=_r_pte_T_6 ? 1'h0:r_pte_a; 
  assign _r_pte_T_9_g=_r_pte_T_6 ? 1'h0:r_pte_g; 
  assign _r_pte_T_9_u=_r_pte_T_6 ? 1'h0:r_pte_u; 
  assign _r_pte_T_9_x=_r_pte_T_6 ? 1'h0:r_pte_x; 
  assign _r_pte_T_9_w=_r_pte_T_6 ? 1'h0:r_pte_w; 
  assign _r_pte_T_9_r=_r_pte_T_6 ? 1'h0:r_pte_r; 
  assign _r_pte_T_9_v=_r_pte_T_6 ? 1'h0:r_pte_v; 
  assign _r_pte_T_10_ppn=_r_pte_T_4 ? fragmented_superpage_ppn:_r_pte_T_9_ppn; 
  assign _r_pte_T_10_d=_r_pte_T_4 ? r_pte_d:_r_pte_T_9_d; 
  assign _r_pte_T_10_a=_r_pte_T_4 ? r_pte_a:_r_pte_T_9_a; 
  assign _r_pte_T_10_g=_r_pte_T_4 ? r_pte_g:_r_pte_T_9_g; 
  assign _r_pte_T_10_u=_r_pte_T_4 ? r_pte_u:_r_pte_T_9_u; 
  assign _r_pte_T_10_x=_r_pte_T_4 ? r_pte_x:_r_pte_T_9_x; 
  assign _r_pte_T_10_w=_r_pte_T_4 ? r_pte_w:_r_pte_T_9_w; 
  assign _r_pte_T_10_r=_r_pte_T_4 ? r_pte_r:_r_pte_T_9_r; 
  assign _r_pte_T_10_v=_r_pte_T_4 ? r_pte_v:_r_pte_T_9_v; 
  assign _GEN_90=~r_req_dest|_GEN_87; 
  assign _GEN_91=r_req_dest|_GEN_88; 
  assign _T_121=state==3'h5; 
  assign _T_123=_T_121|reset; 
  assign _l2_refill_T_1=res_v&~invalid_paddr; 
  assign _l2_refill_T_3=_l2_refill_T_1&_pte_addr_vpn_idx_T_2; 
  assign ae=res_v&invalid_paddr; 
  assign _GEN_102=traverse ? 3'h1:3'h0; 
  assign _GEN_104=traverse ? 1'h0:_l2_refill_T_3; 
  assign _GEN_108=mem_resp_valid ? _GEN_102:_GEN_82; 
  assign _T_131=state==3'h4; 
  assign _T_133=_T_131|reset; 
  assign io_requestor_0_req_ready=arb_io_in_0_ready; 
  assign io_requestor_0_resp_valid=resp_valid_0; 
  assign io_requestor_0_resp_bits_ae=resp_ae; 
  assign io_requestor_0_resp_bits_pte_ppn=r_pte_ppn; 
  assign io_requestor_0_resp_bits_pte_d=r_pte_d; 
  assign io_requestor_0_resp_bits_pte_a=r_pte_a; 
  assign io_requestor_0_resp_bits_pte_g=r_pte_g; 
  assign io_requestor_0_resp_bits_pte_u=r_pte_u; 
  assign io_requestor_0_resp_bits_pte_x=r_pte_x; 
  assign io_requestor_0_resp_bits_pte_w=r_pte_w; 
  assign io_requestor_0_resp_bits_pte_r=r_pte_r; 
  assign io_requestor_0_resp_bits_pte_v=r_pte_v; 
  assign io_requestor_0_resp_bits_level=count; 
  assign io_requestor_0_resp_bits_homogeneous=pmaHomogeneous&pmpHomogeneous; 
  assign io_requestor_0_ptbr_mode=io_dpath_ptbr_mode; 
  assign io_requestor_0_status_debug=io_dpath_status_debug; 
  assign io_requestor_0_status_dprv=io_dpath_status_dprv; 
  assign io_requestor_0_status_mxr=io_dpath_status_mxr; 
  assign io_requestor_0_status_sum=io_dpath_status_sum; 
  assign io_requestor_0_pmp_0_cfg_l=io_dpath_pmp_0_cfg_l; 
  assign io_requestor_0_pmp_0_cfg_a=io_dpath_pmp_0_cfg_a; 
  assign io_requestor_0_pmp_0_cfg_x=io_dpath_pmp_0_cfg_x; 
  assign io_requestor_0_pmp_0_cfg_w=io_dpath_pmp_0_cfg_w; 
  assign io_requestor_0_pmp_0_cfg_r=io_dpath_pmp_0_cfg_r; 
  assign io_requestor_0_pmp_0_addr=io_dpath_pmp_0_addr; 
  assign io_requestor_0_pmp_0_mask=io_dpath_pmp_0_mask; 
  assign io_requestor_0_pmp_1_cfg_l=io_dpath_pmp_1_cfg_l; 
  assign io_requestor_0_pmp_1_cfg_a=io_dpath_pmp_1_cfg_a; 
  assign io_requestor_0_pmp_1_cfg_x=io_dpath_pmp_1_cfg_x; 
  assign io_requestor_0_pmp_1_cfg_w=io_dpath_pmp_1_cfg_w; 
  assign io_requestor_0_pmp_1_cfg_r=io_dpath_pmp_1_cfg_r; 
  assign io_requestor_0_pmp_1_addr=io_dpath_pmp_1_addr; 
  assign io_requestor_0_pmp_1_mask=io_dpath_pmp_1_mask; 
  assign io_requestor_0_pmp_2_cfg_l=io_dpath_pmp_2_cfg_l; 
  assign io_requestor_0_pmp_2_cfg_a=io_dpath_pmp_2_cfg_a; 
  assign io_requestor_0_pmp_2_cfg_x=io_dpath_pmp_2_cfg_x; 
  assign io_requestor_0_pmp_2_cfg_w=io_dpath_pmp_2_cfg_w; 
  assign io_requestor_0_pmp_2_cfg_r=io_dpath_pmp_2_cfg_r; 
  assign io_requestor_0_pmp_2_addr=io_dpath_pmp_2_addr; 
  assign io_requestor_0_pmp_2_mask=io_dpath_pmp_2_mask; 
  assign io_requestor_0_pmp_3_cfg_l=io_dpath_pmp_3_cfg_l; 
  assign io_requestor_0_pmp_3_cfg_a=io_dpath_pmp_3_cfg_a; 
  assign io_requestor_0_pmp_3_cfg_x=io_dpath_pmp_3_cfg_x; 
  assign io_requestor_0_pmp_3_cfg_w=io_dpath_pmp_3_cfg_w; 
  assign io_requestor_0_pmp_3_cfg_r=io_dpath_pmp_3_cfg_r; 
  assign io_requestor_0_pmp_3_addr=io_dpath_pmp_3_addr; 
  assign io_requestor_0_pmp_3_mask=io_dpath_pmp_3_mask; 
  assign io_requestor_0_pmp_4_cfg_l=io_dpath_pmp_4_cfg_l; 
  assign io_requestor_0_pmp_4_cfg_a=io_dpath_pmp_4_cfg_a; 
  assign io_requestor_0_pmp_4_cfg_x=io_dpath_pmp_4_cfg_x; 
  assign io_requestor_0_pmp_4_cfg_w=io_dpath_pmp_4_cfg_w; 
  assign io_requestor_0_pmp_4_cfg_r=io_dpath_pmp_4_cfg_r; 
  assign io_requestor_0_pmp_4_addr=io_dpath_pmp_4_addr; 
  assign io_requestor_0_pmp_4_mask=io_dpath_pmp_4_mask; 
  assign io_requestor_0_pmp_5_cfg_l=io_dpath_pmp_5_cfg_l; 
  assign io_requestor_0_pmp_5_cfg_a=io_dpath_pmp_5_cfg_a; 
  assign io_requestor_0_pmp_5_cfg_x=io_dpath_pmp_5_cfg_x; 
  assign io_requestor_0_pmp_5_cfg_w=io_dpath_pmp_5_cfg_w; 
  assign io_requestor_0_pmp_5_cfg_r=io_dpath_pmp_5_cfg_r; 
  assign io_requestor_0_pmp_5_addr=io_dpath_pmp_5_addr; 
  assign io_requestor_0_pmp_5_mask=io_dpath_pmp_5_mask; 
  assign io_requestor_0_pmp_6_cfg_l=io_dpath_pmp_6_cfg_l; 
  assign io_requestor_0_pmp_6_cfg_a=io_dpath_pmp_6_cfg_a; 
  assign io_requestor_0_pmp_6_cfg_x=io_dpath_pmp_6_cfg_x; 
  assign io_requestor_0_pmp_6_cfg_w=io_dpath_pmp_6_cfg_w; 
  assign io_requestor_0_pmp_6_cfg_r=io_dpath_pmp_6_cfg_r; 
  assign io_requestor_0_pmp_6_addr=io_dpath_pmp_6_addr; 
  assign io_requestor_0_pmp_6_mask=io_dpath_pmp_6_mask; 
  assign io_requestor_0_pmp_7_cfg_l=io_dpath_pmp_7_cfg_l; 
  assign io_requestor_0_pmp_7_cfg_a=io_dpath_pmp_7_cfg_a; 
  assign io_requestor_0_pmp_7_cfg_x=io_dpath_pmp_7_cfg_x; 
  assign io_requestor_0_pmp_7_cfg_w=io_dpath_pmp_7_cfg_w; 
  assign io_requestor_0_pmp_7_cfg_r=io_dpath_pmp_7_cfg_r; 
  assign io_requestor_0_pmp_7_addr=io_dpath_pmp_7_addr; 
  assign io_requestor_0_pmp_7_mask=io_dpath_pmp_7_mask; 
  assign io_requestor_1_req_ready=arb_io_in_1_ready; 
  assign io_requestor_1_resp_valid=resp_valid_1; 
  assign io_requestor_1_resp_bits_ae=resp_ae; 
  assign io_requestor_1_resp_bits_pte_ppn=r_pte_ppn; 
  assign io_requestor_1_resp_bits_pte_d=r_pte_d; 
  assign io_requestor_1_resp_bits_pte_a=r_pte_a; 
  assign io_requestor_1_resp_bits_pte_g=r_pte_g; 
  assign io_requestor_1_resp_bits_pte_u=r_pte_u; 
  assign io_requestor_1_resp_bits_pte_x=r_pte_x; 
  assign io_requestor_1_resp_bits_pte_w=r_pte_w; 
  assign io_requestor_1_resp_bits_pte_r=r_pte_r; 
  assign io_requestor_1_resp_bits_pte_v=r_pte_v; 
  assign io_requestor_1_resp_bits_level=count; 
  assign io_requestor_1_resp_bits_homogeneous=pmaHomogeneous&pmpHomogeneous; 
  assign io_requestor_1_ptbr_mode=io_dpath_ptbr_mode; 
  assign io_requestor_1_status_debug=io_dpath_status_debug; 
  assign io_requestor_1_status_prv=io_dpath_status_prv; 
  assign io_requestor_1_pmp_0_cfg_l=io_dpath_pmp_0_cfg_l; 
  assign io_requestor_1_pmp_0_cfg_a=io_dpath_pmp_0_cfg_a; 
  assign io_requestor_1_pmp_0_cfg_x=io_dpath_pmp_0_cfg_x; 
  assign io_requestor_1_pmp_0_cfg_w=io_dpath_pmp_0_cfg_w; 
  assign io_requestor_1_pmp_0_cfg_r=io_dpath_pmp_0_cfg_r; 
  assign io_requestor_1_pmp_0_addr=io_dpath_pmp_0_addr; 
  assign io_requestor_1_pmp_0_mask=io_dpath_pmp_0_mask; 
  assign io_requestor_1_pmp_1_cfg_l=io_dpath_pmp_1_cfg_l; 
  assign io_requestor_1_pmp_1_cfg_a=io_dpath_pmp_1_cfg_a; 
  assign io_requestor_1_pmp_1_cfg_x=io_dpath_pmp_1_cfg_x; 
  assign io_requestor_1_pmp_1_cfg_w=io_dpath_pmp_1_cfg_w; 
  assign io_requestor_1_pmp_1_cfg_r=io_dpath_pmp_1_cfg_r; 
  assign io_requestor_1_pmp_1_addr=io_dpath_pmp_1_addr; 
  assign io_requestor_1_pmp_1_mask=io_dpath_pmp_1_mask; 
  assign io_requestor_1_pmp_2_cfg_l=io_dpath_pmp_2_cfg_l; 
  assign io_requestor_1_pmp_2_cfg_a=io_dpath_pmp_2_cfg_a; 
  assign io_requestor_1_pmp_2_cfg_x=io_dpath_pmp_2_cfg_x; 
  assign io_requestor_1_pmp_2_cfg_w=io_dpath_pmp_2_cfg_w; 
  assign io_requestor_1_pmp_2_cfg_r=io_dpath_pmp_2_cfg_r; 
  assign io_requestor_1_pmp_2_addr=io_dpath_pmp_2_addr; 
  assign io_requestor_1_pmp_2_mask=io_dpath_pmp_2_mask; 
  assign io_requestor_1_pmp_3_cfg_l=io_dpath_pmp_3_cfg_l; 
  assign io_requestor_1_pmp_3_cfg_a=io_dpath_pmp_3_cfg_a; 
  assign io_requestor_1_pmp_3_cfg_x=io_dpath_pmp_3_cfg_x; 
  assign io_requestor_1_pmp_3_cfg_w=io_dpath_pmp_3_cfg_w; 
  assign io_requestor_1_pmp_3_cfg_r=io_dpath_pmp_3_cfg_r; 
  assign io_requestor_1_pmp_3_addr=io_dpath_pmp_3_addr; 
  assign io_requestor_1_pmp_3_mask=io_dpath_pmp_3_mask; 
  assign io_requestor_1_pmp_4_cfg_l=io_dpath_pmp_4_cfg_l; 
  assign io_requestor_1_pmp_4_cfg_a=io_dpath_pmp_4_cfg_a; 
  assign io_requestor_1_pmp_4_cfg_x=io_dpath_pmp_4_cfg_x; 
  assign io_requestor_1_pmp_4_cfg_w=io_dpath_pmp_4_cfg_w; 
  assign io_requestor_1_pmp_4_cfg_r=io_dpath_pmp_4_cfg_r; 
  assign io_requestor_1_pmp_4_addr=io_dpath_pmp_4_addr; 
  assign io_requestor_1_pmp_4_mask=io_dpath_pmp_4_mask; 
  assign io_requestor_1_pmp_5_cfg_l=io_dpath_pmp_5_cfg_l; 
  assign io_requestor_1_pmp_5_cfg_a=io_dpath_pmp_5_cfg_a; 
  assign io_requestor_1_pmp_5_cfg_x=io_dpath_pmp_5_cfg_x; 
  assign io_requestor_1_pmp_5_cfg_w=io_dpath_pmp_5_cfg_w; 
  assign io_requestor_1_pmp_5_cfg_r=io_dpath_pmp_5_cfg_r; 
  assign io_requestor_1_pmp_5_addr=io_dpath_pmp_5_addr; 
  assign io_requestor_1_pmp_5_mask=io_dpath_pmp_5_mask; 
  assign io_requestor_1_pmp_6_cfg_l=io_dpath_pmp_6_cfg_l; 
  assign io_requestor_1_pmp_6_cfg_a=io_dpath_pmp_6_cfg_a; 
  assign io_requestor_1_pmp_6_cfg_x=io_dpath_pmp_6_cfg_x; 
  assign io_requestor_1_pmp_6_cfg_w=io_dpath_pmp_6_cfg_w; 
  assign io_requestor_1_pmp_6_cfg_r=io_dpath_pmp_6_cfg_r; 
  assign io_requestor_1_pmp_6_addr=io_dpath_pmp_6_addr; 
  assign io_requestor_1_pmp_6_mask=io_dpath_pmp_6_mask; 
  assign io_requestor_1_pmp_7_cfg_l=io_dpath_pmp_7_cfg_l; 
  assign io_requestor_1_pmp_7_cfg_a=io_dpath_pmp_7_cfg_a; 
  assign io_requestor_1_pmp_7_cfg_x=io_dpath_pmp_7_cfg_x; 
  assign io_requestor_1_pmp_7_cfg_w=io_dpath_pmp_7_cfg_w; 
  assign io_requestor_1_pmp_7_cfg_r=io_dpath_pmp_7_cfg_r; 
  assign io_requestor_1_pmp_7_addr=io_dpath_pmp_7_addr; 
  assign io_requestor_1_pmp_7_mask=io_dpath_pmp_7_mask; 
  assign io_requestor_1_customCSRs_csrs_0_value=io_dpath_customCSRs_csrs_0_value; 
  assign io_mem_req_valid=_T_55|_io_mem_req_valid_T_1; 
  assign io_mem_req_bits_addr=pte_addr[39:0]; 
  assign io_mem_s1_kill=state!=3'h2; 
  assign io_dpath_perf_l2hit=1'h0; 
  assign io_dpath_perf_pte_miss=_T_100 ? 1'h0:_GEN_77; 
  assign io_dpath_perf_pte_hit=_io_dpath_perf_pte_hit_T_1&~io_dpath_perf_l2hit; 
  assign arb_io_in_0_valid=io_requestor_0_req_valid; 
  assign arb_io_in_0_bits_bits_addr=io_requestor_0_req_bits_bits_addr; 
  assign arb_io_in_1_valid=io_requestor_1_req_valid; 
  assign arb_io_in_1_bits_valid=io_requestor_1_req_bits_valid; 
  assign arb_io_in_1_bits_bits_addr=io_requestor_1_req_bits_bits_addr; 
  assign arb_io_out_ready=_arb_io_out_ready_T&~l2_refill; 
  assign state_barrier_io_x=io_mem_s2_nack ? 3'h1:_GEN_108; 
  assign r_pte_barrier_io_x_ppn=mem_resp_valid ? res_ppn:_r_pte_T_10_ppn; 
  assign r_pte_barrier_io_x_d=mem_resp_valid ? tmp_d:_r_pte_T_10_d; 
  assign r_pte_barrier_io_x_a=mem_resp_valid ? tmp_a:_r_pte_T_10_a; 
  assign r_pte_barrier_io_x_g=mem_resp_valid ? tmp_g:_r_pte_T_10_g; 
  assign r_pte_barrier_io_x_u=mem_resp_valid ? tmp_u:_r_pte_T_10_u; 
  assign r_pte_barrier_io_x_x=mem_resp_valid ? tmp_x:_r_pte_T_10_x; 
  assign r_pte_barrier_io_x_w=mem_resp_valid ? tmp_w:_r_pte_T_10_w; 
  assign r_pte_barrier_io_x_r=mem_resp_valid ? tmp_r:_r_pte_T_10_r; 
  assign r_pte_barrier_io_x_v=mem_resp_valid ? res_v:_r_pte_T_10_v; 
  assign PTW_cov_read_addr=PTW_state; 
  assign PTW_cov_read_data=PTW_cov[PTW_cov_read_addr]; 
  assign PTW_cov_write_data=1'h1; 
  assign PTW_cov_write_addr=PTW_state; 
  assign PTW_cov_write_mask=1'h1; 
  assign PTW_cov_write_en=1'h1; 
  assign valid_shl={valid,3'h0}; 
  assign valid_pad={9'h0,valid_shl}; 
  assign count_shl={count,16'h0}; 
  assign count_pad={2'h0,count_shl}; 
  assign state_reg_shl={state_reg,2'h0}; 
  assign state_reg_pad={11'h0,state_reg_shl}; 
  assign mem_resp_valid_shl={mem_resp_valid,6'h0}; 
  assign mem_resp_valid_pad={13'h0,mem_resp_valid_shl}; 
  assign state_shl={state,7'h0}; 
  assign state_pad={10'h0,state_shl}; 
  assign invalidated_shl={invalidated,13'h0}; 
  assign invalidated_pad={6'h0,invalidated_shl}; 
  assign PTW_xor4=count_pad^state_reg_pad; 
  assign PTW_xor1=valid_pad^PTW_xor4; 
  assign PTW_xor6=state_pad^invalidated_pad; 
  assign PTW_xor2=mem_resp_valid_pad^PTW_xor6; 
  assign PTW_xor0=PTW_xor1^PTW_xor2; 
  assign arb_sum=PTW_covSum+arb_io_covSum; 
  assign state_barrier_sum=arb_sum+state_barrier_io_covSum; 
  assign r_pte_barrier_sum=state_barrier_sum+r_pte_barrier_io_covSum; 
  assign io_covSum=r_pte_barrier_sum; 
  assign stopEn0=~_T_98; 
  assign stopEn1=mem_resp_valid&~_T_123; 
  assign stopEn2=io_mem_s2_nack&~_T_133; 
  assign arb_metaAssert_wire=arb_metaAssert; 
  assign state_barrier_metaAssert_wire=state_barrier_metaAssert; 
  assign r_pte_barrier_metaAssert_wire=r_pte_barrier_metaAssert; 
  assign PTW_or4=stopEn1|stopEn2; 
  assign PTW_or1=stopEn0|PTW_or4; 
  assign PTW_or6=state_barrier_metaAssert_wire|r_pte_barrier_metaAssert_wire; 
  assign PTW_or2=arb_metaAssert_wire|PTW_or6; 
  assign PTW_or0=PTW_or1|PTW_or2; 
  assign metaAssert=PTW_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              state <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 state <=3'h0;
               end 
             else 
               begin 
                 state <=state_barrier_io_y;
               end 
         if (metaReset)
            begin 
              l2_refill <=1'h0;
            end 
          else 
            begin 
              l2_refill <=mem_resp_valid&_GEN_104;
            end 
         if (metaReset)
            begin 
              resp_valid_0 <=1'h0;
            end 
          else 
            if (mem_resp_valid)
               begin 
                 if (traverse)
                    begin 
                      if (_T_100)
                         begin 
                           resp_valid_0 <=1'h0;
                         end 
                       else 
                         if (_T_102)
                            begin 
                              resp_valid_0 <=1'h0;
                            end 
                          else 
                            if (_T_103)
                               begin 
                                 resp_valid_0 <=1'h0;
                               end 
                             else 
                               if (_T_104)
                                  begin 
                                    resp_valid_0 <=_GEN_48;
                                  end 
                                else 
                                  begin 
                                    resp_valid_0 <=_GEN_55;
                                  end 
                    end 
                  else 
                    begin 
                      resp_valid_0 <=_GEN_90;
                    end 
               end 
             else 
               if (_T_100)
                  begin 
                    resp_valid_0 <=1'h0;
                  end 
                else 
                  if (_T_102)
                     begin 
                       resp_valid_0 <=1'h0;
                     end 
                   else 
                     if (_T_103)
                        begin 
                          resp_valid_0 <=1'h0;
                        end 
                      else 
                        if (_T_104)
                           begin 
                             resp_valid_0 <=_GEN_48;
                           end 
                         else 
                           begin 
                             resp_valid_0 <=_GEN_55;
                           end 
         if (metaReset)
            begin 
              resp_valid_1 <=1'h0;
            end 
          else 
            if (mem_resp_valid)
               begin 
                 if (traverse)
                    begin 
                      if (_T_100)
                         begin 
                           resp_valid_1 <=1'h0;
                         end 
                       else 
                         if (_T_102)
                            begin 
                              resp_valid_1 <=1'h0;
                            end 
                          else 
                            if (_T_103)
                               begin 
                                 resp_valid_1 <=1'h0;
                               end 
                             else 
                               if (_T_104)
                                  begin 
                                    resp_valid_1 <=_GEN_49;
                                  end 
                                else 
                                  begin 
                                    resp_valid_1 <=_GEN_56;
                                  end 
                    end 
                  else 
                    begin 
                      resp_valid_1 <=_GEN_91;
                    end 
               end 
             else 
               if (_T_100)
                  begin 
                    resp_valid_1 <=1'h0;
                  end 
                else 
                  if (_T_102)
                     begin 
                       resp_valid_1 <=1'h0;
                     end 
                   else 
                     if (_T_103)
                        begin 
                          resp_valid_1 <=1'h0;
                        end 
                      else 
                        if (_T_104)
                           begin 
                             resp_valid_1 <=_GEN_49;
                           end 
                         else 
                           begin 
                             resp_valid_1 <=_GEN_56;
                           end 
         if (metaReset)
            begin 
              invalidated <=1'h0;
            end 
          else 
            begin 
              invalidated <=io_dpath_sfence_valid|_invalidated_T_1;
            end 
         if (metaReset)
            begin 
              count <=2'h0;
            end 
          else 
            if (mem_resp_valid)
               begin 
                 if (traverse)
                    begin 
                      count <=_count_T_3;
                    end 
                  else 
                    if (_T_100)
                       begin 
                         count <={1'b0,_count_T_1};
                       end 
                     else 
                       if (_T_102)
                          begin 
                            if (pte_cache_hit)
                               begin 
                                 count <=_count_T_3;
                               end 
                          end 
                        else 
                          if (!(_T_103))
                             begin 
                               if (!(_T_104))
                                  begin 
                                    if (_T_107)
                                       begin 
                                         if (~homogeneous)
                                            begin 
                                              count <=2'h2;
                                            end 
                                       end 
                                  end 
                             end 
               end 
             else 
               if (_T_100)
                  begin 
                    count <={1'b0,_count_T_1};
                  end 
                else 
                  if (_T_102)
                     begin 
                       if (pte_cache_hit)
                          begin 
                            count <=_count_T_3;
                          end 
                     end 
                   else 
                     if (!(_T_103))
                        begin 
                          if (!(_T_104))
                             begin 
                               if (_T_107)
                                  begin 
                                    if (~homogeneous)
                                       begin 
                                         count <=2'h2;
                                       end 
                                  end 
                             end 
                        end 
         if (metaReset)
            begin 
              resp_ae <=1'h0;
            end 
          else 
            if (mem_resp_valid)
               begin 
                 if (traverse)
                    begin 
                      if (_T_100)
                         begin 
                           resp_ae <=1'h0;
                         end 
                       else 
                         if (_T_102)
                            begin 
                              resp_ae <=1'h0;
                            end 
                          else 
                            if (_T_103)
                               begin 
                                 resp_ae <=1'h0;
                               end 
                             else 
                               begin 
                                 resp_ae <=_GEN_62;
                               end 
                    end 
                  else 
                    begin 
                      resp_ae <=ae;
                    end 
               end 
             else 
               if (_T_100)
                  begin 
                    resp_ae <=1'h0;
                  end 
                else 
                  if (_T_102)
                     begin 
                       resp_ae <=1'h0;
                     end 
                   else 
                     if (_T_103)
                        begin 
                          resp_ae <=1'h0;
                        end 
                      else 
                        begin 
                          resp_ae <=_GEN_62;
                        end 
         if (metaReset)
            begin 
              r_req_addr <=27'h0;
            end 
          else 
            if (_T_22)
               begin 
                 r_req_addr <=arb_io_out_bits_bits_addr;
               end 
         if (metaReset)
            begin 
              r_req_dest <=1'h0;
            end 
          else 
            if (_T_22)
               begin 
                 r_req_dest <=arb_io_chosen;
               end 
         if (metaReset)
            begin 
              r_pte_ppn <=54'h0;
            end 
          else 
            begin 
              r_pte_ppn <=r_pte_barrier_io_y_ppn;
            end 
         if (metaReset)
            begin 
              r_pte_d <=1'h0;
            end 
          else 
            begin 
              r_pte_d <=r_pte_barrier_io_y_d;
            end 
         if (metaReset)
            begin 
              r_pte_a <=1'h0;
            end 
          else 
            begin 
              r_pte_a <=r_pte_barrier_io_y_a;
            end 
         if (metaReset)
            begin 
              r_pte_g <=1'h0;
            end 
          else 
            begin 
              r_pte_g <=r_pte_barrier_io_y_g;
            end 
         if (metaReset)
            begin 
              r_pte_u <=1'h0;
            end 
          else 
            begin 
              r_pte_u <=r_pte_barrier_io_y_u;
            end 
         if (metaReset)
            begin 
              r_pte_x <=1'h0;
            end 
          else 
            begin 
              r_pte_x <=r_pte_barrier_io_y_x;
            end 
         if (metaReset)
            begin 
              r_pte_w <=1'h0;
            end 
          else 
            begin 
              r_pte_w <=r_pte_barrier_io_y_w;
            end 
         if (metaReset)
            begin 
              r_pte_r <=1'h0;
            end 
          else 
            begin 
              r_pte_r <=r_pte_barrier_io_y_r;
            end 
         if (metaReset)
            begin 
              r_pte_v <=1'h0;
            end 
          else 
            begin 
              r_pte_v <=r_pte_barrier_io_y_v;
            end 
         if (metaReset)
            begin 
              mem_resp_valid <=1'h0;
            end 
          else 
            begin 
              mem_resp_valid <=io_mem_resp_valid;
            end 
         if (metaReset)
            begin 
              mem_resp_data <=64'h0;
            end 
          else 
            begin 
              mem_resp_data <=io_mem_resp_bits_data;
            end 
         if (metaReset)
            begin 
              state_reg <=7'h0;
            end 
          else 
            if (reset)
               begin 
                 state_reg <=7'h0;
               end 
             else 
               if (_T_56)
                  begin 
                    state_reg <=_state_reg_T_16;
                  end 
         if (metaReset)
            begin 
              valid <=8'h0;
            end 
          else 
            if (reset)
               begin 
                 valid <=8'h0;
               end 
             else 
               if (_T_61)
                  begin 
                    valid <=8'h0;
                  end 
                else 
                  if (_T_28)
                     begin 
                       valid <=_T_54;
                     end 
         if (metaReset)
            begin 
              tags_0 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h0==r)
                    begin 
                      tags_0 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              tags_1 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h1==r)
                    begin 
                      tags_1 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              tags_2 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h2==r)
                    begin 
                      tags_2 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              tags_3 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h3==r)
                    begin 
                      tags_3 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              tags_4 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h4==r)
                    begin 
                      tags_4 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              tags_5 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h5==r)
                    begin 
                      tags_5 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              tags_6 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h6==r)
                    begin 
                      tags_6 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              tags_7 <=32'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h7==r)
                    begin 
                      tags_7 <=pte_addr[31:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_0 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h0==r)
                    begin 
                      data_0 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_1 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h1==r)
                    begin 
                      data_1 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_2 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h2==r)
                    begin 
                      data_2 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_3 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h3==r)
                    begin 
                      data_3 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_4 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h4==r)
                    begin 
                      data_4 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_5 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h5==r)
                    begin 
                      data_5 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_6 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h6==r)
                    begin 
                      data_6 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              data_7 <=20'h0;
            end 
          else 
            if (_T_28)
               begin 
                 if (3'h7==r)
                    begin 
                      data_7 <=res_ppn[19:0];
                    end 
               end 
         if (metaReset)
            begin 
              pte_hit <=1'h0;
            end 
          else 
            if (_T_100)
               begin 
                 pte_hit <=1'h0;
               end 
             else 
               begin 
                 pte_hit <=_GEN_75;
               end 
         if (~_T_98)
            begin $display("Assertion failed: PTE Cache Hit/Miss Performance Monitor Events are lower priority than L2TLB Hit event\n    at PTW.scala:198 assert(!(io.dpath.perf.l2hit && (io.dpath.perf.pte_miss || io.dpath.perf.pte_hit)),\n");
            end 
         if (~_T_98)
            begin $display("fatal");
            end 
         if (mem_resp_valid&~_T_123)
            begin $display("Assertion failed\n    at PTW.scala:389 assert(state === s_wait3)\n");
            end 
         if (mem_resp_valid&~_T_123)
            begin $display("fatal");
            end 
         if (io_mem_s2_nack&~_T_133)
            begin $display("Assertion failed\n    at PTW.scala:406 assert(state === s_wait2)\n");
            end 
         if (io_mem_s2_nack&~_T_133)
            begin $display("fatal");
            end 
         PTW_state <=PTW_xor0;
         if (!(PTW_cov_read_data))
            begin 
              PTW_covSum <=PTW_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              PTW_metaAssert <=1'h0;
            end 
          else 
            begin 
              PTW_metaAssert <=PTW_metaAssert|PTW_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (PTW_cov_write_en&PTW_cov_write_mask)
            begin 
              PTW_cov [PTW_cov_write_addr]<=PTW_cov_write_data;
            end 
       end
  
endmodule
 
module Rocket (
  input clock,
  input reset,
  input io_hartid,
  input io_interrupts_debug,
  input io_interrupts_mtip,
  input io_interrupts_msip,
  input io_interrupts_meip,
  input io_interrupts_seip,
  output io_imem_might_request,
  output io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output io_imem_req_bits_speculative,
  output io_imem_sfence_valid,
  output io_imem_sfence_bits_rs1,
  output io_imem_sfence_bits_rs2,
  output [38:0] io_imem_sfence_bits_addr,
  output io_imem_resp_ready,
  input io_imem_resp_valid,
  input io_imem_resp_bits_btb_taken,
  input io_imem_resp_bits_btb_bridx,
  input [4:0] io_imem_resp_bits_btb_entry,
  input [7:0] io_imem_resp_bits_btb_bht_history,
  input [39:0] io_imem_resp_bits_pc,
  input [31:0] io_imem_resp_bits_data,
  input io_imem_resp_bits_xcpt_pf_inst,
  input io_imem_resp_bits_xcpt_ae_inst,
  input io_imem_resp_bits_replay,
  output io_imem_btb_update_valid,
  output [4:0] io_imem_btb_update_bits_prediction_entry,
  output [38:0] io_imem_btb_update_bits_pc,
  output io_imem_btb_update_bits_isValid,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output [1:0] io_imem_btb_update_bits_cfiType,
  output io_imem_bht_update_valid,
  output [7:0] io_imem_bht_update_bits_prediction_history,
  output [38:0] io_imem_bht_update_bits_pc,
  output io_imem_bht_update_bits_branch,
  output io_imem_bht_update_bits_taken,
  output io_imem_bht_update_bits_mispredict,
  output io_imem_flush_icache,
  input io_dmem_req_ready,
  output io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [6:0] io_dmem_req_bits_tag,
  output [4:0] io_dmem_req_bits_cmd,
  output [1:0] io_dmem_req_bits_size,
  output io_dmem_req_bits_signed,
  output io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data_data,
  input io_dmem_s2_nack,
  input io_dmem_resp_valid,
  input [6:0] io_dmem_resp_bits_tag,
  input [1:0] io_dmem_resp_bits_size,
  input [63:0] io_dmem_resp_bits_data,
  input io_dmem_resp_bits_replay,
  input io_dmem_resp_bits_has_data,
  input [63:0] io_dmem_resp_bits_data_word_bypass,
  input io_dmem_replay_next,
  input io_dmem_s2_xcpt_ma_ld,
  input io_dmem_s2_xcpt_ma_st,
  input io_dmem_s2_xcpt_pf_ld,
  input io_dmem_s2_xcpt_pf_st,
  input io_dmem_s2_xcpt_ae_ld,
  input io_dmem_s2_xcpt_ae_st,
  input io_dmem_ordered,
  input io_dmem_perf_release,
  input io_dmem_perf_grant,
  output [3:0] io_ptw_ptbr_mode,
  output [43:0] io_ptw_ptbr_ppn,
  output io_ptw_sfence_valid,
  output io_ptw_sfence_bits_rs1,
  output io_ptw_status_debug,
  output [1:0] io_ptw_status_dprv,
  output [1:0] io_ptw_status_prv,
  output io_ptw_status_mxr,
  output io_ptw_status_sum,
  output io_ptw_pmp_0_cfg_l,
  output [1:0] io_ptw_pmp_0_cfg_a,
  output io_ptw_pmp_0_cfg_x,
  output io_ptw_pmp_0_cfg_w,
  output io_ptw_pmp_0_cfg_r,
  output [29:0] io_ptw_pmp_0_addr,
  output [31:0] io_ptw_pmp_0_mask,
  output io_ptw_pmp_1_cfg_l,
  output [1:0] io_ptw_pmp_1_cfg_a,
  output io_ptw_pmp_1_cfg_x,
  output io_ptw_pmp_1_cfg_w,
  output io_ptw_pmp_1_cfg_r,
  output [29:0] io_ptw_pmp_1_addr,
  output [31:0] io_ptw_pmp_1_mask,
  output io_ptw_pmp_2_cfg_l,
  output [1:0] io_ptw_pmp_2_cfg_a,
  output io_ptw_pmp_2_cfg_x,
  output io_ptw_pmp_2_cfg_w,
  output io_ptw_pmp_2_cfg_r,
  output [29:0] io_ptw_pmp_2_addr,
  output [31:0] io_ptw_pmp_2_mask,
  output io_ptw_pmp_3_cfg_l,
  output [1:0] io_ptw_pmp_3_cfg_a,
  output io_ptw_pmp_3_cfg_x,
  output io_ptw_pmp_3_cfg_w,
  output io_ptw_pmp_3_cfg_r,
  output [29:0] io_ptw_pmp_3_addr,
  output [31:0] io_ptw_pmp_3_mask,
  output io_ptw_pmp_4_cfg_l,
  output [1:0] io_ptw_pmp_4_cfg_a,
  output io_ptw_pmp_4_cfg_x,
  output io_ptw_pmp_4_cfg_w,
  output io_ptw_pmp_4_cfg_r,
  output [29:0] io_ptw_pmp_4_addr,
  output [31:0] io_ptw_pmp_4_mask,
  output io_ptw_pmp_5_cfg_l,
  output [1:0] io_ptw_pmp_5_cfg_a,
  output io_ptw_pmp_5_cfg_x,
  output io_ptw_pmp_5_cfg_w,
  output io_ptw_pmp_5_cfg_r,
  output [29:0] io_ptw_pmp_5_addr,
  output [31:0] io_ptw_pmp_5_mask,
  output io_ptw_pmp_6_cfg_l,
  output [1:0] io_ptw_pmp_6_cfg_a,
  output io_ptw_pmp_6_cfg_x,
  output io_ptw_pmp_6_cfg_w,
  output io_ptw_pmp_6_cfg_r,
  output [29:0] io_ptw_pmp_6_addr,
  output [31:0] io_ptw_pmp_6_mask,
  output io_ptw_pmp_7_cfg_l,
  output [1:0] io_ptw_pmp_7_cfg_a,
  output io_ptw_pmp_7_cfg_x,
  output io_ptw_pmp_7_cfg_w,
  output io_ptw_pmp_7_cfg_r,
  output [29:0] io_ptw_pmp_7_addr,
  output [31:0] io_ptw_pmp_7_mask,
  output [63:0] io_ptw_customCSRs_csrs_0_value,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0] io_fpu_fcsr_rm,
  input io_fpu_fcsr_flags_valid,
  input [4:0] io_fpu_fcsr_flags_bits,
  input [63:0] io_fpu_store_data,
  input [63:0] io_fpu_toint_data,
  output io_fpu_dmem_resp_val,
  output [2:0] io_fpu_dmem_resp_type,
  output [4:0] io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output io_fpu_valid,
  input io_fpu_fcsr_rdy,
  input io_fpu_nack_mem,
  input io_fpu_illegal_rm,
  output io_fpu_killx,
  output io_fpu_killm,
  input io_fpu_dec_wen,
  input io_fpu_dec_ren1,
  input io_fpu_dec_ren2,
  input io_fpu_dec_ren3,
  input io_fpu_sboard_set,
  input io_fpu_sboard_clr,
  input [4:0] io_fpu_sboard_clra,
  output io_trace_0_valid,
  output [39:0] io_trace_0_iaddr,
  output [31:0] io_trace_0_insn,
  output [2:0] io_trace_0_priv,
  output io_trace_0_exception,
  output io_trace_0_interrupt,
  output [63:0] io_trace_0_cause,
  output [39:0] io_trace_0_tval,
  output io_wfi,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input PlusArgTimeout_halt,
  input csr_halt,
  input ibuf_halt,
  input div_halt) ; 
   wire ibuf_clock ;  
   wire ibuf_reset ;  
   wire ibuf_io_imem_ready ;  
   wire ibuf_io_imem_valid ;  
   wire ibuf_io_imem_bits_btb_taken ;  
   wire ibuf_io_imem_bits_btb_bridx ;  
   wire [4:0] ibuf_io_imem_bits_btb_entry ;  
   wire [7:0] ibuf_io_imem_bits_btb_bht_history ;  
   wire [39:0] ibuf_io_imem_bits_pc ;  
   wire [31:0] ibuf_io_imem_bits_data ;  
   wire ibuf_io_imem_bits_xcpt_pf_inst ;  
   wire ibuf_io_imem_bits_xcpt_ae_inst ;  
   wire ibuf_io_imem_bits_replay ;  
   wire ibuf_io_kill ;  
   wire [39:0] ibuf_io_pc ;  
   wire [4:0] ibuf_io_btb_resp_entry ;  
   wire [7:0] ibuf_io_btb_resp_bht_history ;  
   wire ibuf_io_inst_0_ready ;  
   wire ibuf_io_inst_0_valid ;  
   wire ibuf_io_inst_0_bits_xcpt0_pf_inst ;  
   wire ibuf_io_inst_0_bits_xcpt0_ae_inst ;  
   wire ibuf_io_inst_0_bits_xcpt1_pf_inst ;  
   wire ibuf_io_inst_0_bits_xcpt1_ae_inst ;  
   wire ibuf_io_inst_0_bits_replay ;  
   wire ibuf_io_inst_0_bits_rvc ;  
   wire [31:0] ibuf_io_inst_0_bits_inst_bits ;  
   wire [4:0] ibuf_io_inst_0_bits_inst_rd ;  
   wire [4:0] ibuf_io_inst_0_bits_inst_rs1 ;  
   wire [4:0] ibuf_io_inst_0_bits_inst_rs2 ;  
   wire [4:0] ibuf_io_inst_0_bits_inst_rs3 ;  
   wire [31:0] ibuf_io_inst_0_bits_raw ;  
   wire [29:0] ibuf_io_covSum ;  
   wire ibuf_metaAssert ;  
   wire ibuf_metaReset ;  
   reg [63:0] rf[0:30] ;  
   reg [63:0] _RAND_0 ;  
   wire [63:0] rf_id_rs_MPORT_data ;  
   wire [4:0] rf_id_rs_MPORT_addr ;  
   reg [63:0] _RAND_1 ;  
   wire [63:0] rf_id_rs_MPORT_1_data ;  
   wire [4:0] rf_id_rs_MPORT_1_addr ;  
   reg [63:0] _RAND_2 ;  
   wire [63:0] rf_MPORT_data ;  
   wire [4:0] rf_MPORT_addr ;  
   wire rf_MPORT_mask ;  
   wire rf_MPORT_en ;  
   wire csr_clock ;  
   wire csr_reset ;  
   wire csr_io_ungated_clock ;  
   wire csr_io_interrupts_debug ;  
   wire csr_io_interrupts_mtip ;  
   wire csr_io_interrupts_msip ;  
   wire csr_io_interrupts_meip ;  
   wire csr_io_interrupts_seip ;  
   wire csr_io_hartid ;  
   wire [11:0] csr_io_rw_addr ;  
   wire [2:0] csr_io_rw_cmd ;  
   wire [63:0] csr_io_rw_rdata ;  
   wire [63:0] csr_io_rw_wdata ;  
   wire [11:0] csr_io_decode_0_csr ;  
   wire csr_io_decode_0_fp_illegal ;  
   wire csr_io_decode_0_fp_csr ;  
   wire csr_io_decode_0_read_illegal ;  
   wire csr_io_decode_0_write_illegal ;  
   wire csr_io_decode_0_write_flush ;  
   wire csr_io_decode_0_system_illegal ;  
   wire csr_io_csr_stall ;  
   wire csr_io_eret ;  
   wire csr_io_singleStep ;  
   wire csr_io_status_debug ;  
   wire csr_io_status_cease ;  
   wire csr_io_status_wfi ;  
   wire [31:0] csr_io_status_isa ;  
   wire [1:0] csr_io_status_dprv ;  
   wire [1:0] csr_io_status_prv ;  
   wire csr_io_status_sd ;  
   wire [26:0] csr_io_status_zero2 ;  
   wire [1:0] csr_io_status_sxl ;  
   wire [1:0] csr_io_status_uxl ;  
   wire csr_io_status_sd_rv32 ;  
   wire [7:0] csr_io_status_zero1 ;  
   wire csr_io_status_tsr ;  
   wire csr_io_status_tw ;  
   wire csr_io_status_tvm ;  
   wire csr_io_status_mxr ;  
   wire csr_io_status_sum ;  
   wire csr_io_status_mprv ;  
   wire [1:0] csr_io_status_xs ;  
   wire [1:0] csr_io_status_fs ;  
   wire [1:0] csr_io_status_mpp ;  
   wire [1:0] csr_io_status_vs ;  
   wire csr_io_status_spp ;  
   wire csr_io_status_mpie ;  
   wire csr_io_status_hpie ;  
   wire csr_io_status_spie ;  
   wire csr_io_status_upie ;  
   wire csr_io_status_mie ;  
   wire csr_io_status_hie ;  
   wire csr_io_status_sie ;  
   wire csr_io_status_uie ;  
   wire [3:0] csr_io_ptbr_mode ;  
   wire [43:0] csr_io_ptbr_ppn ;  
   wire [39:0] csr_io_evec ;  
   wire csr_io_exception ;  
   wire csr_io_retire ;  
   wire [63:0] csr_io_cause ;  
   wire [39:0] csr_io_pc ;  
   wire [39:0] csr_io_tval ;  
   wire [63:0] csr_io_time ;  
   wire [2:0] csr_io_fcsr_rm ;  
   wire csr_io_fcsr_flags_valid ;  
   wire [4:0] csr_io_fcsr_flags_bits ;  
   wire csr_io_interrupt ;  
   wire [63:0] csr_io_interrupt_cause ;  
   wire csr_io_bp_0_control_action ;  
   wire [1:0] csr_io_bp_0_control_tmatch ;  
   wire csr_io_bp_0_control_m ;  
   wire csr_io_bp_0_control_s ;  
   wire csr_io_bp_0_control_u ;  
   wire csr_io_bp_0_control_x ;  
   wire csr_io_bp_0_control_w ;  
   wire csr_io_bp_0_control_r ;  
   wire [38:0] csr_io_bp_0_address ;  
   wire csr_io_pmp_0_cfg_l ;  
   wire [1:0] csr_io_pmp_0_cfg_a ;  
   wire csr_io_pmp_0_cfg_x ;  
   wire csr_io_pmp_0_cfg_w ;  
   wire csr_io_pmp_0_cfg_r ;  
   wire [29:0] csr_io_pmp_0_addr ;  
   wire [31:0] csr_io_pmp_0_mask ;  
   wire csr_io_pmp_1_cfg_l ;  
   wire [1:0] csr_io_pmp_1_cfg_a ;  
   wire csr_io_pmp_1_cfg_x ;  
   wire csr_io_pmp_1_cfg_w ;  
   wire csr_io_pmp_1_cfg_r ;  
   wire [29:0] csr_io_pmp_1_addr ;  
   wire [31:0] csr_io_pmp_1_mask ;  
   wire csr_io_pmp_2_cfg_l ;  
   wire [1:0] csr_io_pmp_2_cfg_a ;  
   wire csr_io_pmp_2_cfg_x ;  
   wire csr_io_pmp_2_cfg_w ;  
   wire csr_io_pmp_2_cfg_r ;  
   wire [29:0] csr_io_pmp_2_addr ;  
   wire [31:0] csr_io_pmp_2_mask ;  
   wire csr_io_pmp_3_cfg_l ;  
   wire [1:0] csr_io_pmp_3_cfg_a ;  
   wire csr_io_pmp_3_cfg_x ;  
   wire csr_io_pmp_3_cfg_w ;  
   wire csr_io_pmp_3_cfg_r ;  
   wire [29:0] csr_io_pmp_3_addr ;  
   wire [31:0] csr_io_pmp_3_mask ;  
   wire csr_io_pmp_4_cfg_l ;  
   wire [1:0] csr_io_pmp_4_cfg_a ;  
   wire csr_io_pmp_4_cfg_x ;  
   wire csr_io_pmp_4_cfg_w ;  
   wire csr_io_pmp_4_cfg_r ;  
   wire [29:0] csr_io_pmp_4_addr ;  
   wire [31:0] csr_io_pmp_4_mask ;  
   wire csr_io_pmp_5_cfg_l ;  
   wire [1:0] csr_io_pmp_5_cfg_a ;  
   wire csr_io_pmp_5_cfg_x ;  
   wire csr_io_pmp_5_cfg_w ;  
   wire csr_io_pmp_5_cfg_r ;  
   wire [29:0] csr_io_pmp_5_addr ;  
   wire [31:0] csr_io_pmp_5_mask ;  
   wire csr_io_pmp_6_cfg_l ;  
   wire [1:0] csr_io_pmp_6_cfg_a ;  
   wire csr_io_pmp_6_cfg_x ;  
   wire csr_io_pmp_6_cfg_w ;  
   wire csr_io_pmp_6_cfg_r ;  
   wire [29:0] csr_io_pmp_6_addr ;  
   wire [31:0] csr_io_pmp_6_mask ;  
   wire csr_io_pmp_7_cfg_l ;  
   wire [1:0] csr_io_pmp_7_cfg_a ;  
   wire csr_io_pmp_7_cfg_x ;  
   wire csr_io_pmp_7_cfg_w ;  
   wire csr_io_pmp_7_cfg_r ;  
   wire [29:0] csr_io_pmp_7_addr ;  
   wire [31:0] csr_io_pmp_7_mask ;  
   wire csr_io_inhibit_cycle ;  
   wire [31:0] csr_io_inst_0 ;  
   wire csr_io_trace_0_valid ;  
   wire [39:0] csr_io_trace_0_iaddr ;  
   wire [31:0] csr_io_trace_0_insn ;  
   wire [2:0] csr_io_trace_0_priv ;  
   wire csr_io_trace_0_exception ;  
   wire csr_io_trace_0_interrupt ;  
   wire [63:0] csr_io_trace_0_cause ;  
   wire [39:0] csr_io_trace_0_tval ;  
   wire [63:0] csr_io_customCSRs_0_value ;  
   wire [29:0] csr_io_covSum ;  
   wire csr_metaAssert ;  
   wire csr_metaReset ;  
   wire bpu_io_status_debug ;  
   wire [1:0] bpu_io_status_prv ;  
   wire bpu_io_bp_0_control_action ;  
   wire [1:0] bpu_io_bp_0_control_tmatch ;  
   wire bpu_io_bp_0_control_m ;  
   wire bpu_io_bp_0_control_s ;  
   wire bpu_io_bp_0_control_u ;  
   wire bpu_io_bp_0_control_x ;  
   wire bpu_io_bp_0_control_w ;  
   wire bpu_io_bp_0_control_r ;  
   wire [38:0] bpu_io_bp_0_address ;  
   wire [38:0] bpu_io_pc ;  
   wire [38:0] bpu_io_ea ;  
   wire bpu_io_xcpt_if ;  
   wire bpu_io_xcpt_ld ;  
   wire bpu_io_xcpt_st ;  
   wire bpu_io_debug_if ;  
   wire bpu_io_debug_ld ;  
   wire bpu_io_debug_st ;  
   wire [29:0] bpu_io_covSum ;  
   wire bpu_metaAssert ;  
   wire alu_io_dw ;  
   wire [3:0] alu_io_fn ;  
   wire [63:0] alu_io_in2 ;  
   wire [63:0] alu_io_in1 ;  
   wire [63:0] alu_io_out ;  
   wire [63:0] alu_io_adder_out ;  
   wire alu_io_cmp_out ;  
   wire [29:0] alu_io_covSum ;  
   wire alu_metaAssert ;  
   wire div_clock ;  
   wire div_reset ;  
   wire div_io_req_ready ;  
   wire div_io_req_valid ;  
   wire [3:0] div_io_req_bits_fn ;  
   wire div_io_req_bits_dw ;  
   wire [63:0] div_io_req_bits_in1 ;  
   wire [63:0] div_io_req_bits_in2 ;  
   wire [4:0] div_io_req_bits_tag ;  
   wire div_io_kill ;  
   wire div_io_resp_ready ;  
   wire div_io_resp_valid ;  
   wire [63:0] div_io_resp_bits_data ;  
   wire [4:0] div_io_resp_bits_tag ;  
   wire [29:0] div_io_covSum ;  
   wire div_metaAssert ;  
   wire div_metaReset ;  
   wire PlusArgTimeout_clock ;  
   wire PlusArgTimeout_reset ;  
   wire [31:0] PlusArgTimeout_io_count ;  
   wire [29:0] PlusArgTimeout_io_covSum ;  
   wire PlusArgTimeout_metaAssert ;  
   wire PlusArgTimeout_metaReset ;  
   reg id_reg_pause ;  
   reg [31:0] _RAND_3 ;  
   reg imem_might_request_reg ;  
   reg [31:0] _RAND_4 ;  
   reg ex_ctrl_fp ;  
   reg [31:0] _RAND_5 ;  
   reg ex_ctrl_branch ;  
   reg [31:0] _RAND_6 ;  
   reg ex_ctrl_jal ;  
   reg [31:0] _RAND_7 ;  
   reg ex_ctrl_jalr ;  
   reg [31:0] _RAND_8 ;  
   reg ex_ctrl_rxs2 ;  
   reg [31:0] _RAND_9 ;  
   reg [1:0] ex_ctrl_sel_alu2 ;  
   reg [31:0] _RAND_10 ;  
   reg [1:0] ex_ctrl_sel_alu1 ;  
   reg [31:0] _RAND_11 ;  
   reg [2:0] ex_ctrl_sel_imm ;  
   reg [31:0] _RAND_12 ;  
   reg ex_ctrl_alu_dw ;  
   reg [31:0] _RAND_13 ;  
   reg [3:0] ex_ctrl_alu_fn ;  
   reg [31:0] _RAND_14 ;  
   reg ex_ctrl_mem ;  
   reg [31:0] _RAND_15 ;  
   reg [4:0] ex_ctrl_mem_cmd ;  
   reg [31:0] _RAND_16 ;  
   reg ex_ctrl_wfd ;  
   reg [31:0] _RAND_17 ;  
   reg ex_ctrl_div ;  
   reg [31:0] _RAND_18 ;  
   reg ex_ctrl_wxd ;  
   reg [31:0] _RAND_19 ;  
   reg [2:0] ex_ctrl_csr ;  
   reg [31:0] _RAND_20 ;  
   reg ex_ctrl_fence_i ;  
   reg [31:0] _RAND_21 ;  
   reg mem_ctrl_fp ;  
   reg [31:0] _RAND_22 ;  
   reg mem_ctrl_branch ;  
   reg [31:0] _RAND_23 ;  
   reg mem_ctrl_jal ;  
   reg [31:0] _RAND_24 ;  
   reg mem_ctrl_jalr ;  
   reg [31:0] _RAND_25 ;  
   reg mem_ctrl_mem ;  
   reg [31:0] _RAND_26 ;  
   reg mem_ctrl_wfd ;  
   reg [31:0] _RAND_27 ;  
   reg mem_ctrl_div ;  
   reg [31:0] _RAND_28 ;  
   reg mem_ctrl_wxd ;  
   reg [31:0] _RAND_29 ;  
   reg [2:0] mem_ctrl_csr ;  
   reg [31:0] _RAND_30 ;  
   reg mem_ctrl_fence_i ;  
   reg [31:0] _RAND_31 ;  
   reg wb_ctrl_mem ;  
   reg [31:0] _RAND_32 ;  
   reg wb_ctrl_wfd ;  
   reg [31:0] _RAND_33 ;  
   reg wb_ctrl_div ;  
   reg [31:0] _RAND_34 ;  
   reg wb_ctrl_wxd ;  
   reg [31:0] _RAND_35 ;  
   reg [2:0] wb_ctrl_csr ;  
   reg [31:0] _RAND_36 ;  
   reg wb_ctrl_fence_i ;  
   reg [31:0] _RAND_37 ;  
   reg ex_reg_xcpt_interrupt ;  
   reg [31:0] _RAND_38 ;  
   reg ex_reg_valid ;  
   reg [31:0] _RAND_39 ;  
   reg ex_reg_rvc ;  
   reg [31:0] _RAND_40 ;  
   reg [4:0] ex_reg_btb_resp_entry ;  
   reg [31:0] _RAND_41 ;  
   reg [7:0] ex_reg_btb_resp_bht_history ;  
   reg [31:0] _RAND_42 ;  
   reg ex_reg_xcpt ;  
   reg [31:0] _RAND_43 ;  
   reg ex_reg_flush_pipe ;  
   reg [31:0] _RAND_44 ;  
   reg ex_reg_load_use ;  
   reg [31:0] _RAND_45 ;  
   reg [63:0] ex_reg_cause ;  
   reg [63:0] _RAND_46 ;  
   reg ex_reg_replay ;  
   reg [31:0] _RAND_47 ;  
   reg [39:0] ex_reg_pc ;  
   reg [63:0] _RAND_48 ;  
   reg [1:0] ex_reg_mem_size ;  
   reg [31:0] _RAND_49 ;  
   reg [31:0] ex_reg_inst ;  
   reg [31:0] _RAND_50 ;  
   reg [31:0] ex_reg_raw_inst ;  
   reg [31:0] _RAND_51 ;  
   reg mem_reg_xcpt_interrupt ;  
   reg [31:0] _RAND_52 ;  
   reg mem_reg_valid ;  
   reg [31:0] _RAND_53 ;  
   reg mem_reg_rvc ;  
   reg [31:0] _RAND_54 ;  
   reg [4:0] mem_reg_btb_resp_entry ;  
   reg [31:0] _RAND_55 ;  
   reg [7:0] mem_reg_btb_resp_bht_history ;  
   reg [31:0] _RAND_56 ;  
   reg mem_reg_xcpt ;  
   reg [31:0] _RAND_57 ;  
   reg mem_reg_replay ;  
   reg [31:0] _RAND_58 ;  
   reg mem_reg_flush_pipe ;  
   reg [31:0] _RAND_59 ;  
   reg [63:0] mem_reg_cause ;  
   reg [63:0] _RAND_60 ;  
   reg mem_reg_slow_bypass ;  
   reg [31:0] _RAND_61 ;  
   reg mem_reg_load ;  
   reg [31:0] _RAND_62 ;  
   reg mem_reg_store ;  
   reg [31:0] _RAND_63 ;  
   reg mem_reg_sfence ;  
   reg [31:0] _RAND_64 ;  
   reg [39:0] mem_reg_pc ;  
   reg [63:0] _RAND_65 ;  
   reg [31:0] mem_reg_inst ;  
   reg [31:0] _RAND_66 ;  
   reg [1:0] mem_reg_mem_size ;  
   reg [31:0] _RAND_67 ;  
   reg [31:0] mem_reg_raw_inst ;  
   reg [31:0] _RAND_68 ;  
   reg [63:0] mem_reg_wdata ;  
   reg [63:0] _RAND_69 ;  
   reg [63:0] mem_reg_rs2 ;  
   reg [63:0] _RAND_70 ;  
   reg mem_br_taken ;  
   reg [31:0] _RAND_71 ;  
   reg wb_reg_valid ;  
   reg [31:0] _RAND_72 ;  
   reg wb_reg_xcpt ;  
   reg [31:0] _RAND_73 ;  
   reg wb_reg_replay ;  
   reg [31:0] _RAND_74 ;  
   reg wb_reg_flush_pipe ;  
   reg [31:0] _RAND_75 ;  
   reg [63:0] wb_reg_cause ;  
   reg [63:0] _RAND_76 ;  
   reg wb_reg_sfence ;  
   reg [31:0] _RAND_77 ;  
   reg [39:0] wb_reg_pc ;  
   reg [63:0] _RAND_78 ;  
   reg [1:0] wb_reg_mem_size ;  
   reg [31:0] _RAND_79 ;  
   reg [31:0] wb_reg_inst ;  
   reg [31:0] _RAND_80 ;  
   reg [31:0] wb_reg_raw_inst ;  
   reg [31:0] _RAND_81 ;  
   reg [63:0] wb_reg_wdata ;  
   reg [63:0] _RAND_82 ;  
   wire replay_wb_common ;  
   wire _T_83 ;  
   wire _T_84 ;  
   wire _T_95 ;  
   wire _T_86 ;  
   wire _T_96 ;  
   wire _T_88 ;  
   wire _T_97 ;  
   wire _T_90 ;  
   wire _T_98 ;  
   wire _T_92 ;  
   wire _T_99 ;  
   wire _T_94 ;  
   wire wb_xcpt ;  
   wire _take_pc_wb_T ;  
   wire _take_pc_wb_T_1 ;  
   wire take_pc_wb ;  
   wire _ex_pc_valid_T ;  
   wire ex_pc_valid ;  
   wire _mem_npc_T ;  
   wire [24:0] a ;  
   wire _mem_npc_msb_T ;  
   wire _mem_npc_msb_T_1 ;  
   wire _mem_npc_msb_T_2 ;  
   wire msb ;  
   wire [38:0] mem_npc_lo ;  
   wire [39:0] _mem_npc_T_2 ;  
   wire _mem_br_target_T_1 ;  
   wire mem_br_target_sign ;  
   wire mem_br_target_hi_hi_hi ;  
   wire [10:0] mem_br_target_hi_hi_lo ;  
   wire [7:0] mem_br_target_hi_lo_hi ;  
   wire mem_br_target_hi_lo_lo ;  
   wire [5:0] mem_br_target_lo_hi_hi ;  
   wire [3:0] mem_br_target_lo_hi_lo ;  
   wire [31:0] _mem_br_target_T_3 ;  
   wire [7:0] mem_br_target_hi_lo_hi_1 ;  
   wire mem_br_target_hi_lo_lo_1 ;  
   wire [31:0] _mem_br_target_T_5 ;  
   wire [3:0] _mem_br_target_T_6 ;  
   wire [31:0] _mem_br_target_T_7 ;  
   wire [31:0] _mem_br_target_T_8 ;  
   wire [39:0] _GEN_248 ;  
   wire [39:0] mem_br_target ;  
   wire [39:0] _mem_npc_T_3 ;  
   wire [39:0] mem_npc ;  
   wire _mem_wrong_npc_T ;  
   wire _mem_wrong_npc_T_1 ;  
   wire _mem_wrong_npc_T_2 ;  
   wire _mem_wrong_npc_T_3 ;  
   wire mem_wrong_npc ;  
   wire _take_pc_mem_T ;  
   wire take_pc_mem ;  
   wire take_pc_mem_wb ;  
   wire [31:0] _id_ctrl_decoder_bit_T ;  
   wire _id_ctrl_decoder_bit_T_1 ;  
   wire _id_ctrl_decoder_bit_T_3 ;  
   wire _id_ctrl_decoder_bit_T_5 ;  
   wire _id_ctrl_decoder_bit_T_7 ;  
   wire _id_ctrl_decoder_bit_T_9 ;  
   wire _id_ctrl_decoder_bit_T_11 ;  
   wire _id_ctrl_decoder_bit_T_13 ;  
   wire _id_ctrl_decoder_bit_T_15 ;  
   wire _id_ctrl_decoder_bit_T_17 ;  
   wire _id_ctrl_decoder_bit_T_19 ;  
   wire _id_ctrl_decoder_bit_T_21 ;  
   wire _id_ctrl_decoder_bit_T_23 ;  
   wire _id_ctrl_decoder_bit_T_25 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_26 ;  
   wire _id_ctrl_decoder_bit_T_27 ;  
   wire _id_ctrl_decoder_bit_T_29 ;  
   wire _id_ctrl_decoder_bit_T_31 ;  
   wire _id_ctrl_decoder_bit_T_33 ;  
   wire _id_ctrl_decoder_bit_T_35 ;  
   wire _id_ctrl_decoder_bit_T_37 ;  
   wire _id_ctrl_decoder_bit_T_39 ;  
   wire _id_ctrl_decoder_bit_T_41 ;  
   wire _id_ctrl_decoder_bit_T_43 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_44 ;  
   wire _id_ctrl_decoder_bit_T_45 ;  
   wire _id_ctrl_decoder_bit_T_47 ;  
   wire _id_ctrl_decoder_bit_T_49 ;  
   wire _id_ctrl_decoder_bit_T_51 ;  
   wire _id_ctrl_decoder_bit_T_53 ;  
   wire _id_ctrl_decoder_bit_T_55 ;  
   wire _id_ctrl_decoder_bit_T_57 ;  
   wire _id_ctrl_decoder_bit_T_59 ;  
   wire _id_ctrl_decoder_bit_T_61 ;  
   wire _id_ctrl_decoder_bit_T_63 ;  
   wire _id_ctrl_decoder_bit_T_65 ;  
   wire _id_ctrl_decoder_bit_T_67 ;  
   wire _id_ctrl_decoder_bit_T_69 ;  
   wire _id_ctrl_decoder_bit_T_71 ;  
   wire _id_ctrl_decoder_bit_T_73 ;  
   wire _id_ctrl_decoder_bit_T_75 ;  
   wire _id_ctrl_decoder_bit_T_77 ;  
   wire _id_ctrl_decoder_bit_T_79 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_80 ;  
   wire _id_ctrl_decoder_bit_T_81 ;  
   wire _id_ctrl_decoder_bit_T_83 ;  
   wire _id_ctrl_decoder_bit_T_85 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_86 ;  
   wire _id_ctrl_decoder_bit_T_87 ;  
   wire _id_ctrl_decoder_bit_T_89 ;  
   wire _id_ctrl_decoder_bit_T_91 ;  
   wire _id_ctrl_decoder_bit_T_93 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_94 ;  
   wire _id_ctrl_decoder_bit_T_95 ;  
   wire _id_ctrl_decoder_bit_T_97 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_98 ;  
   wire _id_ctrl_decoder_bit_T_99 ;  
   wire _id_ctrl_decoder_bit_T_101 ;  
   wire _id_ctrl_decoder_bit_T_103 ;  
   wire _id_ctrl_decoder_bit_T_105 ;  
   wire _id_ctrl_decoder_bit_T_107 ;  
   wire _id_ctrl_decoder_bit_T_109 ;  
   wire _id_ctrl_decoder_bit_T_111 ;  
   wire _id_ctrl_decoder_bit_T_113 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_114 ;  
   wire _id_ctrl_decoder_bit_T_115 ;  
   wire _id_ctrl_decoder_bit_T_117 ;  
   wire _id_ctrl_decoder_bit_T_119 ;  
   wire _id_ctrl_decoder_bit_T_121 ;  
   wire _id_ctrl_decoder_bit_T_123 ;  
   wire _id_ctrl_decoder_bit_T_125 ;  
   wire _id_ctrl_decoder_bit_T_127 ;  
   wire _id_ctrl_decoder_bit_T_129 ;  
   wire _id_ctrl_decoder_bit_T_131 ;  
   wire _id_ctrl_decoder_bit_T_133 ;  
   wire _id_ctrl_decoder_bit_T_135 ;  
   wire _id_ctrl_decoder_bit_T_137 ;  
   wire _id_ctrl_decoder_bit_T_139 ;  
   wire _id_ctrl_decoder_bit_T_141 ;  
   wire _id_ctrl_decoder_bit_T_143 ;  
   wire _id_ctrl_decoder_bit_T_145 ;  
   wire _id_ctrl_decoder_bit_T_147 ;  
   wire _id_ctrl_decoder_bit_T_149 ;  
   wire _id_ctrl_decoder_bit_T_151 ;  
   wire _id_ctrl_decoder_bit_T_153 ;  
   wire _id_ctrl_decoder_bit_T_155 ;  
   wire _id_ctrl_decoder_bit_T_157 ;  
   wire _id_ctrl_decoder_bit_T_159 ;  
   wire _id_ctrl_decoder_bit_T_161 ;  
   wire _id_ctrl_decoder_bit_T_163 ;  
   wire _id_ctrl_decoder_bit_T_165 ;  
   wire _id_ctrl_decoder_bit_T_167 ;  
   wire _id_ctrl_decoder_bit_T_169 ;  
   wire _id_ctrl_decoder_bit_T_171 ;  
   wire _id_ctrl_decoder_bit_T_173 ;  
   wire _id_ctrl_decoder_bit_T_175 ;  
   wire _id_ctrl_decoder_bit_T_177 ;  
   wire _id_ctrl_decoder_bit_T_179 ;  
   wire _id_ctrl_decoder_bit_T_181 ;  
   wire _id_ctrl_decoder_bit_T_183 ;  
   wire _id_ctrl_decoder_bit_T_185 ;  
   wire _id_ctrl_decoder_bit_T_187 ;  
   wire _id_ctrl_decoder_bit_T_189 ;  
   wire _id_ctrl_decoder_bit_T_191 ;  
   wire _id_ctrl_decoder_bit_T_193 ;  
   wire _id_ctrl_decoder_bit_T_195 ;  
   wire _id_ctrl_decoder_bit_T_197 ;  
   wire _id_ctrl_decoder_bit_T_199 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_200 ;  
   wire _id_ctrl_decoder_bit_T_201 ;  
   wire _id_ctrl_decoder_bit_T_203 ;  
   wire _id_ctrl_decoder_bit_T_205 ;  
   wire _id_ctrl_decoder_bit_T_207 ;  
   wire _id_ctrl_decoder_bit_T_209 ;  
   wire _id_ctrl_decoder_bit_T_211 ;  
   wire _id_ctrl_decoder_bit_T_213 ;  
   wire _id_ctrl_decoder_bit_T_215 ;  
   wire _id_ctrl_decoder_bit_T_217 ;  
   wire _id_ctrl_decoder_bit_T_219 ;  
   wire _id_ctrl_decoder_bit_T_221 ;  
   wire _id_ctrl_decoder_bit_T_223 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_224 ;  
   wire _id_ctrl_decoder_bit_T_225 ;  
   wire _id_ctrl_decoder_bit_T_226 ;  
   wire _id_ctrl_decoder_bit_T_227 ;  
   wire _id_ctrl_decoder_bit_T_229 ;  
   wire _id_ctrl_decoder_bit_T_231 ;  
   wire _id_ctrl_decoder_bit_T_233 ;  
   wire _id_ctrl_decoder_bit_T_235 ;  
   wire _id_ctrl_decoder_bit_T_237 ;  
   wire _id_ctrl_decoder_bit_T_239 ;  
   wire _id_ctrl_decoder_bit_T_241 ;  
   wire [31:0] _id_ctrl_decoder_bit_T_242 ;  
   wire _id_ctrl_decoder_bit_T_243 ;  
   wire _id_ctrl_decoder_bit_T_245 ;  
   wire _id_ctrl_decoder_bit_T_247 ;  
   wire _id_ctrl_decoder_bit_T_249 ;  
   wire _id_ctrl_decoder_bit_T_251 ;  
   wire _id_ctrl_decoder_bit_T_253 ;  
   wire _id_ctrl_decoder_bit_T_255 ;  
   wire _id_ctrl_decoder_bit_T_257 ;  
   wire _id_ctrl_decoder_bit_T_259 ;  
   wire _id_ctrl_decoder_bit_T_261 ;  
   wire _id_ctrl_decoder_bit_T_263 ;  
   wire _id_ctrl_decoder_bit_T_265 ;  
   wire _id_ctrl_decoder_bit_T_267 ;  
   wire _id_ctrl_decoder_bit_T_269 ;  
   wire _id_ctrl_decoder_bit_T_271 ;  
   wire _id_ctrl_decoder_bit_T_273 ;  
   wire _id_ctrl_decoder_bit_T_275 ;  
   wire _id_ctrl_decoder_bit_T_277 ;  
   wire _id_ctrl_decoder_bit_T_279 ;  
   wire _id_ctrl_decoder_bit_T_281 ;  
   wire _id_ctrl_decoder_bit_T_283 ;  
   wire _id_ctrl_decoder_bit_T_285 ;  
   wire _id_ctrl_decoder_bit_T_287 ;  
   wire _id_ctrl_decoder_bit_T_289 ;  
   wire _id_ctrl_decoder_bit_T_291 ;  
   wire _id_ctrl_decoder_bit_T_293 ;  
   wire _id_ctrl_decoder_bit_T_295 ;  
   wire _id_ctrl_decoder_bit_T_297 ;  
   wire _id_ctrl_decoder_bit_T_299 ;  
   wire _id_ctrl_decoder_bit_T_300 ;  
   wire _id_ctrl_decoder_bit_T_301 ;  
   wire _id_ctrl_decoder_bit_T_302 ;  
   wire _id_ctrl_decoder_bit_T_303 ;  
   wire _id_ctrl_decoder_bit_T_304 ;  
   wire _id_ctrl_decoder_bit_T_306 ;  
   wire _id_ctrl_decoder_bit_T_308 ;  
   wire _id_ctrl_decoder_bit_T_310 ;  
   wire _id_ctrl_decoder_bit_T_312 ;  
   wire _id_ctrl_decoder_bit_T_314 ;  
   wire _id_ctrl_decoder_bit_T_316 ;  
   wire _id_ctrl_decoder_bit_T_318 ;  
   wire _id_ctrl_decoder_bit_T_319 ;  
   wire _id_ctrl_decoder_bit_T_320 ;  
   wire _id_ctrl_decoder_bit_T_321 ;  
   wire _id_ctrl_decoder_bit_T_322 ;  
   wire _id_ctrl_decoder_bit_T_323 ;  
   wire _id_ctrl_decoder_bit_T_324 ;  
   wire _id_ctrl_decoder_bit_T_325 ;  
   wire _id_ctrl_decoder_bit_T_326 ;  
   wire _id_ctrl_decoder_bit_T_327 ;  
   wire _id_ctrl_decoder_bit_T_328 ;  
   wire _id_ctrl_decoder_bit_T_329 ;  
   wire _id_ctrl_decoder_bit_T_330 ;  
   wire _id_ctrl_decoder_bit_T_331 ;  
   wire _id_ctrl_decoder_bit_T_332 ;  
   wire _id_ctrl_decoder_bit_T_333 ;  
   wire _id_ctrl_decoder_bit_T_334 ;  
   wire _id_ctrl_decoder_bit_T_335 ;  
   wire _id_ctrl_decoder_bit_T_336 ;  
   wire _id_ctrl_decoder_bit_T_337 ;  
   wire _id_ctrl_decoder_bit_T_338 ;  
   wire _id_ctrl_decoder_bit_T_339 ;  
   wire _id_ctrl_decoder_bit_T_340 ;  
   wire _id_ctrl_decoder_bit_T_341 ;  
   wire _id_ctrl_decoder_bit_T_342 ;  
   wire _id_ctrl_decoder_bit_T_343 ;  
   wire _id_ctrl_decoder_bit_T_344 ;  
   wire _id_ctrl_decoder_bit_T_345 ;  
   wire _id_ctrl_decoder_bit_T_346 ;  
   wire _id_ctrl_decoder_bit_T_347 ;  
   wire _id_ctrl_decoder_bit_T_348 ;  
   wire _id_ctrl_decoder_bit_T_349 ;  
   wire _id_ctrl_decoder_bit_T_350 ;  
   wire _id_ctrl_decoder_bit_T_351 ;  
   wire _id_ctrl_decoder_bit_T_352 ;  
   wire _id_ctrl_decoder_bit_T_353 ;  
   wire _id_ctrl_decoder_bit_T_354 ;  
   wire _id_ctrl_decoder_bit_T_355 ;  
   wire _id_ctrl_decoder_bit_T_356 ;  
   wire _id_ctrl_decoder_bit_T_357 ;  
   wire _id_ctrl_decoder_bit_T_358 ;  
   wire _id_ctrl_decoder_bit_T_359 ;  
   wire _id_ctrl_decoder_bit_T_360 ;  
   wire _id_ctrl_decoder_bit_T_361 ;  
   wire _id_ctrl_decoder_bit_T_362 ;  
   wire _id_ctrl_decoder_bit_T_363 ;  
   wire _id_ctrl_decoder_bit_T_364 ;  
   wire _id_ctrl_decoder_bit_T_365 ;  
   wire _id_ctrl_decoder_bit_T_366 ;  
   wire _id_ctrl_decoder_bit_T_367 ;  
   wire _id_ctrl_decoder_bit_T_368 ;  
   wire _id_ctrl_decoder_bit_T_369 ;  
   wire _id_ctrl_decoder_bit_T_370 ;  
   wire _id_ctrl_decoder_bit_T_371 ;  
   wire _id_ctrl_decoder_bit_T_372 ;  
   wire _id_ctrl_decoder_bit_T_373 ;  
   wire _id_ctrl_decoder_bit_T_374 ;  
   wire _id_ctrl_decoder_bit_T_375 ;  
   wire _id_ctrl_decoder_bit_T_376 ;  
   wire _id_ctrl_decoder_bit_T_377 ;  
   wire _id_ctrl_decoder_bit_T_378 ;  
   wire _id_ctrl_decoder_bit_T_379 ;  
   wire _id_ctrl_decoder_bit_T_380 ;  
   wire _id_ctrl_decoder_bit_T_381 ;  
   wire _id_ctrl_decoder_bit_T_382 ;  
   wire _id_ctrl_decoder_bit_T_383 ;  
   wire _id_ctrl_decoder_bit_T_384 ;  
   wire _id_ctrl_decoder_bit_T_385 ;  
   wire _id_ctrl_decoder_bit_T_386 ;  
   wire _id_ctrl_decoder_bit_T_387 ;  
   wire _id_ctrl_decoder_bit_T_388 ;  
   wire _id_ctrl_decoder_bit_T_389 ;  
   wire _id_ctrl_decoder_bit_T_390 ;  
   wire _id_ctrl_decoder_bit_T_391 ;  
   wire _id_ctrl_decoder_bit_T_392 ;  
   wire _id_ctrl_decoder_bit_T_393 ;  
   wire _id_ctrl_decoder_bit_T_394 ;  
   wire _id_ctrl_decoder_bit_T_395 ;  
   wire _id_ctrl_decoder_bit_T_396 ;  
   wire _id_ctrl_decoder_bit_T_397 ;  
   wire _id_ctrl_decoder_bit_T_398 ;  
   wire _id_ctrl_decoder_bit_T_399 ;  
   wire _id_ctrl_decoder_bit_T_400 ;  
   wire _id_ctrl_decoder_bit_T_401 ;  
   wire _id_ctrl_decoder_bit_T_402 ;  
   wire _id_ctrl_decoder_bit_T_403 ;  
   wire _id_ctrl_decoder_bit_T_404 ;  
   wire _id_ctrl_decoder_bit_T_405 ;  
   wire _id_ctrl_decoder_bit_T_406 ;  
   wire _id_ctrl_decoder_bit_T_407 ;  
   wire _id_ctrl_decoder_bit_T_408 ;  
   wire _id_ctrl_decoder_bit_T_409 ;  
   wire _id_ctrl_decoder_bit_T_410 ;  
   wire _id_ctrl_decoder_bit_T_411 ;  
   wire _id_ctrl_decoder_bit_T_412 ;  
   wire _id_ctrl_decoder_bit_T_413 ;  
   wire _id_ctrl_decoder_bit_T_414 ;  
   wire _id_ctrl_decoder_bit_T_415 ;  
   wire _id_ctrl_decoder_bit_T_416 ;  
   wire _id_ctrl_decoder_bit_T_417 ;  
   wire _id_ctrl_decoder_bit_T_418 ;  
   wire _id_ctrl_decoder_bit_T_419 ;  
   wire _id_ctrl_decoder_bit_T_420 ;  
   wire _id_ctrl_decoder_bit_T_421 ;  
   wire _id_ctrl_decoder_bit_T_422 ;  
   wire _id_ctrl_decoder_bit_T_423 ;  
   wire _id_ctrl_decoder_bit_T_424 ;  
   wire _id_ctrl_decoder_bit_T_425 ;  
   wire _id_ctrl_decoder_bit_T_426 ;  
   wire _id_ctrl_decoder_bit_T_427 ;  
   wire _id_ctrl_decoder_bit_T_428 ;  
   wire _id_ctrl_decoder_bit_T_429 ;  
   wire _id_ctrl_decoder_bit_T_430 ;  
   wire _id_ctrl_decoder_bit_T_431 ;  
   wire _id_ctrl_decoder_bit_T_432 ;  
   wire _id_ctrl_decoder_bit_T_433 ;  
   wire _id_ctrl_decoder_bit_T_434 ;  
   wire _id_ctrl_decoder_bit_T_435 ;  
   wire _id_ctrl_decoder_bit_T_436 ;  
   wire _id_ctrl_decoder_bit_T_437 ;  
   wire _id_ctrl_decoder_bit_T_438 ;  
   wire _id_ctrl_decoder_bit_T_439 ;  
   wire _id_ctrl_decoder_bit_T_440 ;  
   wire _id_ctrl_decoder_bit_T_441 ;  
   wire _id_ctrl_decoder_bit_T_442 ;  
   wire _id_ctrl_decoder_bit_T_443 ;  
   wire _id_ctrl_decoder_bit_T_444 ;  
   wire _id_ctrl_decoder_bit_T_445 ;  
   wire _id_ctrl_decoder_bit_T_446 ;  
   wire _id_ctrl_decoder_bit_T_447 ;  
   wire _id_ctrl_decoder_bit_T_448 ;  
   wire _id_ctrl_decoder_bit_T_449 ;  
   wire _id_ctrl_decoder_bit_T_450 ;  
   wire _id_ctrl_decoder_bit_T_451 ;  
   wire _id_ctrl_decoder_bit_T_452 ;  
   wire _id_ctrl_decoder_bit_T_453 ;  
   wire _id_ctrl_decoder_bit_T_454 ;  
   wire _id_ctrl_decoder_bit_T_455 ;  
   wire _id_ctrl_decoder_bit_T_456 ;  
   wire _id_ctrl_decoder_bit_T_457 ;  
   wire _id_ctrl_decoder_bit_T_458 ;  
   wire _id_ctrl_decoder_bit_T_459 ;  
   wire _id_ctrl_decoder_bit_T_460 ;  
   wire _id_ctrl_decoder_bit_T_461 ;  
   wire _id_ctrl_decoder_bit_T_462 ;  
   wire _id_ctrl_decoder_bit_T_463 ;  
   wire _id_ctrl_decoder_bit_T_464 ;  
   wire _id_ctrl_decoder_bit_T_465 ;  
   wire _id_ctrl_decoder_bit_T_466 ;  
   wire _id_ctrl_decoder_bit_T_467 ;  
   wire _id_ctrl_decoder_bit_T_468 ;  
   wire _id_ctrl_decoder_bit_T_469 ;  
   wire _id_ctrl_decoder_bit_T_470 ;  
   wire _id_ctrl_decoder_bit_T_471 ;  
   wire _id_ctrl_decoder_bit_T_472 ;  
   wire _id_ctrl_decoder_bit_T_473 ;  
   wire _id_ctrl_decoder_bit_T_474 ;  
   wire _id_ctrl_decoder_bit_T_475 ;  
   wire _id_ctrl_decoder_bit_T_476 ;  
   wire _id_ctrl_decoder_bit_T_477 ;  
   wire id_ctrl_decoder_0 ;  
   wire [31:0] _id_ctrl_decoder_T ;  
   wire _id_ctrl_decoder_T_1 ;  
   wire [31:0] _id_ctrl_decoder_T_2 ;  
   wire _id_ctrl_decoder_T_3 ;  
   wire id_ctrl_decoder_1 ;  
   wire [31:0] _id_ctrl_decoder_T_5 ;  
   wire id_ctrl_decoder_3 ;  
   wire [31:0] _id_ctrl_decoder_T_7 ;  
   wire id_ctrl_decoder_4 ;  
   wire [31:0] _id_ctrl_decoder_T_9 ;  
   wire id_ctrl_decoder_5 ;  
   wire [31:0] _id_ctrl_decoder_T_11 ;  
   wire _id_ctrl_decoder_T_12 ;  
   wire [31:0] _id_ctrl_decoder_T_13 ;  
   wire _id_ctrl_decoder_T_14 ;  
   wire [31:0] _id_ctrl_decoder_T_15 ;  
   wire _id_ctrl_decoder_T_16 ;  
   wire [31:0] _id_ctrl_decoder_T_17 ;  
   wire _id_ctrl_decoder_T_18 ;  
   wire _id_ctrl_decoder_T_20 ;  
   wire _id_ctrl_decoder_T_21 ;  
   wire id_ctrl_decoder_6 ;  
   wire [31:0] _id_ctrl_decoder_T_22 ;  
   wire _id_ctrl_decoder_T_23 ;  
   wire [31:0] _id_ctrl_decoder_T_24 ;  
   wire _id_ctrl_decoder_T_25 ;  
   wire [31:0] _id_ctrl_decoder_T_26 ;  
   wire _id_ctrl_decoder_T_27 ;  
   wire [31:0] _id_ctrl_decoder_T_28 ;  
   wire _id_ctrl_decoder_T_29 ;  
   wire [31:0] _id_ctrl_decoder_T_30 ;  
   wire _id_ctrl_decoder_T_31 ;  
   wire _id_ctrl_decoder_T_33 ;  
   wire _id_ctrl_decoder_T_34 ;  
   wire _id_ctrl_decoder_T_35 ;  
   wire id_ctrl_decoder_7 ;  
   wire [31:0] _id_ctrl_decoder_T_36 ;  
   wire _id_ctrl_decoder_T_37 ;  
   wire [31:0] _id_ctrl_decoder_T_38 ;  
   wire _id_ctrl_decoder_T_39 ;  
   wire [31:0] _id_ctrl_decoder_T_40 ;  
   wire _id_ctrl_decoder_T_41 ;  
   wire [31:0] _id_ctrl_decoder_T_42 ;  
   wire _id_ctrl_decoder_T_43 ;  
   wire [31:0] _id_ctrl_decoder_T_44 ;  
   wire _id_ctrl_decoder_T_45 ;  
   wire _id_ctrl_decoder_T_47 ;  
   wire _id_ctrl_decoder_T_48 ;  
   wire _id_ctrl_decoder_T_49 ;  
   wire id_ctrl_decoder_lo ;  
   wire _id_ctrl_decoder_T_51 ;  
   wire [31:0] _id_ctrl_decoder_T_52 ;  
   wire _id_ctrl_decoder_T_53 ;  
   wire [31:0] _id_ctrl_decoder_T_54 ;  
   wire _id_ctrl_decoder_T_55 ;  
   wire _id_ctrl_decoder_T_57 ;  
   wire _id_ctrl_decoder_T_58 ;  
   wire id_ctrl_decoder_hi ;  
   wire [1:0] id_ctrl_decoder_9 ;  
   wire [31:0] _id_ctrl_decoder_T_59 ;  
   wire _id_ctrl_decoder_T_60 ;  
   wire [31:0] _id_ctrl_decoder_T_61 ;  
   wire _id_ctrl_decoder_T_62 ;  
   wire [31:0] _id_ctrl_decoder_T_63 ;  
   wire _id_ctrl_decoder_T_64 ;  
   wire _id_ctrl_decoder_T_66 ;  
   wire _id_ctrl_decoder_T_67 ;  
   wire _id_ctrl_decoder_T_68 ;  
   wire id_ctrl_decoder_lo_1 ;  
   wire _id_ctrl_decoder_T_70 ;  
   wire id_ctrl_decoder_hi_1 ;  
   wire [1:0] id_ctrl_decoder_10 ;  
   wire _id_ctrl_decoder_T_73 ;  
   wire _id_ctrl_decoder_T_75 ;  
   wire id_ctrl_decoder_lo_2 ;  
   wire [31:0] _id_ctrl_decoder_T_77 ;  
   wire _id_ctrl_decoder_T_78 ;  
   wire id_ctrl_decoder_hi_lo ;  
   wire [31:0] _id_ctrl_decoder_T_80 ;  
   wire _id_ctrl_decoder_T_81 ;  
   wire [31:0] _id_ctrl_decoder_T_82 ;  
   wire _id_ctrl_decoder_T_83 ;  
   wire _id_ctrl_decoder_T_85 ;  
   wire _id_ctrl_decoder_T_87 ;  
   wire id_ctrl_decoder_hi_hi ;  
   wire [2:0] id_ctrl_decoder_11 ;  
   wire [31:0] _id_ctrl_decoder_T_88 ;  
   wire _id_ctrl_decoder_T_89 ;  
   wire [31:0] _id_ctrl_decoder_T_90 ;  
   wire _id_ctrl_decoder_T_91 ;  
   wire id_ctrl_decoder_12 ;  
   wire [31:0] _id_ctrl_decoder_T_93 ;  
   wire _id_ctrl_decoder_T_94 ;  
   wire [31:0] _id_ctrl_decoder_T_95 ;  
   wire _id_ctrl_decoder_T_96 ;  
   wire [31:0] _id_ctrl_decoder_T_97 ;  
   wire _id_ctrl_decoder_T_98 ;  
   wire [31:0] _id_ctrl_decoder_T_99 ;  
   wire _id_ctrl_decoder_T_100 ;  
   wire _id_ctrl_decoder_T_102 ;  
   wire _id_ctrl_decoder_T_103 ;  
   wire id_ctrl_decoder_lo_lo ;  
   wire [31:0] _id_ctrl_decoder_T_104 ;  
   wire _id_ctrl_decoder_T_105 ;  
   wire [31:0] _id_ctrl_decoder_T_106 ;  
   wire _id_ctrl_decoder_T_107 ;  
   wire _id_ctrl_decoder_T_109 ;  
   wire [31:0] _id_ctrl_decoder_T_110 ;  
   wire _id_ctrl_decoder_T_111 ;  
   wire [31:0] _id_ctrl_decoder_T_112 ;  
   wire _id_ctrl_decoder_T_113 ;  
   wire [31:0] _id_ctrl_decoder_T_114 ;  
   wire _id_ctrl_decoder_T_115 ;  
   wire [31:0] _id_ctrl_decoder_T_116 ;  
   wire _id_ctrl_decoder_T_117 ;  
   wire _id_ctrl_decoder_T_119 ;  
   wire _id_ctrl_decoder_T_120 ;  
   wire _id_ctrl_decoder_T_121 ;  
   wire _id_ctrl_decoder_T_122 ;  
   wire _id_ctrl_decoder_T_123 ;  
   wire id_ctrl_decoder_lo_hi ;  
   wire [31:0] _id_ctrl_decoder_T_124 ;  
   wire _id_ctrl_decoder_T_125 ;  
   wire [31:0] _id_ctrl_decoder_T_126 ;  
   wire _id_ctrl_decoder_T_127 ;  
   wire [31:0] _id_ctrl_decoder_T_128 ;  
   wire _id_ctrl_decoder_T_129 ;  
   wire [31:0] _id_ctrl_decoder_T_130 ;  
   wire _id_ctrl_decoder_T_131 ;  
   wire [31:0] _id_ctrl_decoder_T_132 ;  
   wire _id_ctrl_decoder_T_133 ;  
   wire _id_ctrl_decoder_T_135 ;  
   wire _id_ctrl_decoder_T_136 ;  
   wire _id_ctrl_decoder_T_137 ;  
   wire id_ctrl_decoder_hi_lo_1 ;  
   wire [31:0] _id_ctrl_decoder_T_138 ;  
   wire _id_ctrl_decoder_T_139 ;  
   wire [31:0] _id_ctrl_decoder_T_140 ;  
   wire _id_ctrl_decoder_T_141 ;  
   wire [31:0] _id_ctrl_decoder_T_142 ;  
   wire _id_ctrl_decoder_T_143 ;  
   wire _id_ctrl_decoder_T_145 ;  
   wire _id_ctrl_decoder_T_146 ;  
   wire _id_ctrl_decoder_T_147 ;  
   wire id_ctrl_decoder_hi_hi_1 ;  
   wire [3:0] id_ctrl_decoder_13 ;  
   wire _id_ctrl_decoder_bit_T_479 ;  
   wire _id_ctrl_decoder_bit_T_480 ;  
   wire _id_ctrl_decoder_bit_T_481 ;  
   wire _id_ctrl_decoder_bit_T_482 ;  
   wire _id_ctrl_decoder_bit_T_483 ;  
   wire _id_ctrl_decoder_bit_T_484 ;  
   wire _id_ctrl_decoder_bit_T_485 ;  
   wire _id_ctrl_decoder_bit_T_486 ;  
   wire _id_ctrl_decoder_bit_T_487 ;  
   wire _id_ctrl_decoder_bit_T_488 ;  
   wire _id_ctrl_decoder_bit_T_489 ;  
   wire _id_ctrl_decoder_bit_T_490 ;  
   wire _id_ctrl_decoder_bit_T_491 ;  
   wire _id_ctrl_decoder_bit_T_492 ;  
   wire _id_ctrl_decoder_bit_T_493 ;  
   wire _id_ctrl_decoder_bit_T_494 ;  
   wire _id_ctrl_decoder_bit_T_495 ;  
   wire _id_ctrl_decoder_bit_T_496 ;  
   wire _id_ctrl_decoder_bit_T_497 ;  
   wire _id_ctrl_decoder_bit_T_498 ;  
   wire _id_ctrl_decoder_bit_T_499 ;  
   wire _id_ctrl_decoder_bit_T_500 ;  
   wire _id_ctrl_decoder_bit_T_501 ;  
   wire _id_ctrl_decoder_bit_T_502 ;  
   wire _id_ctrl_decoder_bit_T_503 ;  
   wire _id_ctrl_decoder_bit_T_504 ;  
   wire _id_ctrl_decoder_bit_T_505 ;  
   wire _id_ctrl_decoder_bit_T_506 ;  
   wire _id_ctrl_decoder_bit_T_507 ;  
   wire _id_ctrl_decoder_bit_T_508 ;  
   wire _id_ctrl_decoder_bit_T_509 ;  
   wire _id_ctrl_decoder_bit_T_510 ;  
   wire _id_ctrl_decoder_bit_T_511 ;  
   wire _id_ctrl_decoder_bit_T_512 ;  
   wire _id_ctrl_decoder_bit_T_513 ;  
   wire _id_ctrl_decoder_bit_T_514 ;  
   wire id_ctrl_decoder_14 ;  
   wire _id_ctrl_decoder_T_149 ;  
   wire [31:0] _id_ctrl_decoder_T_150 ;  
   wire _id_ctrl_decoder_T_151 ;  
   wire [31:0] _id_ctrl_decoder_T_152 ;  
   wire _id_ctrl_decoder_T_153 ;  
   wire _id_ctrl_decoder_T_155 ;  
   wire id_ctrl_decoder_lo_lo_1 ;  
   wire [31:0] _id_ctrl_decoder_T_156 ;  
   wire _id_ctrl_decoder_T_157 ;  
   wire [31:0] _id_ctrl_decoder_T_158 ;  
   wire _id_ctrl_decoder_T_159 ;  
   wire id_ctrl_decoder_lo_hi_1 ;  
   wire [31:0] _id_ctrl_decoder_T_161 ;  
   wire id_ctrl_decoder_hi_hi_hi ;  
   wire [31:0] _id_ctrl_decoder_T_163 ;  
   wire _id_ctrl_decoder_T_164 ;  
   wire [31:0] _id_ctrl_decoder_T_165 ;  
   wire _id_ctrl_decoder_T_166 ;  
   wire _id_ctrl_decoder_T_168 ;  
   wire _id_ctrl_decoder_T_169 ;  
   wire id_ctrl_decoder_hi_lo_2 ;  
   wire [31:0] _id_ctrl_decoder_T_170 ;  
   wire id_ctrl_decoder_hi_hi_lo ;  
   wire [4:0] id_ctrl_decoder_15 ;  
   wire [31:0] _id_ctrl_decoder_T_172 ;  
   wire _id_ctrl_decoder_T_173 ;  
   wire [31:0] _id_ctrl_decoder_T_174 ;  
   wire [31:0] _id_ctrl_decoder_T_176 ;  
   wire id_ctrl_decoder_18 ;  
   wire [31:0] _id_ctrl_decoder_T_189 ;  
   wire _id_ctrl_decoder_T_190 ;  
   wire _id_ctrl_decoder_T_192 ;  
   wire _id_ctrl_decoder_T_194 ;  
   wire _id_ctrl_decoder_T_195 ;  
   wire id_ctrl_decoder_19 ;  
   wire [31:0] _id_ctrl_decoder_T_196 ;  
   wire id_ctrl_decoder_21 ;  
   wire _id_ctrl_decoder_T_199 ;  
   wire _id_ctrl_decoder_T_201 ;  
   wire [31:0] _id_ctrl_decoder_T_202 ;  
   wire _id_ctrl_decoder_T_203 ;  
   wire [31:0] _id_ctrl_decoder_T_204 ;  
   wire _id_ctrl_decoder_T_205 ;  
   wire [31:0] _id_ctrl_decoder_T_206 ;  
   wire _id_ctrl_decoder_T_207 ;  
   wire [31:0] _id_ctrl_decoder_T_208 ;  
   wire _id_ctrl_decoder_T_209 ;  
   wire [31:0] _id_ctrl_decoder_T_210 ;  
   wire _id_ctrl_decoder_T_211 ;  
   wire _id_ctrl_decoder_T_213 ;  
   wire _id_ctrl_decoder_T_214 ;  
   wire _id_ctrl_decoder_T_215 ;  
   wire _id_ctrl_decoder_T_216 ;  
   wire _id_ctrl_decoder_T_217 ;  
   wire id_ctrl_decoder_22 ;  
   wire [31:0] _id_ctrl_decoder_T_218 ;  
   wire id_ctrl_decoder_lo_5 ;  
   wire [31:0] _id_ctrl_decoder_T_220 ;  
   wire id_ctrl_decoder_hi_lo_3 ;  
   wire [31:0] _id_ctrl_decoder_T_222 ;  
   wire _id_ctrl_decoder_T_223 ;  
   wire [31:0] _id_ctrl_decoder_T_224 ;  
   wire _id_ctrl_decoder_T_225 ;  
   wire [31:0] _id_ctrl_decoder_T_226 ;  
   wire _id_ctrl_decoder_T_227 ;  
   wire _id_ctrl_decoder_T_229 ;  
   wire _id_ctrl_decoder_T_230 ;  
   wire _id_ctrl_decoder_T_231 ;  
   wire id_ctrl_decoder_hi_hi_3 ;  
   wire [2:0] id_ctrl_decoder_23 ;  
   wire [31:0] _id_ctrl_decoder_T_232 ;  
   wire id_ctrl_decoder_24 ;  
   wire id_ctrl_decoder_25 ;  
   wire [31:0] _id_ctrl_decoder_T_236 ;  
   wire id_ctrl_decoder_26 ;  
   wire [31:0] _id_ctrl_decoder_T_238 ;  
   wire _id_ctrl_decoder_T_239 ;  
   wire [31:0] _id_ctrl_decoder_T_240 ;  
   wire _id_ctrl_decoder_T_241 ;  
   wire [31:0] _id_ctrl_decoder_T_242 ;  
   wire _id_ctrl_decoder_T_243 ;  
   wire _id_ctrl_decoder_T_245 ;  
   wire id_ctrl_decoder_27 ;  
   wire [4:0] id_raddr3 ;  
   wire [4:0] id_raddr2 ;  
   wire [4:0] id_raddr1 ;  
   wire [4:0] id_waddr ;  
   reg id_reg_fence ;  
   reg [31:0] _RAND_83 ;  
   wire [63:0] _id_rs_T_4 ;  
   wire [63:0] _id_rs_T_9 ;  
   wire _id_csr_en_T ;  
   wire _id_csr_en_T_1 ;  
   wire _id_csr_en_T_2 ;  
   wire _id_csr_en_T_3 ;  
   wire id_csr_en ;  
   wire id_system_insn ;  
   wire _id_csr_ren_T_3 ;  
   wire id_csr_ren ;  
   wire _id_sfence_T ;  
   wire id_sfence ;  
   wire _id_csr_flush_T ;  
   wire _id_csr_flush_T_2 ;  
   wire _id_csr_flush_T_3 ;  
   wire id_csr_flush ;  
   wire _id_illegal_insn_T_4 ;  
   wire _id_illegal_insn_T_5 ;  
   wire _id_illegal_insn_T_8 ;  
   wire _id_illegal_insn_T_9 ;  
   wire _id_illegal_insn_T_10 ;  
   wire _id_illegal_insn_T_11 ;  
   wire _id_illegal_insn_T_12 ;  
   wire _id_illegal_insn_T_15 ;  
   wire _id_illegal_insn_T_16 ;  
   wire _id_illegal_insn_T_19 ;  
   wire _id_illegal_insn_T_20 ;  
   wire _id_illegal_insn_T_40 ;  
   wire _id_illegal_insn_T_41 ;  
   wire _id_illegal_insn_T_42 ;  
   wire _id_illegal_insn_T_43 ;  
   wire _id_illegal_insn_T_46 ;  
   wire _id_illegal_insn_T_47 ;  
   wire id_illegal_insn ;  
   wire id_amo_aq ;  
   wire id_amo_rl ;  
   wire [3:0] id_fence_succ ;  
   wire _id_fence_next_T ;  
   wire id_fence_next ;  
   wire id_mem_busy ;  
   wire _GEN_0 ;  
   wire _id_do_fence_x8_T_1 ;  
   wire _id_do_fence_x8_T_2 ;  
   wire _id_do_fence_x8_T_4 ;  
   wire _id_do_fence_x8_T_5 ;  
   wire id_do_fence_x8 ;  
   wire _T_1 ;  
   wire _T_2 ;  
   wire _T_3 ;  
   wire _T_4 ;  
   wire _T_5 ;  
   wire _T_6 ;  
   wire id_xcpt ;  
   wire [1:0] _T_7 ;  
   wire [3:0] _T_8 ;  
   wire [3:0] _T_9 ;  
   wire [3:0] _T_10 ;  
   wire [3:0] _T_11 ;  
   wire [3:0] _T_12 ;  
   wire [4:0] ex_waddr ;  
   wire [4:0] mem_waddr ;  
   wire [4:0] wb_waddr ;  
   wire _T_23 ;  
   wire _T_24 ;  
   wire _T_26 ;  
   wire id_bypass_src_0_0 ;  
   wire _id_bypass_src_T_1 ;  
   wire id_bypass_src_0_1 ;  
   wire _id_bypass_src_T_2 ;  
   wire id_bypass_src_0_2 ;  
   wire id_bypass_src_0_3 ;  
   wire id_bypass_src_1_0 ;  
   wire _id_bypass_src_T_5 ;  
   wire id_bypass_src_1_1 ;  
   wire _id_bypass_src_T_6 ;  
   wire id_bypass_src_1_2 ;  
   wire id_bypass_src_1_3 ;  
   reg ex_reg_rs_bypass_0 ;  
   reg [31:0] _RAND_84 ;  
   reg ex_reg_rs_bypass_1 ;  
   reg [31:0] _RAND_85 ;  
   reg [1:0] ex_reg_rs_lsb_0 ;  
   reg [31:0] _RAND_86 ;  
   reg [1:0] ex_reg_rs_lsb_1 ;  
   reg [31:0] _RAND_87 ;  
   reg [61:0] ex_reg_rs_msb_0 ;  
   reg [63:0] _RAND_88 ;  
   reg [61:0] ex_reg_rs_msb_1 ;  
   reg [63:0] _RAND_89 ;  
   wire _ex_rs_T ;  
   wire [63:0] _ex_rs_T_1 ;  
   wire _ex_rs_T_2 ;  
   wire [63:0] _ex_rs_T_3 ;  
   wire _ex_rs_T_4 ;  
   wire [63:0] _ex_rs_T_5 ;  
   wire [63:0] _ex_rs_T_6 ;  
   wire _ex_rs_T_7 ;  
   wire [63:0] _ex_rs_T_8 ;  
   wire _ex_rs_T_9 ;  
   wire [63:0] _ex_rs_T_10 ;  
   wire _ex_rs_T_11 ;  
   wire [63:0] _ex_rs_T_12 ;  
   wire [63:0] _ex_rs_T_13 ;  
   wire [63:0] ex_rs_1 ;  
   wire _ex_imm_sign_T ;  
   wire _ex_imm_sign_T_2 ;  
   wire ex_imm_sign ;  
   wire _ex_imm_b30_20_T ;  
   wire [10:0] _ex_imm_b30_20_T_2 ;  
   wire _ex_imm_b19_12_T ;  
   wire _ex_imm_b19_12_T_1 ;  
   wire _ex_imm_b19_12_T_2 ;  
   wire [7:0] _ex_imm_b19_12_T_4 ;  
   wire _ex_imm_b11_T_2 ;  
   wire _ex_imm_b11_T_3 ;  
   wire _ex_imm_b11_T_5 ;  
   wire _ex_imm_b11_T_6 ;  
   wire _ex_imm_b11_T_8 ;  
   wire _ex_imm_b11_T_9 ;  
   wire _ex_imm_b11_T_10 ;  
   wire [5:0] ex_imm_lo_hi_hi ;  
   wire _ex_imm_b4_1_T_1 ;  
   wire _ex_imm_b4_1_T_3 ;  
   wire [3:0] _ex_imm_b4_1_T_8 ;  
   wire [3:0] _ex_imm_b4_1_T_9 ;  
   wire [3:0] ex_imm_lo_hi_lo ;  
   wire _ex_imm_b0_T_2 ;  
   wire _ex_imm_b0_T_6 ;  
   wire _ex_imm_b0_T_7 ;  
   wire ex_imm_lo_lo ;  
   wire ex_imm_hi_lo_lo ;  
   wire [7:0] ex_imm_hi_lo_hi ;  
   wire [10:0] ex_imm_hi_hi_lo ;  
   wire ex_imm_hi_hi_hi ;  
   wire [31:0] ex_imm ;  
   wire [63:0] _ex_op1_T ;  
   wire _ex_op1_T_2 ;  
   wire [63:0] _ex_op1_T_3 ;  
   wire _ex_op1_T_4 ;  
   wire [63:0] _ex_op2_T ;  
   wire [3:0] _ex_op2_T_1 ;  
   wire _ex_op2_T_2 ;  
   wire [63:0] _ex_op2_T_3 ;  
   wire _ex_op2_T_4 ;  
   wire [63:0] _ex_op2_T_5 ;  
   wire _ex_op2_T_6 ;  
   wire _ctrl_killd_T_1 ;  
   wire _ctrl_killd_T_2 ;  
   wire _T_123 ;  
   wire _T_124 ;  
   wire _data_hazard_ex_T ;  
   wire _data_hazard_ex_T_1 ;  
   wire _T_125 ;  
   wire _T_126 ;  
   wire _data_hazard_ex_T_2 ;  
   wire _data_hazard_ex_T_3 ;  
   wire _data_hazard_ex_T_6 ;  
   wire _T_127 ;  
   wire _T_128 ;  
   wire _data_hazard_ex_T_4 ;  
   wire _data_hazard_ex_T_5 ;  
   wire _data_hazard_ex_T_7 ;  
   wire data_hazard_ex ;  
   wire _ex_cannot_bypass_T ;  
   wire _ex_cannot_bypass_T_1 ;  
   wire _ex_cannot_bypass_T_2 ;  
   wire _ex_cannot_bypass_T_4 ;  
   wire ex_cannot_bypass ;  
   wire _id_ex_hazard_T ;  
   wire _fp_data_hazard_ex_T_1 ;  
   wire _fp_data_hazard_ex_T_3 ;  
   wire _fp_data_hazard_ex_T_8 ;  
   wire _fp_data_hazard_ex_T_4 ;  
   wire _fp_data_hazard_ex_T_5 ;  
   wire _fp_data_hazard_ex_T_9 ;  
   wire _fp_data_hazard_ex_T_7 ;  
   wire _fp_data_hazard_ex_T_10 ;  
   wire fp_data_hazard_ex ;  
   wire _id_ex_hazard_T_1 ;  
   wire id_ex_hazard ;  
   wire _data_hazard_mem_T ;  
   wire _data_hazard_mem_T_1 ;  
   wire _data_hazard_mem_T_2 ;  
   wire _data_hazard_mem_T_3 ;  
   wire _data_hazard_mem_T_6 ;  
   wire _data_hazard_mem_T_4 ;  
   wire _data_hazard_mem_T_5 ;  
   wire _data_hazard_mem_T_7 ;  
   wire data_hazard_mem ;  
   wire _mem_cannot_bypass_T ;  
   wire _mem_cannot_bypass_T_1 ;  
   wire _mem_cannot_bypass_T_2 ;  
   wire _mem_cannot_bypass_T_4 ;  
   wire mem_cannot_bypass ;  
   wire _id_mem_hazard_T ;  
   wire _fp_data_hazard_mem_T_1 ;  
   wire _fp_data_hazard_mem_T_3 ;  
   wire _fp_data_hazard_mem_T_8 ;  
   wire _fp_data_hazard_mem_T_4 ;  
   wire _fp_data_hazard_mem_T_5 ;  
   wire _fp_data_hazard_mem_T_9 ;  
   wire _fp_data_hazard_mem_T_7 ;  
   wire _fp_data_hazard_mem_T_10 ;  
   wire fp_data_hazard_mem ;  
   wire _id_mem_hazard_T_1 ;  
   wire id_mem_hazard ;  
   wire _ctrl_stalld_T ;  
   wire _data_hazard_wb_T ;  
   wire _data_hazard_wb_T_1 ;  
   wire _data_hazard_wb_T_2 ;  
   wire _data_hazard_wb_T_3 ;  
   wire _data_hazard_wb_T_6 ;  
   wire _data_hazard_wb_T_4 ;  
   wire _data_hazard_wb_T_5 ;  
   wire _data_hazard_wb_T_7 ;  
   wire data_hazard_wb ;  
   wire wb_dcache_miss ;  
   wire wb_set_sboard ;  
   wire _id_wb_hazard_T ;  
   wire _fp_data_hazard_wb_T_1 ;  
   wire _fp_data_hazard_wb_T_3 ;  
   wire _fp_data_hazard_wb_T_8 ;  
   wire _fp_data_hazard_wb_T_4 ;  
   wire _fp_data_hazard_wb_T_5 ;  
   wire _fp_data_hazard_wb_T_9 ;  
   wire _fp_data_hazard_wb_T_7 ;  
   wire _fp_data_hazard_wb_T_10 ;  
   wire fp_data_hazard_wb ;  
   wire _id_wb_hazard_T_1 ;  
   wire id_wb_hazard ;  
   wire _ctrl_stalld_T_1 ;  
   reg [31:0] _r ;  
   reg [31:0] _RAND_90 ;  
   wire [31:0] r ;  
   wire [31:0] _id_sboard_hazard_T ;  
   wire dmem_resp_valid ;  
   wire dmem_resp_replay ;  
   wire dmem_resp_xpu ;  
   wire _T_117 ;  
   wire ll_wen_x1 ;  
   wire ll_wen ;  
   wire [4:0] dmem_resp_waddr ;  
   wire [4:0] ll_waddr ;  
   wire _id_sboard_hazard_T_2 ;  
   wire _id_sboard_hazard_T_3 ;  
   wire _id_sboard_hazard_T_5 ;  
   wire _id_sboard_hazard_T_6 ;  
   wire [31:0] _id_sboard_hazard_T_7 ;  
   wire _id_sboard_hazard_T_9 ;  
   wire _id_sboard_hazard_T_10 ;  
   wire _id_sboard_hazard_T_12 ;  
   wire _id_sboard_hazard_T_13 ;  
   wire _id_sboard_hazard_T_21 ;  
   wire [31:0] _id_sboard_hazard_T_14 ;  
   wire _id_sboard_hazard_T_16 ;  
   wire _id_sboard_hazard_T_17 ;  
   wire _id_sboard_hazard_T_19 ;  
   wire _id_sboard_hazard_T_20 ;  
   wire id_sboard_hazard ;  
   wire _ctrl_stalld_T_2 ;  
   wire _ctrl_stalld_T_3 ;  
   wire _ctrl_stalld_T_4 ;  
   wire _ctrl_stalld_T_5 ;  
   wire _ctrl_stalld_T_6 ;  
   wire _ctrl_stalld_T_7 ;  
   wire _ctrl_stalld_T_9 ;  
   wire _ctrl_stalld_T_10 ;  
   reg [31:0] id_stall_fpu__r ;  
   reg [31:0] _RAND_91 ;  
   wire [31:0] _id_stall_fpu_T_18 ;  
   wire _id_stall_fpu_T_20 ;  
   wire [31:0] _id_stall_fpu_T_21 ;  
   wire _id_stall_fpu_T_23 ;  
   wire _id_stall_fpu_T_30 ;  
   wire [31:0] _id_stall_fpu_T_24 ;  
   wire _id_stall_fpu_T_26 ;  
   wire _id_stall_fpu_T_31 ;  
   wire [31:0] _id_stall_fpu_T_27 ;  
   wire _id_stall_fpu_T_29 ;  
   wire id_stall_fpu ;  
   wire _ctrl_stalld_T_11 ;  
   wire _ctrl_stalld_T_12 ;  
   reg blocked ;  
   reg [31:0] _RAND_92 ;  
   wire dcache_blocked ;  
   wire _ctrl_stalld_T_13 ;  
   wire _ctrl_stalld_T_14 ;  
   wire wb_wxd ;  
   wire _ctrl_stalld_T_18 ;  
   wire _ctrl_stalld_T_19 ;  
   wire _ctrl_stalld_T_21 ;  
   wire _ctrl_stalld_T_22 ;  
   wire _ctrl_stalld_T_23 ;  
   wire _ctrl_stalld_T_26 ;  
   wire _ctrl_stalld_T_27 ;  
   wire ctrl_stalld ;  
   wire _ctrl_killd_T_3 ;  
   wire ctrl_killd ;  
   wire _ex_reg_replay_T_1 ;  
   wire _T_29 ;  
   wire _T_30 ;  
   wire _GEN_1 ;  
   wire _GEN_2 ;  
   wire [1:0] _T_31 ;  
   wire _T_32 ;  
   wire _GEN_5 ;  
   wire [1:0] _T_33 ;  
   wire _T_34 ;  
   wire _T_35 ;  
   wire _GEN_9 ;  
   wire _ex_reg_flush_pipe_T ;  
   wire _T_37 ;  
   wire _T_38 ;  
   wire [1:0] _ex_reg_mem_size_T_1 ;  
   wire _do_bypass_T ;  
   wire _do_bypass_T_1 ;  
   wire do_bypass ;  
   wire _T_40 ;  
   wire _wb_valid_T_1 ;  
   wire wb_valid ;  
   wire wb_wen ;  
   wire rf_wen ;  
   wire [4:0] rf_waddr ;  
   wire _T_118 ;  
   wire _T_121 ;  
   wire _rf_wdata_T ;  
   wire [63:0] ll_wdata ;  
   wire _rf_wdata_T_2 ;  
   wire [63:0] _rf_wdata_T_4 ;  
   wire [63:0] _rf_wdata_T_5 ;  
   wire [63:0] rf_wdata ;  
   wire [63:0] _GEN_226 ;  
   wire [63:0] _GEN_233 ;  
   wire [63:0] id_rs_0 ;  
   wire _do_bypass_T_2 ;  
   wire _do_bypass_T_3 ;  
   wire do_bypass_1 ;  
   wire _T_42 ;  
   wire _T_122 ;  
   wire [63:0] _GEN_227 ;  
   wire [63:0] _GEN_234 ;  
   wire [63:0] id_rs_1 ;  
   wire [31:0] inst ;  
   wire _id_load_use_T ;  
   wire id_load_use ;  
   wire _T_44 ;  
   wire _T_45 ;  
   wire _replay_ex_structural_T_1 ;  
   wire _replay_ex_structural_T_3 ;  
   wire replay_ex_structural ;  
   wire replay_ex_load_use ;  
   wire _replay_ex_T ;  
   wire _replay_ex_T_1 ;  
   wire replay_ex ;  
   wire _ctrl_killx_T ;  
   wire ctrl_killx ;  
   wire _ex_slow_bypass_T ;  
   wire _ex_slow_bypass_T_1 ;  
   wire ex_slow_bypass ;  
   wire _ex_sfence_T_1 ;  
   wire ex_sfence ;  
   wire ex_xcpt ;  
   wire _mem_pc_valid_T ;  
   wire mem_pc_valid ;  
   wire _mem_npc_misaligned_T_3 ;  
   wire mem_npc_misaligned ;  
   wire _mem_int_wdata_T_1 ;  
   wire _mem_int_wdata_T_2 ;  
   wire [63:0] mem_int_wdata ;  
   wire _mem_cfi_T ;  
   wire mem_cfi ;  
   wire _mem_cfi_taken_T_1 ;  
   wire mem_cfi_taken ;  
   wire _T_56 ;  
   wire _mem_reg_load_T ;  
   wire _mem_reg_load_T_1 ;  
   wire _mem_reg_load_T_2 ;  
   wire _mem_reg_load_T_4 ;  
   wire _mem_reg_load_T_5 ;  
   wire _mem_reg_load_T_6 ;  
   wire _mem_reg_load_T_7 ;  
   wire _mem_reg_load_T_8 ;  
   wire _mem_reg_load_T_9 ;  
   wire _mem_reg_load_T_10 ;  
   wire _mem_reg_load_T_11 ;  
   wire _mem_reg_load_T_12 ;  
   wire _mem_reg_load_T_13 ;  
   wire _mem_reg_load_T_14 ;  
   wire _mem_reg_load_T_15 ;  
   wire _mem_reg_load_T_16 ;  
   wire _mem_reg_load_T_17 ;  
   wire _mem_reg_load_T_18 ;  
   wire _mem_reg_load_T_19 ;  
   wire _mem_reg_load_T_20 ;  
   wire _mem_reg_load_T_21 ;  
   wire _mem_reg_load_T_22 ;  
   wire _mem_reg_load_T_23 ;  
   wire _mem_reg_store_T ;  
   wire _mem_reg_store_T_1 ;  
   wire _mem_reg_store_T_2 ;  
   wire _mem_reg_store_T_4 ;  
   wire _mem_reg_store_T_22 ;  
   wire _mem_reg_store_T_23 ;  
   wire [63:0] _mem_reg_wdata_T ;  
   wire _T_58 ;  
   wire _T_59 ;  
   wire _mem_reg_rs2_T ;  
   wire [7:0] mem_reg_rs2_hi ;  
   wire [63:0] _mem_reg_rs2_T_1 ;  
   wire _mem_reg_rs2_T_2 ;  
   wire [15:0] mem_reg_rs2_hi_3 ;  
   wire [63:0] _mem_reg_rs2_T_3 ;  
   wire _mem_reg_rs2_T_4 ;  
   wire [31:0] mem_reg_rs2_hi_5 ;  
   wire [63:0] _mem_reg_rs2_T_5 ;  
   wire _T_60 ;  
   wire _GEN_77 ;  
   wire _GEN_78 ;  
   wire _mem_breakpoint_T ;  
   wire _mem_breakpoint_T_1 ;  
   wire mem_breakpoint ;  
   wire _mem_debug_breakpoint_T ;  
   wire _mem_debug_breakpoint_T_1 ;  
   wire mem_debug_breakpoint ;  
   wire mem_ldst_xcpt ;  
   wire [3:0] mem_ldst_cause ;  
   wire _T_61 ;  
   wire _T_62 ;  
   wire _T_63 ;  
   wire _T_64 ;  
   wire mem_xcpt ;  
   wire [3:0] _T_65 ;  
   wire dcache_kill_mem ;  
   wire _fpu_kill_mem_T ;  
   wire fpu_kill_mem ;  
   wire _replay_mem_T ;  
   wire replay_mem ;  
   wire _killm_common_T ;  
   wire _killm_common_T_1 ;  
   wire killm_common ;  
   reg div_io_kill_REG ;  
   reg [31:0] _RAND_93 ;  
   wire _ctrl_killm_T ;  
   wire ctrl_killm ;  
   wire _wb_reg_wdata_T_1 ;  
   wire _wb_reg_wdata_T_2 ;  
   wire [2:0] _T_100 ;  
   wire [3:0] _T_101 ;  
   wire [3:0] _T_102 ;  
   wire [3:0] _T_103 ;  
   wire [3:0] _T_104 ;  
   wire [63:0] wb_cause ;  
   wire _T_105 ;  
   wire _T_107 ;  
   wire _T_109 ;  
   wire _T_111 ;  
   wire _T_113 ;  
   wire _T_115 ;  
   wire _csr_io_inst_0_T_1 ;  
   wire [15:0] csr_io_inst_0_hi ;  
   wire [15:0] csr_io_inst_0_lo ;  
   wire _tval_valid_T ;  
   wire _tval_valid_T_1 ;  
   wire _tval_valid_T_6 ;  
   wire _tval_valid_T_9 ;  
   wire _tval_valid_T_10 ;  
   wire _tval_valid_T_11 ;  
   wire _tval_valid_T_12 ;  
   wire _tval_valid_T_13 ;  
   wire _tval_valid_T_14 ;  
   wire _tval_valid_T_15 ;  
   wire _tval_valid_T_16 ;  
   wire _tval_valid_T_17 ;  
   wire _tval_valid_T_18 ;  
   wire tval_valid ;  
   wire [24:0] a_1 ;  
   wire _csr_io_tval_msb_T ;  
   wire _csr_io_tval_msb_T_1 ;  
   wire _csr_io_tval_msb_T_2 ;  
   wire msb_1 ;  
   wire [38:0] csr_io_tval_lo ;  
   wire [39:0] _csr_io_tval_T ;  
   wire [2:0] _csr_io_rw_cmd_T ;  
   wire [31:0] _T_129 ;  
   wire [31:0] _T_130 ;  
   wire [31:0] _T_132 ;  
   wire _T_134 ;  
   wire [31:0] _T_135 ;  
   wire [31:0] _T_136 ;  
   wire [31:0] _T_137 ;  
   wire _T_138 ;  
   wire _id_stall_fpu_T ;  
   wire _id_stall_fpu_T_1 ;  
   wire _id_stall_fpu_T_2 ;  
   wire [31:0] _id_stall_fpu_T_4 ;  
   wire [31:0] _id_stall_fpu_T_5 ;  
   wire _id_stall_fpu_T_7 ;  
   wire [31:0] _id_stall_fpu_T_8 ;  
   wire [31:0] _id_stall_fpu_T_9 ;  
   wire [31:0] _id_stall_fpu_T_11 ;  
   wire _id_stall_fpu_T_12 ;  
   wire [31:0] _id_stall_fpu_T_13 ;  
   wire [31:0] _id_stall_fpu_T_14 ;  
   wire [31:0] _id_stall_fpu_T_16 ;  
   wire _id_stall_fpu_T_17 ;  
   wire _dcache_blocked_blocked_T_3 ;  
   wire _dcache_blocked_blocked_T_4 ;  
   wire _dcache_blocked_blocked_T_5 ;  
   wire _io_imem_req_bits_pc_T ;  
   wire [39:0] _io_imem_req_bits_pc_T_1 ;  
   wire _io_imem_flush_icache_T ;  
   wire _io_imem_might_request_imem_might_request_reg_T ;  
   wire _io_imem_btb_update_valid_T_1 ;  
   wire _io_imem_btb_update_valid_T_2 ;  
   wire _io_imem_btb_update_valid_T_4 ;  
   wire _io_imem_btb_update_bits_cfiType_T ;  
   wire _io_imem_btb_update_bits_cfiType_T_2 ;  
   wire [4:0] _io_imem_btb_update_bits_cfiType_T_5 ;  
   wire _io_imem_btb_update_bits_cfiType_T_6 ;  
   wire _io_imem_btb_update_bits_cfiType_T_7 ;  
   wire [1:0] _io_imem_btb_update_bits_cfiType_T_10 ;  
   wire [1:0] _io_imem_btb_update_bits_br_pc_T ;  
   wire [39:0] _GEN_250 ;  
   wire [39:0] _io_imem_btb_update_bits_br_pc_T_2 ;  
   wire [38:0] _io_imem_btb_update_bits_pc_T_1 ;  
   wire [5:0] ex_dcache_tag ;  
   wire [24:0] a_2 ;  
   wire _io_dmem_req_bits_addr_msb_T ;  
   wire _io_dmem_req_bits_addr_msb_T_1 ;  
   wire _io_dmem_req_bits_addr_msb_T_2 ;  
   wire msb_2 ;  
   wire [38:0] io_dmem_req_bits_addr_lo ;  
   wire _io_dmem_s1_kill_T ;  
   wire _unpause_T_1 ;  
   wire _unpause_T_2 ;  
   wire _unpause_T_3 ;  
   wire unpause ;  
   wire coreMonitorBundle_valid ;  
   wire coreMonitorBundle_wrenx ;  
   wire [5:0] _GEN_251 ;  
   wire [5:0] _T_142 ;  
   wire _T_145 ;  
   wire _T_146 ;  
   wire _T_147 ;  
   wire _T_153 ;  
   wire _T_159 ;  
   wire _GEN_254 ;  
   wire _GEN_256 ;  
   wire _GEN_257 ;  
   wire _GEN_261 ;  
   wire _GEN_262 ;  
   wire _GEN_268 ;  
   reg [19:0] Rocket_state ;  
   reg [31:0] _RAND_94 ;  
   reg Rocket_cov[0:1048575] ;  
   reg [31:0] _RAND_95 ;  
   wire Rocket_cov_read_data ;  
   wire [19:0] Rocket_cov_read_addr ;  
   wire Rocket_cov_write_data ;  
   wire [19:0] Rocket_cov_write_addr ;  
   wire Rocket_cov_write_mask ;  
   wire Rocket_cov_write_en ;  
   reg [29:0] Rocket_covSum ;  
   reg [31:0] _RAND_96 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire mux_cond_4 ;  
   wire mux_cond_5 ;  
   wire [10:0] ex_ctrl_wfd_shl ;  
   wire [19:0] ex_ctrl_wfd_pad ;  
   wire [15:0] ex_ctrl_fp_shl ;  
   wire [19:0] ex_ctrl_fp_pad ;  
   wire [15:0] mem_ctrl_jalr_shl ;  
   wire [19:0] mem_ctrl_jalr_pad ;  
   wire [11:0] wb_ctrl_mem_shl ;  
   wire [19:0] wb_ctrl_mem_pad ;  
   wire [6:0] ex_ctrl_wxd_shl ;  
   wire [19:0] ex_ctrl_wxd_pad ;  
   wire [19:0] ex_ctrl_mem_shl ;  
   wire [19:0] ex_ctrl_mem_pad ;  
   wire [19:0] ex_ctrl_sel_alu1_shl ;  
   wire [19:0] ex_ctrl_sel_alu1_pad ;  
   wire [11:0] mem_reg_replay_shl ;  
   wire [19:0] mem_reg_replay_pad ;  
   wire [16:0] blocked_shl ;  
   wire [19:0] blocked_pad ;  
   wire [2:0] wb_ctrl_div_shl ;  
   wire [19:0] wb_ctrl_div_pad ;  
   wire [15:0] wb_reg_flush_pipe_shl ;  
   wire [19:0] wb_reg_flush_pipe_pad ;  
   wire [11:0] mem_ctrl_jal_shl ;  
   wire [19:0] mem_ctrl_jal_pad ;  
   wire [9:0] ex_ctrl_sel_imm_shl ;  
   wire [19:0] ex_ctrl_sel_imm_pad ;  
   wire [8:0] wb_ctrl_wfd_shl ;  
   wire [19:0] wb_ctrl_wfd_pad ;  
   wire [19:0] mem_reg_slow_bypass_shl ;  
   wire [19:0] mem_reg_slow_bypass_pad ;  
   wire [16:0] mem_reg_sfence_shl ;  
   wire [19:0] mem_reg_sfence_pad ;  
   wire [2:0] wb_reg_xcpt_shl ;  
   wire [19:0] wb_reg_xcpt_pad ;  
   wire [15:0] id_reg_pause_shl ;  
   wire [19:0] id_reg_pause_pad ;  
   wire [8:0] ex_reg_rvc_shl ;  
   wire [19:0] ex_reg_rvc_pad ;  
   wire [3:0] wb_reg_valid_shl ;  
   wire [19:0] wb_reg_valid_pad ;  
   wire [13:0] mem_br_taken_shl ;  
   wire [19:0] mem_br_taken_pad ;  
   wire [18:0] mem_reg_flush_pipe_shl ;  
   wire [19:0] mem_reg_flush_pipe_pad ;  
   wire [17:0] ex_ctrl_div_shl ;  
   wire [19:0] ex_ctrl_div_pad ;  
   wire [15:0] mem_ctrl_fp_shl ;  
   wire [19:0] mem_ctrl_fp_pad ;  
   wire [5:0] mem_reg_xcpt_shl ;  
   wire [19:0] mem_reg_xcpt_pad ;  
   wire [14:0] mem_ctrl_wxd_shl ;  
   wire [19:0] mem_ctrl_wxd_pad ;  
   wire [8:0] mem_ctrl_mem_shl ;  
   wire [19:0] mem_ctrl_mem_pad ;  
   wire [16:0] ex_reg_mem_size_shl ;  
   wire [19:0] ex_reg_mem_size_pad ;  
   wire [8:0] ex_ctrl_sel_alu2_shl ;  
   wire [19:0] ex_ctrl_sel_alu2_pad ;  
   wire [2:0] ex_ctrl_rxs2_shl ;  
   wire [19:0] ex_ctrl_rxs2_pad ;  
   wire [3:0] ex_ctrl_jalr_shl ;  
   wire [19:0] ex_ctrl_jalr_pad ;  
   wire [4:0] ex_reg_replay_shl ;  
   wire [19:0] ex_reg_replay_pad ;  
   wire [3:0] ex_reg_valid_shl ;  
   wire [19:0] ex_reg_valid_pad ;  
   wire [6:0] mem_reg_valid_shl ;  
   wire [19:0] mem_reg_valid_pad ;  
   wire mem_reg_rvc_shl ;  
   wire [19:0] mem_reg_rvc_pad ;  
   wire mem_ctrl_wfd_shl ;  
   wire [19:0] mem_ctrl_wfd_pad ;  
   wire [11:0] id_reg_fence_shl ;  
   wire [19:0] id_reg_fence_pad ;  
   wire [8:0] mem_reg_load_shl ;  
   wire [19:0] mem_reg_load_pad ;  
   wire [18:0] wb_ctrl_wxd_shl ;  
   wire [19:0] wb_ctrl_wxd_pad ;  
   wire [1:0] wb_reg_replay_shl ;  
   wire [19:0] wb_reg_replay_pad ;  
   wire [10:0] ex_reg_xcpt_interrupt_shl ;  
   wire [19:0] ex_reg_xcpt_interrupt_pad ;  
   wire [6:0] mem_ctrl_branch_shl ;  
   wire [19:0] mem_ctrl_branch_pad ;  
   wire [1:0] mem_reg_xcpt_interrupt_shl ;  
   wire [19:0] mem_reg_xcpt_interrupt_pad ;  
   wire [4:0] mem_reg_store_shl ;  
   wire [19:0] mem_reg_store_pad ;  
   wire [5:0] mem_ctrl_div_shl ;  
   wire [19:0] mem_ctrl_div_pad ;  
   wire [17:0] mux_cond_0_shl ;  
   wire [19:0] mux_cond_0_pad ;  
   wire [8:0] mux_cond_1_shl ;  
   wire [19:0] mux_cond_1_pad ;  
   wire [15:0] mux_cond_2_shl ;  
   wire [19:0] mux_cond_2_pad ;  
   wire [4:0] mux_cond_3_shl ;  
   wire [19:0] mux_cond_3_pad ;  
   wire [9:0] mux_cond_4_shl ;  
   wire [19:0] mux_cond_4_pad ;  
   wire [17:0] mux_cond_5_shl ;  
   wire [19:0] mux_cond_5_pad ;  
   wire [12:0] ex_reg_rs_lsb_0_shl ;  
   wire [19:0] ex_reg_rs_lsb_0_pad ;  
   wire [12:0] ex_reg_rs_lsb_1_shl ;  
   wire [19:0] ex_reg_rs_lsb_1_pad ;  
   wire [10:0] ex_reg_rs_bypass_0_shl ;  
   wire [19:0] ex_reg_rs_bypass_0_pad ;  
   wire [10:0] ex_reg_rs_bypass_1_shl ;  
   wire [19:0] ex_reg_rs_bypass_1_pad ;  
   wire [19:0] Rocket_xor32 ;  
   wire [19:0] Rocket_xor15 ;  
   wire [19:0] Rocket_xor34 ;  
   wire [19:0] Rocket_xor16 ;  
   wire [19:0] Rocket_xor7 ;  
   wire [19:0] Rocket_xor36 ;  
   wire [19:0] Rocket_xor17 ;  
   wire [19:0] Rocket_xor37 ;  
   wire [19:0] Rocket_xor38 ;  
   wire [19:0] Rocket_xor18 ;  
   wire [19:0] Rocket_xor8 ;  
   wire [19:0] Rocket_xor3 ;  
   wire [19:0] Rocket_xor40 ;  
   wire [19:0] Rocket_xor19 ;  
   wire [19:0] Rocket_xor41 ;  
   wire [19:0] Rocket_xor42 ;  
   wire [19:0] Rocket_xor20 ;  
   wire [19:0] Rocket_xor9 ;  
   wire [19:0] Rocket_xor44 ;  
   wire [19:0] Rocket_xor21 ;  
   wire [19:0] Rocket_xor45 ;  
   wire [19:0] Rocket_xor46 ;  
   wire [19:0] Rocket_xor22 ;  
   wire [19:0] Rocket_xor10 ;  
   wire [19:0] Rocket_xor4 ;  
   wire [19:0] Rocket_xor1 ;  
   wire [19:0] Rocket_xor48 ;  
   wire [19:0] Rocket_xor23 ;  
   wire [19:0] Rocket_xor49 ;  
   wire [19:0] Rocket_xor50 ;  
   wire [19:0] Rocket_xor24 ;  
   wire [19:0] Rocket_xor11 ;  
   wire [19:0] Rocket_xor52 ;  
   wire [19:0] Rocket_xor25 ;  
   wire [19:0] Rocket_xor53 ;  
   wire [19:0] Rocket_xor54 ;  
   wire [19:0] Rocket_xor26 ;  
   wire [19:0] Rocket_xor12 ;  
   wire [19:0] Rocket_xor5 ;  
   wire [19:0] Rocket_xor56 ;  
   wire [19:0] Rocket_xor27 ;  
   wire [19:0] Rocket_xor57 ;  
   wire [19:0] Rocket_xor58 ;  
   wire [19:0] Rocket_xor28 ;  
   wire [19:0] Rocket_xor13 ;  
   wire [19:0] Rocket_xor60 ;  
   wire [19:0] Rocket_xor29 ;  
   wire [19:0] Rocket_xor61 ;  
   wire [19:0] Rocket_xor62 ;  
   wire [19:0] Rocket_xor30 ;  
   wire [19:0] Rocket_xor14 ;  
   wire [19:0] Rocket_xor6 ;  
   wire [19:0] Rocket_xor2 ;  
   wire [19:0] Rocket_xor0 ;  
   wire [29:0] PlusArgTimeout_sum ;  
   wire [29:0] csr_sum ;  
   wire [29:0] bpu_sum ;  
   wire [29:0] ibuf_sum ;  
   wire [29:0] div_sum ;  
   wire [29:0] alu_sum ;  
   wire alu_metaAssert_wire ;  
   wire div_metaAssert_wire ;  
   wire bpu_metaAssert_wire ;  
   wire PlusArgTimeout_metaAssert_wire ;  
   wire ibuf_metaAssert_wire ;  
   wire csr_metaAssert_wire ;  
   wire Rocket_or4 ;  
   wire Rocket_or1 ;  
   wire Rocket_or6 ;  
   wire Rocket_or2 ;  
   wire Rocket_or0 ;  
   reg Rocket_metaAssert ;  
   reg [31:0] _RAND_97 ;  
  IBuf ibuf(.clock(ibuf_clock),.reset(ibuf_reset),.io_imem_ready(ibuf_io_imem_ready),.io_imem_valid(ibuf_io_imem_valid),.io_imem_bits_btb_taken(ibuf_io_imem_bits_btb_taken),.io_imem_bits_btb_bridx(ibuf_io_imem_bits_btb_bridx),.io_imem_bits_btb_entry(ibuf_io_imem_bits_btb_entry),.io_imem_bits_btb_bht_history(ibuf_io_imem_bits_btb_bht_history),.io_imem_bits_pc(ibuf_io_imem_bits_pc),.io_imem_bits_data(ibuf_io_imem_bits_data),.io_imem_bits_xcpt_pf_inst(ibuf_io_imem_bits_xcpt_pf_inst),.io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),.io_imem_bits_replay(ibuf_io_imem_bits_replay),.io_kill(ibuf_io_kill),.io_pc(ibuf_io_pc),.io_btb_resp_entry(ibuf_io_btb_resp_entry),.io_btb_resp_bht_history(ibuf_io_btb_resp_bht_history),.io_inst_0_ready(ibuf_io_inst_0_ready),.io_inst_0_valid(ibuf_io_inst_0_valid),.io_inst_0_bits_xcpt0_pf_inst(ibuf_io_inst_0_bits_xcpt0_pf_inst),.io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),.io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),.io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),.io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),.io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),.io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),.io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),.io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),.io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),.io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3),.io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw),.io_covSum(ibuf_io_covSum),.metaAssert(ibuf_metaAssert),.metaReset(ibuf_metaReset)); 
  CSRFile csr(.clock(csr_clock),.reset(csr_reset),.io_ungated_clock(csr_io_ungated_clock),.io_interrupts_debug(csr_io_interrupts_debug),.io_interrupts_mtip(csr_io_interrupts_mtip),.io_interrupts_msip(csr_io_interrupts_msip),.io_interrupts_meip(csr_io_interrupts_meip),.io_interrupts_seip(csr_io_interrupts_seip),.io_hartid(csr_io_hartid),.io_rw_addr(csr_io_rw_addr),.io_rw_cmd(csr_io_rw_cmd),.io_rw_rdata(csr_io_rw_rdata),.io_rw_wdata(csr_io_rw_wdata),.io_decode_0_csr(csr_io_decode_0_csr),.io_decode_0_fp_illegal(csr_io_decode_0_fp_illegal),.io_decode_0_fp_csr(csr_io_decode_0_fp_csr),.io_decode_0_read_illegal(csr_io_decode_0_read_illegal),.io_decode_0_write_illegal(csr_io_decode_0_write_illegal),.io_decode_0_write_flush(csr_io_decode_0_write_flush),.io_decode_0_system_illegal(csr_io_decode_0_system_illegal),.io_csr_stall(csr_io_csr_stall),.io_eret(csr_io_eret),.io_singleStep(csr_io_singleStep),.io_status_debug(csr_io_status_debug),.io_status_cease(csr_io_status_cease),.io_status_wfi(csr_io_status_wfi),.io_status_isa(csr_io_status_isa),.io_status_dprv(csr_io_status_dprv),.io_status_prv(csr_io_status_prv),.io_status_sd(csr_io_status_sd),.io_status_zero2(csr_io_status_zero2),.io_status_sxl(csr_io_status_sxl),.io_status_uxl(csr_io_status_uxl),.io_status_sd_rv32(csr_io_status_sd_rv32),.io_status_zero1(csr_io_status_zero1),.io_status_tsr(csr_io_status_tsr),.io_status_tw(csr_io_status_tw),.io_status_tvm(csr_io_status_tvm),.io_status_mxr(csr_io_status_mxr),.io_status_sum(csr_io_status_sum),.io_status_mprv(csr_io_status_mprv),.io_status_xs(csr_io_status_xs),.io_status_fs(csr_io_status_fs),.io_status_mpp(csr_io_status_mpp),.io_status_vs(csr_io_status_vs),.io_status_spp(csr_io_status_spp),.io_status_mpie(csr_io_status_mpie),.io_status_hpie(csr_io_status_hpie),.io_status_spie(csr_io_status_spie),.io_status_upie(csr_io_status_upie),.io_status_mie(csr_io_status_mie),.io_status_hie(csr_io_status_hie),.io_status_sie(csr_io_status_sie),.io_status_uie(csr_io_status_uie),.io_ptbr_mode(csr_io_ptbr_mode),.io_ptbr_ppn(csr_io_ptbr_ppn),.io_evec(csr_io_evec),.io_exception(csr_io_exception),.io_retire(csr_io_retire),.io_cause(csr_io_cause),.io_pc(csr_io_pc),.io_tval(csr_io_tval),.io_time(csr_io_time),.io_fcsr_rm(csr_io_fcsr_rm),.io_fcsr_flags_valid(csr_io_fcsr_flags_valid),.io_fcsr_flags_bits(csr_io_fcsr_flags_bits),.io_interrupt(csr_io_interrupt),.io_interrupt_cause(csr_io_interrupt_cause),.io_bp_0_control_action(csr_io_bp_0_control_action),.io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),.io_bp_0_control_m(csr_io_bp_0_control_m),.io_bp_0_control_s(csr_io_bp_0_control_s),.io_bp_0_control_u(csr_io_bp_0_control_u),.io_bp_0_control_x(csr_io_bp_0_control_x),.io_bp_0_control_w(csr_io_bp_0_control_w),.io_bp_0_control_r(csr_io_bp_0_control_r),.io_bp_0_address(csr_io_bp_0_address),.io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),.io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),.io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),.io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),.io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),.io_pmp_0_addr(csr_io_pmp_0_addr),.io_pmp_0_mask(csr_io_pmp_0_mask),.io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),.io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),.io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),.io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),.io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),.io_pmp_1_addr(csr_io_pmp_1_addr),.io_pmp_1_mask(csr_io_pmp_1_mask),.io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),.io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),.io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),.io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),.io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),.io_pmp_2_addr(csr_io_pmp_2_addr),.io_pmp_2_mask(csr_io_pmp_2_mask),.io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),.io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),.io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),.io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),.io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),.io_pmp_3_addr(csr_io_pmp_3_addr),.io_pmp_3_mask(csr_io_pmp_3_mask),.io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),.io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),.io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),.io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),.io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),.io_pmp_4_addr(csr_io_pmp_4_addr),.io_pmp_4_mask(csr_io_pmp_4_mask),.io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),.io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),.io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),.io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),.io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),.io_pmp_5_addr(csr_io_pmp_5_addr),.io_pmp_5_mask(csr_io_pmp_5_mask),.io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),.io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),.io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),.io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),.io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),.io_pmp_6_addr(csr_io_pmp_6_addr),.io_pmp_6_mask(csr_io_pmp_6_mask),.io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),.io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),.io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),.io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),.io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),.io_pmp_7_addr(csr_io_pmp_7_addr),.io_pmp_7_mask(csr_io_pmp_7_mask),.io_inhibit_cycle(csr_io_inhibit_cycle),.io_inst_0(csr_io_inst_0),.io_trace_0_valid(csr_io_trace_0_valid),.io_trace_0_iaddr(csr_io_trace_0_iaddr),.io_trace_0_insn(csr_io_trace_0_insn),.io_trace_0_priv(csr_io_trace_0_priv),.io_trace_0_exception(csr_io_trace_0_exception),.io_trace_0_interrupt(csr_io_trace_0_interrupt),.io_trace_0_cause(csr_io_trace_0_cause),.io_trace_0_tval(csr_io_trace_0_tval),.io_customCSRs_0_value(csr_io_customCSRs_0_value),.io_covSum(csr_io_covSum),.metaAssert(csr_metaAssert),.metaReset(csr_metaReset)); 
  BreakpointUnit bpu(.io_status_debug(bpu_io_status_debug),.io_status_prv(bpu_io_status_prv),.io_bp_0_control_action(bpu_io_bp_0_control_action),.io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),.io_bp_0_control_m(bpu_io_bp_0_control_m),.io_bp_0_control_s(bpu_io_bp_0_control_s),.io_bp_0_control_u(bpu_io_bp_0_control_u),.io_bp_0_control_x(bpu_io_bp_0_control_x),.io_bp_0_control_w(bpu_io_bp_0_control_w),.io_bp_0_control_r(bpu_io_bp_0_control_r),.io_bp_0_address(bpu_io_bp_0_address),.io_pc(bpu_io_pc),.io_ea(bpu_io_ea),.io_xcpt_if(bpu_io_xcpt_if),.io_xcpt_ld(bpu_io_xcpt_ld),.io_xcpt_st(bpu_io_xcpt_st),.io_debug_if(bpu_io_debug_if),.io_debug_ld(bpu_io_debug_ld),.io_debug_st(bpu_io_debug_st),.io_covSum(bpu_io_covSum),.metaAssert(bpu_metaAssert)); 
  ALU alu(.io_dw(alu_io_dw),.io_fn(alu_io_fn),.io_in2(alu_io_in2),.io_in1(alu_io_in1),.io_out(alu_io_out),.io_adder_out(alu_io_adder_out),.io_cmp_out(alu_io_cmp_out),.io_covSum(alu_io_covSum),.metaAssert(alu_metaAssert)); 
  MulDiv div(.clock(div_clock),.reset(div_reset),.io_req_ready(div_io_req_ready),.io_req_valid(div_io_req_valid),.io_req_bits_fn(div_io_req_bits_fn),.io_req_bits_dw(div_io_req_bits_dw),.io_req_bits_in1(div_io_req_bits_in1),.io_req_bits_in2(div_io_req_bits_in2),.io_req_bits_tag(div_io_req_bits_tag),.io_kill(div_io_kill),.io_resp_ready(div_io_resp_ready),.io_resp_valid(div_io_resp_valid),.io_resp_bits_data(div_io_resp_bits_data),.io_resp_bits_tag(div_io_resp_bits_tag),.io_covSum(div_io_covSum),.metaAssert(div_metaAssert),.metaReset(div_metaReset)); 
  PlusArgTimeout PlusArgTimeout(.clock(PlusArgTimeout_clock),.reset(PlusArgTimeout_reset),.io_count(PlusArgTimeout_io_count),.io_covSum(PlusArgTimeout_io_covSum),.metaAssert(PlusArgTimeout_metaAssert),.metaReset(PlusArgTimeout_metaReset)); 
  assign rf_id_rs_MPORT_addr=~id_raddr1; 
  assign rf_id_rs_MPORT_data=rf[rf_id_rs_MPORT_addr]; 
  assign rf_id_rs_MPORT_1_addr=~id_raddr2; 
  assign rf_id_rs_MPORT_1_data=rf[rf_id_rs_MPORT_1_addr]; 
  assign rf_MPORT_data=_rf_wdata_T ? io_dmem_resp_bits_data:_rf_wdata_T_5; 
  assign rf_MPORT_addr=~rf_waddr; 
  assign rf_MPORT_mask=1'h1; 
  assign rf_MPORT_en=rf_wen&_T_118; 
  assign replay_wb_common=io_dmem_s2_nack|wb_reg_replay; 
  assign _T_83=wb_reg_valid&wb_ctrl_mem; 
  assign _T_84=_T_83&io_dmem_s2_xcpt_ma_st; 
  assign _T_95=wb_reg_xcpt|_T_84; 
  assign _T_86=_T_83&io_dmem_s2_xcpt_ma_ld; 
  assign _T_96=_T_95|_T_86; 
  assign _T_88=_T_83&io_dmem_s2_xcpt_pf_st; 
  assign _T_97=_T_96|_T_88; 
  assign _T_90=_T_83&io_dmem_s2_xcpt_pf_ld; 
  assign _T_98=_T_97|_T_90; 
  assign _T_92=_T_83&io_dmem_s2_xcpt_ae_st; 
  assign _T_99=_T_98|_T_92; 
  assign _T_94=_T_83&io_dmem_s2_xcpt_ae_ld; 
  assign wb_xcpt=_T_99|_T_94; 
  assign _take_pc_wb_T=replay_wb_common|wb_xcpt; 
  assign _take_pc_wb_T_1=_take_pc_wb_T|csr_io_eret; 
  assign take_pc_wb=_take_pc_wb_T_1|wb_reg_flush_pipe; 
  assign _ex_pc_valid_T=ex_reg_valid|ex_reg_replay; 
  assign ex_pc_valid=_ex_pc_valid_T|ex_reg_xcpt_interrupt; 
  assign _mem_npc_T=mem_ctrl_jalr|mem_reg_sfence; 
  assign a=mem_reg_wdata[63:39]; 
  assign _mem_npc_msb_T=$signed(a)==25'sh0; 
  assign _mem_npc_msb_T_1=$signed(a)==-25'sh1; 
  assign _mem_npc_msb_T_2=_mem_npc_msb_T|_mem_npc_msb_T_1; 
  assign msb=_mem_npc_msb_T_2 ? mem_reg_wdata[39]:~mem_reg_wdata[38]; 
  assign mem_npc_lo=mem_reg_wdata[38:0]; 
  assign _mem_npc_T_2={msb,mem_npc_lo}; 
  assign _mem_br_target_T_1=mem_ctrl_branch&mem_br_taken; 
  assign mem_br_target_sign=mem_reg_inst[31]; 
  assign mem_br_target_hi_hi_hi=mem_reg_inst[31]; 
  assign mem_br_target_hi_hi_lo={11{mem_br_target_sign}}; 
  assign mem_br_target_hi_lo_hi={8{mem_br_target_sign}}; 
  assign mem_br_target_hi_lo_lo=mem_reg_inst[7]; 
  assign mem_br_target_lo_hi_hi=mem_reg_inst[30:25]; 
  assign mem_br_target_lo_hi_lo=mem_reg_inst[11:8]; 
  assign _mem_br_target_T_3={mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi,mem_br_target_hi_lo_lo,mem_br_target_lo_hi_hi,mem_br_target_lo_hi_lo,1'h0}; 
  assign mem_br_target_hi_lo_hi_1=mem_reg_inst[19:12]; 
  assign mem_br_target_hi_lo_lo_1=mem_reg_inst[20]; 
  assign _mem_br_target_T_5={mem_br_target_hi_hi_hi,mem_br_target_hi_hi_lo,mem_br_target_hi_lo_hi_1,mem_br_target_hi_lo_lo_1,mem_br_target_lo_hi_hi,mem_reg_inst[24:21],1'h0}; 
  assign _mem_br_target_T_6=mem_reg_rvc ? $signed(4'sh2):$signed(4'sh4); 
  assign _mem_br_target_T_7=mem_ctrl_jal ? $signed(_mem_br_target_T_5):$signed({{28{_mem_br_target_T_6[3]}},_mem_br_target_T_6}); 
  assign _mem_br_target_T_8=_mem_br_target_T_1 ? $signed(_mem_br_target_T_3):$signed(_mem_br_target_T_7); 
  assign _GEN_248={{8{_mem_br_target_T_8[31]}},_mem_br_target_T_8}; 
  assign mem_br_target=$signed(mem_reg_pc)+$signed(_GEN_248); 
  assign _mem_npc_T_3=_mem_npc_T ? $signed(_mem_npc_T_2):$signed(mem_br_target); 
  assign mem_npc=$signed(_mem_npc_T_3)&-40'sh2; 
  assign _mem_wrong_npc_T=mem_npc!=ex_reg_pc; 
  assign _mem_wrong_npc_T_1=ibuf_io_inst_0_valid|ibuf_io_imem_valid; 
  assign _mem_wrong_npc_T_2=mem_npc!=ibuf_io_pc; 
  assign _mem_wrong_npc_T_3=_mem_wrong_npc_T_1 ? _mem_wrong_npc_T_2:1'h1; 
  assign mem_wrong_npc=ex_pc_valid ? _mem_wrong_npc_T:_mem_wrong_npc_T_3; 
  assign _take_pc_mem_T=mem_wrong_npc|mem_reg_sfence; 
  assign take_pc_mem=mem_reg_valid&_take_pc_mem_T; 
  assign take_pc_mem_wb=take_pc_wb|take_pc_mem; 
  assign _id_ctrl_decoder_bit_T=ibuf_io_inst_0_bits_inst_bits&32'hfe00707f; 
  assign _id_ctrl_decoder_bit_T_1=_id_ctrl_decoder_bit_T==32'h2000033; 
  assign _id_ctrl_decoder_bit_T_3=_id_ctrl_decoder_bit_T==32'h2001033; 
  assign _id_ctrl_decoder_bit_T_5=_id_ctrl_decoder_bit_T==32'h2003033; 
  assign _id_ctrl_decoder_bit_T_7=_id_ctrl_decoder_bit_T==32'h2002033; 
  assign _id_ctrl_decoder_bit_T_9=_id_ctrl_decoder_bit_T==32'h2004033; 
  assign _id_ctrl_decoder_bit_T_11=_id_ctrl_decoder_bit_T==32'h2005033; 
  assign _id_ctrl_decoder_bit_T_13=_id_ctrl_decoder_bit_T==32'h2006033; 
  assign _id_ctrl_decoder_bit_T_15=_id_ctrl_decoder_bit_T==32'h2007033; 
  assign _id_ctrl_decoder_bit_T_17=_id_ctrl_decoder_bit_T==32'h200003b; 
  assign _id_ctrl_decoder_bit_T_19=_id_ctrl_decoder_bit_T==32'h200403b; 
  assign _id_ctrl_decoder_bit_T_21=_id_ctrl_decoder_bit_T==32'h200503b; 
  assign _id_ctrl_decoder_bit_T_23=_id_ctrl_decoder_bit_T==32'h200603b; 
  assign _id_ctrl_decoder_bit_T_25=_id_ctrl_decoder_bit_T==32'h200703b; 
  assign _id_ctrl_decoder_bit_T_26=ibuf_io_inst_0_bits_inst_bits&32'hf800707f; 
  assign _id_ctrl_decoder_bit_T_27=_id_ctrl_decoder_bit_T_26==32'h202f; 
  assign _id_ctrl_decoder_bit_T_29=_id_ctrl_decoder_bit_T_26==32'h2000202f; 
  assign _id_ctrl_decoder_bit_T_31=_id_ctrl_decoder_bit_T_26==32'h800202f; 
  assign _id_ctrl_decoder_bit_T_33=_id_ctrl_decoder_bit_T_26==32'h6000202f; 
  assign _id_ctrl_decoder_bit_T_35=_id_ctrl_decoder_bit_T_26==32'h4000202f; 
  assign _id_ctrl_decoder_bit_T_37=_id_ctrl_decoder_bit_T_26==32'h8000202f; 
  assign _id_ctrl_decoder_bit_T_39=_id_ctrl_decoder_bit_T_26==32'hc000202f; 
  assign _id_ctrl_decoder_bit_T_41=_id_ctrl_decoder_bit_T_26==32'ha000202f; 
  assign _id_ctrl_decoder_bit_T_43=_id_ctrl_decoder_bit_T_26==32'he000202f; 
  assign _id_ctrl_decoder_bit_T_44=ibuf_io_inst_0_bits_inst_bits&32'hf9f0707f; 
  assign _id_ctrl_decoder_bit_T_45=_id_ctrl_decoder_bit_T_44==32'h1000202f; 
  assign _id_ctrl_decoder_bit_T_47=_id_ctrl_decoder_bit_T_26==32'h1800202f; 
  assign _id_ctrl_decoder_bit_T_49=_id_ctrl_decoder_bit_T_26==32'h302f; 
  assign _id_ctrl_decoder_bit_T_51=_id_ctrl_decoder_bit_T_26==32'h800302f; 
  assign _id_ctrl_decoder_bit_T_53=_id_ctrl_decoder_bit_T_26==32'h2000302f; 
  assign _id_ctrl_decoder_bit_T_55=_id_ctrl_decoder_bit_T_26==32'h6000302f; 
  assign _id_ctrl_decoder_bit_T_57=_id_ctrl_decoder_bit_T_26==32'h4000302f; 
  assign _id_ctrl_decoder_bit_T_59=_id_ctrl_decoder_bit_T_26==32'h8000302f; 
  assign _id_ctrl_decoder_bit_T_61=_id_ctrl_decoder_bit_T_26==32'hc000302f; 
  assign _id_ctrl_decoder_bit_T_63=_id_ctrl_decoder_bit_T_26==32'ha000302f; 
  assign _id_ctrl_decoder_bit_T_65=_id_ctrl_decoder_bit_T_26==32'he000302f; 
  assign _id_ctrl_decoder_bit_T_67=_id_ctrl_decoder_bit_T_44==32'h1000302f; 
  assign _id_ctrl_decoder_bit_T_69=_id_ctrl_decoder_bit_T_26==32'h1800302f; 
  assign _id_ctrl_decoder_bit_T_71=_id_ctrl_decoder_bit_T==32'h20000053; 
  assign _id_ctrl_decoder_bit_T_73=_id_ctrl_decoder_bit_T==32'h20002053; 
  assign _id_ctrl_decoder_bit_T_75=_id_ctrl_decoder_bit_T==32'h20001053; 
  assign _id_ctrl_decoder_bit_T_77=_id_ctrl_decoder_bit_T==32'h28000053; 
  assign _id_ctrl_decoder_bit_T_79=_id_ctrl_decoder_bit_T==32'h28001053; 
  assign _id_ctrl_decoder_bit_T_80=ibuf_io_inst_0_bits_inst_bits&32'hfe00007f; 
  assign _id_ctrl_decoder_bit_T_81=_id_ctrl_decoder_bit_T_80==32'h53; 
  assign _id_ctrl_decoder_bit_T_83=_id_ctrl_decoder_bit_T_80==32'h8000053; 
  assign _id_ctrl_decoder_bit_T_85=_id_ctrl_decoder_bit_T_80==32'h10000053; 
  assign _id_ctrl_decoder_bit_T_86=ibuf_io_inst_0_bits_inst_bits&32'h600007f; 
  assign _id_ctrl_decoder_bit_T_87=_id_ctrl_decoder_bit_T_86==32'h43; 
  assign _id_ctrl_decoder_bit_T_89=_id_ctrl_decoder_bit_T_86==32'h47; 
  assign _id_ctrl_decoder_bit_T_91=_id_ctrl_decoder_bit_T_86==32'h4f; 
  assign _id_ctrl_decoder_bit_T_93=_id_ctrl_decoder_bit_T_86==32'h4b; 
  assign _id_ctrl_decoder_bit_T_94=ibuf_io_inst_0_bits_inst_bits&32'hfff0707f; 
  assign _id_ctrl_decoder_bit_T_95=_id_ctrl_decoder_bit_T_94==32'he0001053; 
  assign _id_ctrl_decoder_bit_T_97=_id_ctrl_decoder_bit_T_94==32'he0000053; 
  assign _id_ctrl_decoder_bit_T_98=ibuf_io_inst_0_bits_inst_bits&32'hfff0007f; 
  assign _id_ctrl_decoder_bit_T_99=_id_ctrl_decoder_bit_T_98==32'hc0000053; 
  assign _id_ctrl_decoder_bit_T_101=_id_ctrl_decoder_bit_T_98==32'hc0100053; 
  assign _id_ctrl_decoder_bit_T_103=_id_ctrl_decoder_bit_T==32'ha0002053; 
  assign _id_ctrl_decoder_bit_T_105=_id_ctrl_decoder_bit_T==32'ha0001053; 
  assign _id_ctrl_decoder_bit_T_107=_id_ctrl_decoder_bit_T==32'ha0000053; 
  assign _id_ctrl_decoder_bit_T_109=_id_ctrl_decoder_bit_T_94==32'hf0000053; 
  assign _id_ctrl_decoder_bit_T_111=_id_ctrl_decoder_bit_T_98==32'hd0000053; 
  assign _id_ctrl_decoder_bit_T_113=_id_ctrl_decoder_bit_T_98==32'hd0100053; 
  assign _id_ctrl_decoder_bit_T_114=ibuf_io_inst_0_bits_inst_bits&32'h707f; 
  assign _id_ctrl_decoder_bit_T_115=_id_ctrl_decoder_bit_T_114==32'h2007; 
  assign _id_ctrl_decoder_bit_T_117=_id_ctrl_decoder_bit_T_114==32'h2027; 
  assign _id_ctrl_decoder_bit_T_119=_id_ctrl_decoder_bit_T_80==32'h18000053; 
  assign _id_ctrl_decoder_bit_T_121=_id_ctrl_decoder_bit_T_98==32'h58000053; 
  assign _id_ctrl_decoder_bit_T_123=_id_ctrl_decoder_bit_T_98==32'hc0200053; 
  assign _id_ctrl_decoder_bit_T_125=_id_ctrl_decoder_bit_T_98==32'hc0300053; 
  assign _id_ctrl_decoder_bit_T_127=_id_ctrl_decoder_bit_T_98==32'hd0200053; 
  assign _id_ctrl_decoder_bit_T_129=_id_ctrl_decoder_bit_T_98==32'hd0300053; 
  assign _id_ctrl_decoder_bit_T_131=_id_ctrl_decoder_bit_T_98==32'h40100053; 
  assign _id_ctrl_decoder_bit_T_133=_id_ctrl_decoder_bit_T_98==32'h42000053; 
  assign _id_ctrl_decoder_bit_T_135=_id_ctrl_decoder_bit_T==32'h22000053; 
  assign _id_ctrl_decoder_bit_T_137=_id_ctrl_decoder_bit_T==32'h22002053; 
  assign _id_ctrl_decoder_bit_T_139=_id_ctrl_decoder_bit_T==32'h22001053; 
  assign _id_ctrl_decoder_bit_T_141=_id_ctrl_decoder_bit_T==32'h2a000053; 
  assign _id_ctrl_decoder_bit_T_143=_id_ctrl_decoder_bit_T==32'h2a001053; 
  assign _id_ctrl_decoder_bit_T_145=_id_ctrl_decoder_bit_T_80==32'h2000053; 
  assign _id_ctrl_decoder_bit_T_147=_id_ctrl_decoder_bit_T_80==32'ha000053; 
  assign _id_ctrl_decoder_bit_T_149=_id_ctrl_decoder_bit_T_80==32'h12000053; 
  assign _id_ctrl_decoder_bit_T_151=_id_ctrl_decoder_bit_T_86==32'h2000043; 
  assign _id_ctrl_decoder_bit_T_153=_id_ctrl_decoder_bit_T_86==32'h2000047; 
  assign _id_ctrl_decoder_bit_T_155=_id_ctrl_decoder_bit_T_86==32'h200004f; 
  assign _id_ctrl_decoder_bit_T_157=_id_ctrl_decoder_bit_T_86==32'h200004b; 
  assign _id_ctrl_decoder_bit_T_159=_id_ctrl_decoder_bit_T_94==32'he2001053; 
  assign _id_ctrl_decoder_bit_T_161=_id_ctrl_decoder_bit_T_98==32'hc2000053; 
  assign _id_ctrl_decoder_bit_T_163=_id_ctrl_decoder_bit_T_98==32'hc2100053; 
  assign _id_ctrl_decoder_bit_T_165=_id_ctrl_decoder_bit_T==32'ha2002053; 
  assign _id_ctrl_decoder_bit_T_167=_id_ctrl_decoder_bit_T==32'ha2001053; 
  assign _id_ctrl_decoder_bit_T_169=_id_ctrl_decoder_bit_T==32'ha2000053; 
  assign _id_ctrl_decoder_bit_T_171=_id_ctrl_decoder_bit_T_98==32'hd2000053; 
  assign _id_ctrl_decoder_bit_T_173=_id_ctrl_decoder_bit_T_98==32'hd2100053; 
  assign _id_ctrl_decoder_bit_T_175=_id_ctrl_decoder_bit_T_114==32'h3007; 
  assign _id_ctrl_decoder_bit_T_177=_id_ctrl_decoder_bit_T_114==32'h3027; 
  assign _id_ctrl_decoder_bit_T_179=_id_ctrl_decoder_bit_T_80==32'h1a000053; 
  assign _id_ctrl_decoder_bit_T_181=_id_ctrl_decoder_bit_T_98==32'h5a000053; 
  assign _id_ctrl_decoder_bit_T_183=_id_ctrl_decoder_bit_T_94==32'he2000053; 
  assign _id_ctrl_decoder_bit_T_185=_id_ctrl_decoder_bit_T_98==32'hc2200053; 
  assign _id_ctrl_decoder_bit_T_187=_id_ctrl_decoder_bit_T_98==32'hc2300053; 
  assign _id_ctrl_decoder_bit_T_189=_id_ctrl_decoder_bit_T_94==32'hf2000053; 
  assign _id_ctrl_decoder_bit_T_191=_id_ctrl_decoder_bit_T_98==32'hd2200053; 
  assign _id_ctrl_decoder_bit_T_193=_id_ctrl_decoder_bit_T_98==32'hd2300053; 
  assign _id_ctrl_decoder_bit_T_195=_id_ctrl_decoder_bit_T_114==32'h3003; 
  assign _id_ctrl_decoder_bit_T_197=_id_ctrl_decoder_bit_T_114==32'h6003; 
  assign _id_ctrl_decoder_bit_T_199=_id_ctrl_decoder_bit_T_114==32'h3023; 
  assign _id_ctrl_decoder_bit_T_200=ibuf_io_inst_0_bits_inst_bits&32'hfc00707f; 
  assign _id_ctrl_decoder_bit_T_201=_id_ctrl_decoder_bit_T_200==32'h1013; 
  assign _id_ctrl_decoder_bit_T_203=_id_ctrl_decoder_bit_T_200==32'h5013; 
  assign _id_ctrl_decoder_bit_T_205=_id_ctrl_decoder_bit_T_200==32'h40005013; 
  assign _id_ctrl_decoder_bit_T_207=_id_ctrl_decoder_bit_T_114==32'h1b; 
  assign _id_ctrl_decoder_bit_T_209=_id_ctrl_decoder_bit_T==32'h101b; 
  assign _id_ctrl_decoder_bit_T_211=_id_ctrl_decoder_bit_T==32'h501b; 
  assign _id_ctrl_decoder_bit_T_213=_id_ctrl_decoder_bit_T==32'h4000501b; 
  assign _id_ctrl_decoder_bit_T_215=_id_ctrl_decoder_bit_T==32'h3b; 
  assign _id_ctrl_decoder_bit_T_217=_id_ctrl_decoder_bit_T==32'h4000003b; 
  assign _id_ctrl_decoder_bit_T_219=_id_ctrl_decoder_bit_T==32'h103b; 
  assign _id_ctrl_decoder_bit_T_221=_id_ctrl_decoder_bit_T==32'h503b; 
  assign _id_ctrl_decoder_bit_T_223=_id_ctrl_decoder_bit_T==32'h4000503b; 
  assign _id_ctrl_decoder_bit_T_224=ibuf_io_inst_0_bits_inst_bits&32'hfe007fff; 
  assign _id_ctrl_decoder_bit_T_225=_id_ctrl_decoder_bit_T_224==32'h12000073; 
  assign _id_ctrl_decoder_bit_T_226=ibuf_io_inst_0_bits_inst_bits==32'h10200073; 
  assign _id_ctrl_decoder_bit_T_227=ibuf_io_inst_0_bits_inst_bits==32'h7b200073; 
  assign _id_ctrl_decoder_bit_T_229=_id_ctrl_decoder_bit_T_114==32'h100f; 
  assign _id_ctrl_decoder_bit_T_231=_id_ctrl_decoder_bit_T_114==32'h1063; 
  assign _id_ctrl_decoder_bit_T_233=_id_ctrl_decoder_bit_T_114==32'h63; 
  assign _id_ctrl_decoder_bit_T_235=_id_ctrl_decoder_bit_T_114==32'h4063; 
  assign _id_ctrl_decoder_bit_T_237=_id_ctrl_decoder_bit_T_114==32'h6063; 
  assign _id_ctrl_decoder_bit_T_239=_id_ctrl_decoder_bit_T_114==32'h5063; 
  assign _id_ctrl_decoder_bit_T_241=_id_ctrl_decoder_bit_T_114==32'h7063; 
  assign _id_ctrl_decoder_bit_T_242=ibuf_io_inst_0_bits_inst_bits&32'h7f; 
  assign _id_ctrl_decoder_bit_T_243=_id_ctrl_decoder_bit_T_242==32'h6f; 
  assign _id_ctrl_decoder_bit_T_245=_id_ctrl_decoder_bit_T_114==32'h67; 
  assign _id_ctrl_decoder_bit_T_247=_id_ctrl_decoder_bit_T_242==32'h17; 
  assign _id_ctrl_decoder_bit_T_249=_id_ctrl_decoder_bit_T_114==32'h3; 
  assign _id_ctrl_decoder_bit_T_251=_id_ctrl_decoder_bit_T_114==32'h1003; 
  assign _id_ctrl_decoder_bit_T_253=_id_ctrl_decoder_bit_T_114==32'h2003; 
  assign _id_ctrl_decoder_bit_T_255=_id_ctrl_decoder_bit_T_114==32'h4003; 
  assign _id_ctrl_decoder_bit_T_257=_id_ctrl_decoder_bit_T_114==32'h5003; 
  assign _id_ctrl_decoder_bit_T_259=_id_ctrl_decoder_bit_T_114==32'h23; 
  assign _id_ctrl_decoder_bit_T_261=_id_ctrl_decoder_bit_T_114==32'h1023; 
  assign _id_ctrl_decoder_bit_T_263=_id_ctrl_decoder_bit_T_114==32'h2023; 
  assign _id_ctrl_decoder_bit_T_265=_id_ctrl_decoder_bit_T_242==32'h37; 
  assign _id_ctrl_decoder_bit_T_267=_id_ctrl_decoder_bit_T_114==32'h13; 
  assign _id_ctrl_decoder_bit_T_269=_id_ctrl_decoder_bit_T_114==32'h2013; 
  assign _id_ctrl_decoder_bit_T_271=_id_ctrl_decoder_bit_T_114==32'h3013; 
  assign _id_ctrl_decoder_bit_T_273=_id_ctrl_decoder_bit_T_114==32'h7013; 
  assign _id_ctrl_decoder_bit_T_275=_id_ctrl_decoder_bit_T_114==32'h6013; 
  assign _id_ctrl_decoder_bit_T_277=_id_ctrl_decoder_bit_T_114==32'h4013; 
  assign _id_ctrl_decoder_bit_T_279=_id_ctrl_decoder_bit_T==32'h33; 
  assign _id_ctrl_decoder_bit_T_281=_id_ctrl_decoder_bit_T==32'h40000033; 
  assign _id_ctrl_decoder_bit_T_283=_id_ctrl_decoder_bit_T==32'h2033; 
  assign _id_ctrl_decoder_bit_T_285=_id_ctrl_decoder_bit_T==32'h3033; 
  assign _id_ctrl_decoder_bit_T_287=_id_ctrl_decoder_bit_T==32'h7033; 
  assign _id_ctrl_decoder_bit_T_289=_id_ctrl_decoder_bit_T==32'h6033; 
  assign _id_ctrl_decoder_bit_T_291=_id_ctrl_decoder_bit_T==32'h4033; 
  assign _id_ctrl_decoder_bit_T_293=_id_ctrl_decoder_bit_T==32'h1033; 
  assign _id_ctrl_decoder_bit_T_295=_id_ctrl_decoder_bit_T==32'h5033; 
  assign _id_ctrl_decoder_bit_T_297=_id_ctrl_decoder_bit_T==32'h40005033; 
  assign _id_ctrl_decoder_bit_T_299=_id_ctrl_decoder_bit_T_114==32'hf; 
  assign _id_ctrl_decoder_bit_T_300=ibuf_io_inst_0_bits_inst_bits==32'h73; 
  assign _id_ctrl_decoder_bit_T_301=ibuf_io_inst_0_bits_inst_bits==32'h100073; 
  assign _id_ctrl_decoder_bit_T_302=ibuf_io_inst_0_bits_inst_bits==32'h30200073; 
  assign _id_ctrl_decoder_bit_T_303=ibuf_io_inst_0_bits_inst_bits==32'h10500073; 
  assign _id_ctrl_decoder_bit_T_304=ibuf_io_inst_0_bits_inst_bits==32'h30500073; 
  assign _id_ctrl_decoder_bit_T_306=_id_ctrl_decoder_bit_T_114==32'h1073; 
  assign _id_ctrl_decoder_bit_T_308=_id_ctrl_decoder_bit_T_114==32'h2073; 
  assign _id_ctrl_decoder_bit_T_310=_id_ctrl_decoder_bit_T_114==32'h3073; 
  assign _id_ctrl_decoder_bit_T_312=_id_ctrl_decoder_bit_T_114==32'h5073; 
  assign _id_ctrl_decoder_bit_T_314=_id_ctrl_decoder_bit_T_114==32'h6073; 
  assign _id_ctrl_decoder_bit_T_316=_id_ctrl_decoder_bit_T_114==32'h7073; 
  assign _id_ctrl_decoder_bit_T_318=_id_ctrl_decoder_bit_T_1|_id_ctrl_decoder_bit_T_3; 
  assign _id_ctrl_decoder_bit_T_319=_id_ctrl_decoder_bit_T_318|_id_ctrl_decoder_bit_T_5; 
  assign _id_ctrl_decoder_bit_T_320=_id_ctrl_decoder_bit_T_319|_id_ctrl_decoder_bit_T_7; 
  assign _id_ctrl_decoder_bit_T_321=_id_ctrl_decoder_bit_T_320|_id_ctrl_decoder_bit_T_9; 
  assign _id_ctrl_decoder_bit_T_322=_id_ctrl_decoder_bit_T_321|_id_ctrl_decoder_bit_T_11; 
  assign _id_ctrl_decoder_bit_T_323=_id_ctrl_decoder_bit_T_322|_id_ctrl_decoder_bit_T_13; 
  assign _id_ctrl_decoder_bit_T_324=_id_ctrl_decoder_bit_T_323|_id_ctrl_decoder_bit_T_15; 
  assign _id_ctrl_decoder_bit_T_325=_id_ctrl_decoder_bit_T_324|_id_ctrl_decoder_bit_T_17; 
  assign _id_ctrl_decoder_bit_T_326=_id_ctrl_decoder_bit_T_325|_id_ctrl_decoder_bit_T_19; 
  assign _id_ctrl_decoder_bit_T_327=_id_ctrl_decoder_bit_T_326|_id_ctrl_decoder_bit_T_21; 
  assign _id_ctrl_decoder_bit_T_328=_id_ctrl_decoder_bit_T_327|_id_ctrl_decoder_bit_T_23; 
  assign _id_ctrl_decoder_bit_T_329=_id_ctrl_decoder_bit_T_328|_id_ctrl_decoder_bit_T_25; 
  assign _id_ctrl_decoder_bit_T_330=_id_ctrl_decoder_bit_T_329|_id_ctrl_decoder_bit_T_27; 
  assign _id_ctrl_decoder_bit_T_331=_id_ctrl_decoder_bit_T_330|_id_ctrl_decoder_bit_T_29; 
  assign _id_ctrl_decoder_bit_T_332=_id_ctrl_decoder_bit_T_331|_id_ctrl_decoder_bit_T_31; 
  assign _id_ctrl_decoder_bit_T_333=_id_ctrl_decoder_bit_T_332|_id_ctrl_decoder_bit_T_33; 
  assign _id_ctrl_decoder_bit_T_334=_id_ctrl_decoder_bit_T_333|_id_ctrl_decoder_bit_T_35; 
  assign _id_ctrl_decoder_bit_T_335=_id_ctrl_decoder_bit_T_334|_id_ctrl_decoder_bit_T_37; 
  assign _id_ctrl_decoder_bit_T_336=_id_ctrl_decoder_bit_T_335|_id_ctrl_decoder_bit_T_39; 
  assign _id_ctrl_decoder_bit_T_337=_id_ctrl_decoder_bit_T_336|_id_ctrl_decoder_bit_T_41; 
  assign _id_ctrl_decoder_bit_T_338=_id_ctrl_decoder_bit_T_337|_id_ctrl_decoder_bit_T_43; 
  assign _id_ctrl_decoder_bit_T_339=_id_ctrl_decoder_bit_T_338|_id_ctrl_decoder_bit_T_45; 
  assign _id_ctrl_decoder_bit_T_340=_id_ctrl_decoder_bit_T_339|_id_ctrl_decoder_bit_T_47; 
  assign _id_ctrl_decoder_bit_T_341=_id_ctrl_decoder_bit_T_340|_id_ctrl_decoder_bit_T_49; 
  assign _id_ctrl_decoder_bit_T_342=_id_ctrl_decoder_bit_T_341|_id_ctrl_decoder_bit_T_51; 
  assign _id_ctrl_decoder_bit_T_343=_id_ctrl_decoder_bit_T_342|_id_ctrl_decoder_bit_T_53; 
  assign _id_ctrl_decoder_bit_T_344=_id_ctrl_decoder_bit_T_343|_id_ctrl_decoder_bit_T_55; 
  assign _id_ctrl_decoder_bit_T_345=_id_ctrl_decoder_bit_T_344|_id_ctrl_decoder_bit_T_57; 
  assign _id_ctrl_decoder_bit_T_346=_id_ctrl_decoder_bit_T_345|_id_ctrl_decoder_bit_T_59; 
  assign _id_ctrl_decoder_bit_T_347=_id_ctrl_decoder_bit_T_346|_id_ctrl_decoder_bit_T_61; 
  assign _id_ctrl_decoder_bit_T_348=_id_ctrl_decoder_bit_T_347|_id_ctrl_decoder_bit_T_63; 
  assign _id_ctrl_decoder_bit_T_349=_id_ctrl_decoder_bit_T_348|_id_ctrl_decoder_bit_T_65; 
  assign _id_ctrl_decoder_bit_T_350=_id_ctrl_decoder_bit_T_349|_id_ctrl_decoder_bit_T_67; 
  assign _id_ctrl_decoder_bit_T_351=_id_ctrl_decoder_bit_T_350|_id_ctrl_decoder_bit_T_69; 
  assign _id_ctrl_decoder_bit_T_352=_id_ctrl_decoder_bit_T_351|_id_ctrl_decoder_bit_T_71; 
  assign _id_ctrl_decoder_bit_T_353=_id_ctrl_decoder_bit_T_352|_id_ctrl_decoder_bit_T_73; 
  assign _id_ctrl_decoder_bit_T_354=_id_ctrl_decoder_bit_T_353|_id_ctrl_decoder_bit_T_75; 
  assign _id_ctrl_decoder_bit_T_355=_id_ctrl_decoder_bit_T_354|_id_ctrl_decoder_bit_T_77; 
  assign _id_ctrl_decoder_bit_T_356=_id_ctrl_decoder_bit_T_355|_id_ctrl_decoder_bit_T_79; 
  assign _id_ctrl_decoder_bit_T_357=_id_ctrl_decoder_bit_T_356|_id_ctrl_decoder_bit_T_81; 
  assign _id_ctrl_decoder_bit_T_358=_id_ctrl_decoder_bit_T_357|_id_ctrl_decoder_bit_T_83; 
  assign _id_ctrl_decoder_bit_T_359=_id_ctrl_decoder_bit_T_358|_id_ctrl_decoder_bit_T_85; 
  assign _id_ctrl_decoder_bit_T_360=_id_ctrl_decoder_bit_T_359|_id_ctrl_decoder_bit_T_87; 
  assign _id_ctrl_decoder_bit_T_361=_id_ctrl_decoder_bit_T_360|_id_ctrl_decoder_bit_T_89; 
  assign _id_ctrl_decoder_bit_T_362=_id_ctrl_decoder_bit_T_361|_id_ctrl_decoder_bit_T_91; 
  assign _id_ctrl_decoder_bit_T_363=_id_ctrl_decoder_bit_T_362|_id_ctrl_decoder_bit_T_93; 
  assign _id_ctrl_decoder_bit_T_364=_id_ctrl_decoder_bit_T_363|_id_ctrl_decoder_bit_T_95; 
  assign _id_ctrl_decoder_bit_T_365=_id_ctrl_decoder_bit_T_364|_id_ctrl_decoder_bit_T_97; 
  assign _id_ctrl_decoder_bit_T_366=_id_ctrl_decoder_bit_T_365|_id_ctrl_decoder_bit_T_99; 
  assign _id_ctrl_decoder_bit_T_367=_id_ctrl_decoder_bit_T_366|_id_ctrl_decoder_bit_T_101; 
  assign _id_ctrl_decoder_bit_T_368=_id_ctrl_decoder_bit_T_367|_id_ctrl_decoder_bit_T_103; 
  assign _id_ctrl_decoder_bit_T_369=_id_ctrl_decoder_bit_T_368|_id_ctrl_decoder_bit_T_105; 
  assign _id_ctrl_decoder_bit_T_370=_id_ctrl_decoder_bit_T_369|_id_ctrl_decoder_bit_T_107; 
  assign _id_ctrl_decoder_bit_T_371=_id_ctrl_decoder_bit_T_370|_id_ctrl_decoder_bit_T_109; 
  assign _id_ctrl_decoder_bit_T_372=_id_ctrl_decoder_bit_T_371|_id_ctrl_decoder_bit_T_111; 
  assign _id_ctrl_decoder_bit_T_373=_id_ctrl_decoder_bit_T_372|_id_ctrl_decoder_bit_T_113; 
  assign _id_ctrl_decoder_bit_T_374=_id_ctrl_decoder_bit_T_373|_id_ctrl_decoder_bit_T_115; 
  assign _id_ctrl_decoder_bit_T_375=_id_ctrl_decoder_bit_T_374|_id_ctrl_decoder_bit_T_117; 
  assign _id_ctrl_decoder_bit_T_376=_id_ctrl_decoder_bit_T_375|_id_ctrl_decoder_bit_T_119; 
  assign _id_ctrl_decoder_bit_T_377=_id_ctrl_decoder_bit_T_376|_id_ctrl_decoder_bit_T_121; 
  assign _id_ctrl_decoder_bit_T_378=_id_ctrl_decoder_bit_T_377|_id_ctrl_decoder_bit_T_123; 
  assign _id_ctrl_decoder_bit_T_379=_id_ctrl_decoder_bit_T_378|_id_ctrl_decoder_bit_T_125; 
  assign _id_ctrl_decoder_bit_T_380=_id_ctrl_decoder_bit_T_379|_id_ctrl_decoder_bit_T_127; 
  assign _id_ctrl_decoder_bit_T_381=_id_ctrl_decoder_bit_T_380|_id_ctrl_decoder_bit_T_129; 
  assign _id_ctrl_decoder_bit_T_382=_id_ctrl_decoder_bit_T_381|_id_ctrl_decoder_bit_T_131; 
  assign _id_ctrl_decoder_bit_T_383=_id_ctrl_decoder_bit_T_382|_id_ctrl_decoder_bit_T_133; 
  assign _id_ctrl_decoder_bit_T_384=_id_ctrl_decoder_bit_T_383|_id_ctrl_decoder_bit_T_135; 
  assign _id_ctrl_decoder_bit_T_385=_id_ctrl_decoder_bit_T_384|_id_ctrl_decoder_bit_T_137; 
  assign _id_ctrl_decoder_bit_T_386=_id_ctrl_decoder_bit_T_385|_id_ctrl_decoder_bit_T_139; 
  assign _id_ctrl_decoder_bit_T_387=_id_ctrl_decoder_bit_T_386|_id_ctrl_decoder_bit_T_141; 
  assign _id_ctrl_decoder_bit_T_388=_id_ctrl_decoder_bit_T_387|_id_ctrl_decoder_bit_T_143; 
  assign _id_ctrl_decoder_bit_T_389=_id_ctrl_decoder_bit_T_388|_id_ctrl_decoder_bit_T_145; 
  assign _id_ctrl_decoder_bit_T_390=_id_ctrl_decoder_bit_T_389|_id_ctrl_decoder_bit_T_147; 
  assign _id_ctrl_decoder_bit_T_391=_id_ctrl_decoder_bit_T_390|_id_ctrl_decoder_bit_T_149; 
  assign _id_ctrl_decoder_bit_T_392=_id_ctrl_decoder_bit_T_391|_id_ctrl_decoder_bit_T_151; 
  assign _id_ctrl_decoder_bit_T_393=_id_ctrl_decoder_bit_T_392|_id_ctrl_decoder_bit_T_153; 
  assign _id_ctrl_decoder_bit_T_394=_id_ctrl_decoder_bit_T_393|_id_ctrl_decoder_bit_T_155; 
  assign _id_ctrl_decoder_bit_T_395=_id_ctrl_decoder_bit_T_394|_id_ctrl_decoder_bit_T_157; 
  assign _id_ctrl_decoder_bit_T_396=_id_ctrl_decoder_bit_T_395|_id_ctrl_decoder_bit_T_159; 
  assign _id_ctrl_decoder_bit_T_397=_id_ctrl_decoder_bit_T_396|_id_ctrl_decoder_bit_T_161; 
  assign _id_ctrl_decoder_bit_T_398=_id_ctrl_decoder_bit_T_397|_id_ctrl_decoder_bit_T_163; 
  assign _id_ctrl_decoder_bit_T_399=_id_ctrl_decoder_bit_T_398|_id_ctrl_decoder_bit_T_165; 
  assign _id_ctrl_decoder_bit_T_400=_id_ctrl_decoder_bit_T_399|_id_ctrl_decoder_bit_T_167; 
  assign _id_ctrl_decoder_bit_T_401=_id_ctrl_decoder_bit_T_400|_id_ctrl_decoder_bit_T_169; 
  assign _id_ctrl_decoder_bit_T_402=_id_ctrl_decoder_bit_T_401|_id_ctrl_decoder_bit_T_171; 
  assign _id_ctrl_decoder_bit_T_403=_id_ctrl_decoder_bit_T_402|_id_ctrl_decoder_bit_T_173; 
  assign _id_ctrl_decoder_bit_T_404=_id_ctrl_decoder_bit_T_403|_id_ctrl_decoder_bit_T_175; 
  assign _id_ctrl_decoder_bit_T_405=_id_ctrl_decoder_bit_T_404|_id_ctrl_decoder_bit_T_177; 
  assign _id_ctrl_decoder_bit_T_406=_id_ctrl_decoder_bit_T_405|_id_ctrl_decoder_bit_T_179; 
  assign _id_ctrl_decoder_bit_T_407=_id_ctrl_decoder_bit_T_406|_id_ctrl_decoder_bit_T_181; 
  assign _id_ctrl_decoder_bit_T_408=_id_ctrl_decoder_bit_T_407|_id_ctrl_decoder_bit_T_183; 
  assign _id_ctrl_decoder_bit_T_409=_id_ctrl_decoder_bit_T_408|_id_ctrl_decoder_bit_T_185; 
  assign _id_ctrl_decoder_bit_T_410=_id_ctrl_decoder_bit_T_409|_id_ctrl_decoder_bit_T_187; 
  assign _id_ctrl_decoder_bit_T_411=_id_ctrl_decoder_bit_T_410|_id_ctrl_decoder_bit_T_189; 
  assign _id_ctrl_decoder_bit_T_412=_id_ctrl_decoder_bit_T_411|_id_ctrl_decoder_bit_T_191; 
  assign _id_ctrl_decoder_bit_T_413=_id_ctrl_decoder_bit_T_412|_id_ctrl_decoder_bit_T_193; 
  assign _id_ctrl_decoder_bit_T_414=_id_ctrl_decoder_bit_T_413|_id_ctrl_decoder_bit_T_195; 
  assign _id_ctrl_decoder_bit_T_415=_id_ctrl_decoder_bit_T_414|_id_ctrl_decoder_bit_T_197; 
  assign _id_ctrl_decoder_bit_T_416=_id_ctrl_decoder_bit_T_415|_id_ctrl_decoder_bit_T_199; 
  assign _id_ctrl_decoder_bit_T_417=_id_ctrl_decoder_bit_T_416|_id_ctrl_decoder_bit_T_201; 
  assign _id_ctrl_decoder_bit_T_418=_id_ctrl_decoder_bit_T_417|_id_ctrl_decoder_bit_T_203; 
  assign _id_ctrl_decoder_bit_T_419=_id_ctrl_decoder_bit_T_418|_id_ctrl_decoder_bit_T_205; 
  assign _id_ctrl_decoder_bit_T_420=_id_ctrl_decoder_bit_T_419|_id_ctrl_decoder_bit_T_207; 
  assign _id_ctrl_decoder_bit_T_421=_id_ctrl_decoder_bit_T_420|_id_ctrl_decoder_bit_T_209; 
  assign _id_ctrl_decoder_bit_T_422=_id_ctrl_decoder_bit_T_421|_id_ctrl_decoder_bit_T_211; 
  assign _id_ctrl_decoder_bit_T_423=_id_ctrl_decoder_bit_T_422|_id_ctrl_decoder_bit_T_213; 
  assign _id_ctrl_decoder_bit_T_424=_id_ctrl_decoder_bit_T_423|_id_ctrl_decoder_bit_T_215; 
  assign _id_ctrl_decoder_bit_T_425=_id_ctrl_decoder_bit_T_424|_id_ctrl_decoder_bit_T_217; 
  assign _id_ctrl_decoder_bit_T_426=_id_ctrl_decoder_bit_T_425|_id_ctrl_decoder_bit_T_219; 
  assign _id_ctrl_decoder_bit_T_427=_id_ctrl_decoder_bit_T_426|_id_ctrl_decoder_bit_T_221; 
  assign _id_ctrl_decoder_bit_T_428=_id_ctrl_decoder_bit_T_427|_id_ctrl_decoder_bit_T_223; 
  assign _id_ctrl_decoder_bit_T_429=_id_ctrl_decoder_bit_T_428|_id_ctrl_decoder_bit_T_225; 
  assign _id_ctrl_decoder_bit_T_430=_id_ctrl_decoder_bit_T_429|_id_ctrl_decoder_bit_T_226; 
  assign _id_ctrl_decoder_bit_T_431=_id_ctrl_decoder_bit_T_430|_id_ctrl_decoder_bit_T_227; 
  assign _id_ctrl_decoder_bit_T_432=_id_ctrl_decoder_bit_T_431|_id_ctrl_decoder_bit_T_229; 
  assign _id_ctrl_decoder_bit_T_433=_id_ctrl_decoder_bit_T_432|_id_ctrl_decoder_bit_T_231; 
  assign _id_ctrl_decoder_bit_T_434=_id_ctrl_decoder_bit_T_433|_id_ctrl_decoder_bit_T_233; 
  assign _id_ctrl_decoder_bit_T_435=_id_ctrl_decoder_bit_T_434|_id_ctrl_decoder_bit_T_235; 
  assign _id_ctrl_decoder_bit_T_436=_id_ctrl_decoder_bit_T_435|_id_ctrl_decoder_bit_T_237; 
  assign _id_ctrl_decoder_bit_T_437=_id_ctrl_decoder_bit_T_436|_id_ctrl_decoder_bit_T_239; 
  assign _id_ctrl_decoder_bit_T_438=_id_ctrl_decoder_bit_T_437|_id_ctrl_decoder_bit_T_241; 
  assign _id_ctrl_decoder_bit_T_439=_id_ctrl_decoder_bit_T_438|_id_ctrl_decoder_bit_T_243; 
  assign _id_ctrl_decoder_bit_T_440=_id_ctrl_decoder_bit_T_439|_id_ctrl_decoder_bit_T_245; 
  assign _id_ctrl_decoder_bit_T_441=_id_ctrl_decoder_bit_T_440|_id_ctrl_decoder_bit_T_247; 
  assign _id_ctrl_decoder_bit_T_442=_id_ctrl_decoder_bit_T_441|_id_ctrl_decoder_bit_T_249; 
  assign _id_ctrl_decoder_bit_T_443=_id_ctrl_decoder_bit_T_442|_id_ctrl_decoder_bit_T_251; 
  assign _id_ctrl_decoder_bit_T_444=_id_ctrl_decoder_bit_T_443|_id_ctrl_decoder_bit_T_253; 
  assign _id_ctrl_decoder_bit_T_445=_id_ctrl_decoder_bit_T_444|_id_ctrl_decoder_bit_T_255; 
  assign _id_ctrl_decoder_bit_T_446=_id_ctrl_decoder_bit_T_445|_id_ctrl_decoder_bit_T_257; 
  assign _id_ctrl_decoder_bit_T_447=_id_ctrl_decoder_bit_T_446|_id_ctrl_decoder_bit_T_259; 
  assign _id_ctrl_decoder_bit_T_448=_id_ctrl_decoder_bit_T_447|_id_ctrl_decoder_bit_T_261; 
  assign _id_ctrl_decoder_bit_T_449=_id_ctrl_decoder_bit_T_448|_id_ctrl_decoder_bit_T_263; 
  assign _id_ctrl_decoder_bit_T_450=_id_ctrl_decoder_bit_T_449|_id_ctrl_decoder_bit_T_265; 
  assign _id_ctrl_decoder_bit_T_451=_id_ctrl_decoder_bit_T_450|_id_ctrl_decoder_bit_T_267; 
  assign _id_ctrl_decoder_bit_T_452=_id_ctrl_decoder_bit_T_451|_id_ctrl_decoder_bit_T_269; 
  assign _id_ctrl_decoder_bit_T_453=_id_ctrl_decoder_bit_T_452|_id_ctrl_decoder_bit_T_271; 
  assign _id_ctrl_decoder_bit_T_454=_id_ctrl_decoder_bit_T_453|_id_ctrl_decoder_bit_T_273; 
  assign _id_ctrl_decoder_bit_T_455=_id_ctrl_decoder_bit_T_454|_id_ctrl_decoder_bit_T_275; 
  assign _id_ctrl_decoder_bit_T_456=_id_ctrl_decoder_bit_T_455|_id_ctrl_decoder_bit_T_277; 
  assign _id_ctrl_decoder_bit_T_457=_id_ctrl_decoder_bit_T_456|_id_ctrl_decoder_bit_T_279; 
  assign _id_ctrl_decoder_bit_T_458=_id_ctrl_decoder_bit_T_457|_id_ctrl_decoder_bit_T_281; 
  assign _id_ctrl_decoder_bit_T_459=_id_ctrl_decoder_bit_T_458|_id_ctrl_decoder_bit_T_283; 
  assign _id_ctrl_decoder_bit_T_460=_id_ctrl_decoder_bit_T_459|_id_ctrl_decoder_bit_T_285; 
  assign _id_ctrl_decoder_bit_T_461=_id_ctrl_decoder_bit_T_460|_id_ctrl_decoder_bit_T_287; 
  assign _id_ctrl_decoder_bit_T_462=_id_ctrl_decoder_bit_T_461|_id_ctrl_decoder_bit_T_289; 
  assign _id_ctrl_decoder_bit_T_463=_id_ctrl_decoder_bit_T_462|_id_ctrl_decoder_bit_T_291; 
  assign _id_ctrl_decoder_bit_T_464=_id_ctrl_decoder_bit_T_463|_id_ctrl_decoder_bit_T_293; 
  assign _id_ctrl_decoder_bit_T_465=_id_ctrl_decoder_bit_T_464|_id_ctrl_decoder_bit_T_295; 
  assign _id_ctrl_decoder_bit_T_466=_id_ctrl_decoder_bit_T_465|_id_ctrl_decoder_bit_T_297; 
  assign _id_ctrl_decoder_bit_T_467=_id_ctrl_decoder_bit_T_466|_id_ctrl_decoder_bit_T_299; 
  assign _id_ctrl_decoder_bit_T_468=_id_ctrl_decoder_bit_T_467|_id_ctrl_decoder_bit_T_300; 
  assign _id_ctrl_decoder_bit_T_469=_id_ctrl_decoder_bit_T_468|_id_ctrl_decoder_bit_T_301; 
  assign _id_ctrl_decoder_bit_T_470=_id_ctrl_decoder_bit_T_469|_id_ctrl_decoder_bit_T_302; 
  assign _id_ctrl_decoder_bit_T_471=_id_ctrl_decoder_bit_T_470|_id_ctrl_decoder_bit_T_303; 
  assign _id_ctrl_decoder_bit_T_472=_id_ctrl_decoder_bit_T_471|_id_ctrl_decoder_bit_T_304; 
  assign _id_ctrl_decoder_bit_T_473=_id_ctrl_decoder_bit_T_472|_id_ctrl_decoder_bit_T_306; 
  assign _id_ctrl_decoder_bit_T_474=_id_ctrl_decoder_bit_T_473|_id_ctrl_decoder_bit_T_308; 
  assign _id_ctrl_decoder_bit_T_475=_id_ctrl_decoder_bit_T_474|_id_ctrl_decoder_bit_T_310; 
  assign _id_ctrl_decoder_bit_T_476=_id_ctrl_decoder_bit_T_475|_id_ctrl_decoder_bit_T_312; 
  assign _id_ctrl_decoder_bit_T_477=_id_ctrl_decoder_bit_T_476|_id_ctrl_decoder_bit_T_314; 
  assign id_ctrl_decoder_0=_id_ctrl_decoder_bit_T_477|_id_ctrl_decoder_bit_T_316; 
  assign _id_ctrl_decoder_T=ibuf_io_inst_0_bits_inst_bits&32'h5c; 
  assign _id_ctrl_decoder_T_1=_id_ctrl_decoder_T==32'h4; 
  assign _id_ctrl_decoder_T_2=ibuf_io_inst_0_bits_inst_bits&32'h60; 
  assign _id_ctrl_decoder_T_3=_id_ctrl_decoder_T_2==32'h40; 
  assign id_ctrl_decoder_1=_id_ctrl_decoder_T_1|_id_ctrl_decoder_T_3; 
  assign _id_ctrl_decoder_T_5=ibuf_io_inst_0_bits_inst_bits&32'h74; 
  assign id_ctrl_decoder_3=_id_ctrl_decoder_T_5==32'h60; 
  assign _id_ctrl_decoder_T_7=ibuf_io_inst_0_bits_inst_bits&32'h68; 
  assign id_ctrl_decoder_4=_id_ctrl_decoder_T_7==32'h68; 
  assign _id_ctrl_decoder_T_9=ibuf_io_inst_0_bits_inst_bits&32'h203c; 
  assign id_ctrl_decoder_5=_id_ctrl_decoder_T_9==32'h24; 
  assign _id_ctrl_decoder_T_11=ibuf_io_inst_0_bits_inst_bits&32'h64; 
  assign _id_ctrl_decoder_T_12=_id_ctrl_decoder_T_11==32'h20; 
  assign _id_ctrl_decoder_T_13=ibuf_io_inst_0_bits_inst_bits&32'h34; 
  assign _id_ctrl_decoder_T_14=_id_ctrl_decoder_T_13==32'h20; 
  assign _id_ctrl_decoder_T_15=ibuf_io_inst_0_bits_inst_bits&32'h2048; 
  assign _id_ctrl_decoder_T_16=_id_ctrl_decoder_T_15==32'h2008; 
  assign _id_ctrl_decoder_T_17=ibuf_io_inst_0_bits_inst_bits&32'h42003024; 
  assign _id_ctrl_decoder_T_18=_id_ctrl_decoder_T_17==32'h2000020; 
  assign _id_ctrl_decoder_T_20=_id_ctrl_decoder_T_12|_id_ctrl_decoder_T_14; 
  assign _id_ctrl_decoder_T_21=_id_ctrl_decoder_T_20|_id_ctrl_decoder_T_16; 
  assign id_ctrl_decoder_6=_id_ctrl_decoder_T_21|_id_ctrl_decoder_T_18; 
  assign _id_ctrl_decoder_T_22=ibuf_io_inst_0_bits_inst_bits&32'h44; 
  assign _id_ctrl_decoder_T_23=_id_ctrl_decoder_T_22==32'h0; 
  assign _id_ctrl_decoder_T_24=ibuf_io_inst_0_bits_inst_bits&32'h4024; 
  assign _id_ctrl_decoder_T_25=_id_ctrl_decoder_T_24==32'h20; 
  assign _id_ctrl_decoder_T_26=ibuf_io_inst_0_bits_inst_bits&32'h38; 
  assign _id_ctrl_decoder_T_27=_id_ctrl_decoder_T_26==32'h20; 
  assign _id_ctrl_decoder_T_28=ibuf_io_inst_0_bits_inst_bits&32'h2050; 
  assign _id_ctrl_decoder_T_29=_id_ctrl_decoder_T_28==32'h2000; 
  assign _id_ctrl_decoder_T_30=ibuf_io_inst_0_bits_inst_bits&32'h90000034; 
  assign _id_ctrl_decoder_T_31=_id_ctrl_decoder_T_30==32'h90000010; 
  assign _id_ctrl_decoder_T_33=_id_ctrl_decoder_T_23|_id_ctrl_decoder_T_25; 
  assign _id_ctrl_decoder_T_34=_id_ctrl_decoder_T_33|_id_ctrl_decoder_T_27; 
  assign _id_ctrl_decoder_T_35=_id_ctrl_decoder_T_34|_id_ctrl_decoder_T_29; 
  assign id_ctrl_decoder_7=_id_ctrl_decoder_T_35|_id_ctrl_decoder_T_31; 
  assign _id_ctrl_decoder_T_36=ibuf_io_inst_0_bits_inst_bits&32'h58; 
  assign _id_ctrl_decoder_T_37=_id_ctrl_decoder_T_36==32'h0; 
  assign _id_ctrl_decoder_T_38=ibuf_io_inst_0_bits_inst_bits&32'h20; 
  assign _id_ctrl_decoder_T_39=_id_ctrl_decoder_T_38==32'h0; 
  assign _id_ctrl_decoder_T_40=ibuf_io_inst_0_bits_inst_bits&32'hc; 
  assign _id_ctrl_decoder_T_41=_id_ctrl_decoder_T_40==32'h4; 
  assign _id_ctrl_decoder_T_42=ibuf_io_inst_0_bits_inst_bits&32'h48; 
  assign _id_ctrl_decoder_T_43=_id_ctrl_decoder_T_42==32'h48; 
  assign _id_ctrl_decoder_T_44=ibuf_io_inst_0_bits_inst_bits&32'h4050; 
  assign _id_ctrl_decoder_T_45=_id_ctrl_decoder_T_44==32'h4050; 
  assign _id_ctrl_decoder_T_47=_id_ctrl_decoder_T_37|_id_ctrl_decoder_T_39; 
  assign _id_ctrl_decoder_T_48=_id_ctrl_decoder_T_47|_id_ctrl_decoder_T_41; 
  assign _id_ctrl_decoder_T_49=_id_ctrl_decoder_T_48|_id_ctrl_decoder_T_43; 
  assign id_ctrl_decoder_lo=_id_ctrl_decoder_T_49|_id_ctrl_decoder_T_45; 
  assign _id_ctrl_decoder_T_51=_id_ctrl_decoder_T_42==32'h0; 
  assign _id_ctrl_decoder_T_52=ibuf_io_inst_0_bits_inst_bits&32'h18; 
  assign _id_ctrl_decoder_T_53=_id_ctrl_decoder_T_52==32'h0; 
  assign _id_ctrl_decoder_T_54=ibuf_io_inst_0_bits_inst_bits&32'h4008; 
  assign _id_ctrl_decoder_T_55=_id_ctrl_decoder_T_54==32'h4000; 
  assign _id_ctrl_decoder_T_57=_id_ctrl_decoder_T_51|_id_ctrl_decoder_T_23; 
  assign _id_ctrl_decoder_T_58=_id_ctrl_decoder_T_57|_id_ctrl_decoder_T_53; 
  assign id_ctrl_decoder_hi=_id_ctrl_decoder_T_58|_id_ctrl_decoder_T_55; 
  assign id_ctrl_decoder_9={id_ctrl_decoder_hi,id_ctrl_decoder_lo}; 
  assign _id_ctrl_decoder_T_59=ibuf_io_inst_0_bits_inst_bits&32'h4004; 
  assign _id_ctrl_decoder_T_60=_id_ctrl_decoder_T_59==32'h0; 
  assign _id_ctrl_decoder_T_61=ibuf_io_inst_0_bits_inst_bits&32'h50; 
  assign _id_ctrl_decoder_T_62=_id_ctrl_decoder_T_61==32'h0; 
  assign _id_ctrl_decoder_T_63=ibuf_io_inst_0_bits_inst_bits&32'h24; 
  assign _id_ctrl_decoder_T_64=_id_ctrl_decoder_T_63==32'h0; 
  assign _id_ctrl_decoder_T_66=_id_ctrl_decoder_T_60|_id_ctrl_decoder_T_62; 
  assign _id_ctrl_decoder_T_67=_id_ctrl_decoder_T_66|_id_ctrl_decoder_T_23; 
  assign _id_ctrl_decoder_T_68=_id_ctrl_decoder_T_67|_id_ctrl_decoder_T_64; 
  assign id_ctrl_decoder_lo_1=_id_ctrl_decoder_T_68|_id_ctrl_decoder_T_53; 
  assign _id_ctrl_decoder_T_70=_id_ctrl_decoder_T_13==32'h14; 
  assign id_ctrl_decoder_hi_1=_id_ctrl_decoder_T_70|_id_ctrl_decoder_T_43; 
  assign id_ctrl_decoder_10={id_ctrl_decoder_hi_1,id_ctrl_decoder_lo_1}; 
  assign _id_ctrl_decoder_T_73=_id_ctrl_decoder_T_52==32'h8; 
  assign _id_ctrl_decoder_T_75=_id_ctrl_decoder_T_22==32'h40; 
  assign id_ctrl_decoder_lo_2=_id_ctrl_decoder_T_73|_id_ctrl_decoder_T_75; 
  assign _id_ctrl_decoder_T_77=ibuf_io_inst_0_bits_inst_bits&32'h14; 
  assign _id_ctrl_decoder_T_78=_id_ctrl_decoder_T_77==32'h14; 
  assign id_ctrl_decoder_hi_lo=_id_ctrl_decoder_T_73|_id_ctrl_decoder_T_78; 
  assign _id_ctrl_decoder_T_80=ibuf_io_inst_0_bits_inst_bits&32'h30; 
  assign _id_ctrl_decoder_T_81=_id_ctrl_decoder_T_80==32'h0; 
  assign _id_ctrl_decoder_T_82=ibuf_io_inst_0_bits_inst_bits&32'h201c; 
  assign _id_ctrl_decoder_T_83=_id_ctrl_decoder_T_82==32'h4; 
  assign _id_ctrl_decoder_T_85=_id_ctrl_decoder_T_77==32'h10; 
  assign _id_ctrl_decoder_T_87=_id_ctrl_decoder_T_81|_id_ctrl_decoder_T_83; 
  assign id_ctrl_decoder_hi_hi=_id_ctrl_decoder_T_87|_id_ctrl_decoder_T_85; 
  assign id_ctrl_decoder_11={id_ctrl_decoder_hi_hi,id_ctrl_decoder_hi_lo,id_ctrl_decoder_lo_2}; 
  assign _id_ctrl_decoder_T_88=ibuf_io_inst_0_bits_inst_bits&32'h10; 
  assign _id_ctrl_decoder_T_89=_id_ctrl_decoder_T_88==32'h0; 
  assign _id_ctrl_decoder_T_90=ibuf_io_inst_0_bits_inst_bits&32'h8; 
  assign _id_ctrl_decoder_T_91=_id_ctrl_decoder_T_90==32'h0; 
  assign id_ctrl_decoder_12=_id_ctrl_decoder_T_89|_id_ctrl_decoder_T_91; 
  assign _id_ctrl_decoder_T_93=ibuf_io_inst_0_bits_inst_bits&32'h3054; 
  assign _id_ctrl_decoder_T_94=_id_ctrl_decoder_T_93==32'h1010; 
  assign _id_ctrl_decoder_T_95=ibuf_io_inst_0_bits_inst_bits&32'h1058; 
  assign _id_ctrl_decoder_T_96=_id_ctrl_decoder_T_95==32'h1040; 
  assign _id_ctrl_decoder_T_97=ibuf_io_inst_0_bits_inst_bits&32'h7044; 
  assign _id_ctrl_decoder_T_98=_id_ctrl_decoder_T_97==32'h7000; 
  assign _id_ctrl_decoder_T_99=ibuf_io_inst_0_bits_inst_bits&32'h2001074; 
  assign _id_ctrl_decoder_T_100=_id_ctrl_decoder_T_99==32'h2001030; 
  assign _id_ctrl_decoder_T_102=_id_ctrl_decoder_T_94|_id_ctrl_decoder_T_96; 
  assign _id_ctrl_decoder_T_103=_id_ctrl_decoder_T_102|_id_ctrl_decoder_T_98; 
  assign id_ctrl_decoder_lo_lo=_id_ctrl_decoder_T_103|_id_ctrl_decoder_T_100; 
  assign _id_ctrl_decoder_T_104=ibuf_io_inst_0_bits_inst_bits&32'h4054; 
  assign _id_ctrl_decoder_T_105=_id_ctrl_decoder_T_104==32'h40; 
  assign _id_ctrl_decoder_T_106=ibuf_io_inst_0_bits_inst_bits&32'h2058; 
  assign _id_ctrl_decoder_T_107=_id_ctrl_decoder_T_106==32'h2040; 
  assign _id_ctrl_decoder_T_109=_id_ctrl_decoder_T_93==32'h3010; 
  assign _id_ctrl_decoder_T_110=ibuf_io_inst_0_bits_inst_bits&32'h6054; 
  assign _id_ctrl_decoder_T_111=_id_ctrl_decoder_T_110==32'h6010; 
  assign _id_ctrl_decoder_T_112=ibuf_io_inst_0_bits_inst_bits&32'h2002074; 
  assign _id_ctrl_decoder_T_113=_id_ctrl_decoder_T_112==32'h2002030; 
  assign _id_ctrl_decoder_T_114=ibuf_io_inst_0_bits_inst_bits&32'h40003034; 
  assign _id_ctrl_decoder_T_115=_id_ctrl_decoder_T_114==32'h40000030; 
  assign _id_ctrl_decoder_T_116=ibuf_io_inst_0_bits_inst_bits&32'h40001054; 
  assign _id_ctrl_decoder_T_117=_id_ctrl_decoder_T_116==32'h40001010; 
  assign _id_ctrl_decoder_T_119=_id_ctrl_decoder_T_105|_id_ctrl_decoder_T_107; 
  assign _id_ctrl_decoder_T_120=_id_ctrl_decoder_T_119|_id_ctrl_decoder_T_109; 
  assign _id_ctrl_decoder_T_121=_id_ctrl_decoder_T_120|_id_ctrl_decoder_T_111; 
  assign _id_ctrl_decoder_T_122=_id_ctrl_decoder_T_121|_id_ctrl_decoder_T_113; 
  assign _id_ctrl_decoder_T_123=_id_ctrl_decoder_T_122|_id_ctrl_decoder_T_115; 
  assign id_ctrl_decoder_lo_hi=_id_ctrl_decoder_T_123|_id_ctrl_decoder_T_117; 
  assign _id_ctrl_decoder_T_124=ibuf_io_inst_0_bits_inst_bits&32'h2002054; 
  assign _id_ctrl_decoder_T_125=_id_ctrl_decoder_T_124==32'h2010; 
  assign _id_ctrl_decoder_T_126=ibuf_io_inst_0_bits_inst_bits&32'h2034; 
  assign _id_ctrl_decoder_T_127=_id_ctrl_decoder_T_126==32'h2010; 
  assign _id_ctrl_decoder_T_128=ibuf_io_inst_0_bits_inst_bits&32'h40004054; 
  assign _id_ctrl_decoder_T_129=_id_ctrl_decoder_T_128==32'h4010; 
  assign _id_ctrl_decoder_T_130=ibuf_io_inst_0_bits_inst_bits&32'h5054; 
  assign _id_ctrl_decoder_T_131=_id_ctrl_decoder_T_130==32'h4010; 
  assign _id_ctrl_decoder_T_132=ibuf_io_inst_0_bits_inst_bits&32'h4058; 
  assign _id_ctrl_decoder_T_133=_id_ctrl_decoder_T_132==32'h4040; 
  assign _id_ctrl_decoder_T_135=_id_ctrl_decoder_T_125|_id_ctrl_decoder_T_127; 
  assign _id_ctrl_decoder_T_136=_id_ctrl_decoder_T_135|_id_ctrl_decoder_T_129; 
  assign _id_ctrl_decoder_T_137=_id_ctrl_decoder_T_136|_id_ctrl_decoder_T_131; 
  assign id_ctrl_decoder_hi_lo_1=_id_ctrl_decoder_T_137|_id_ctrl_decoder_T_133; 
  assign _id_ctrl_decoder_T_138=ibuf_io_inst_0_bits_inst_bits&32'h2006054; 
  assign _id_ctrl_decoder_T_139=_id_ctrl_decoder_T_138==32'h2010; 
  assign _id_ctrl_decoder_T_140=ibuf_io_inst_0_bits_inst_bits&32'h6034; 
  assign _id_ctrl_decoder_T_141=_id_ctrl_decoder_T_140==32'h2010; 
  assign _id_ctrl_decoder_T_142=ibuf_io_inst_0_bits_inst_bits&32'h40003054; 
  assign _id_ctrl_decoder_T_143=_id_ctrl_decoder_T_142==32'h40001010; 
  assign _id_ctrl_decoder_T_145=_id_ctrl_decoder_T_139|_id_ctrl_decoder_T_141; 
  assign _id_ctrl_decoder_T_146=_id_ctrl_decoder_T_145|_id_ctrl_decoder_T_133; 
  assign _id_ctrl_decoder_T_147=_id_ctrl_decoder_T_146|_id_ctrl_decoder_T_115; 
  assign id_ctrl_decoder_hi_hi_1=_id_ctrl_decoder_T_147|_id_ctrl_decoder_T_143; 
  assign id_ctrl_decoder_13={id_ctrl_decoder_hi_hi_1,id_ctrl_decoder_hi_lo_1,id_ctrl_decoder_lo_hi,id_ctrl_decoder_lo_lo}; 
  assign _id_ctrl_decoder_bit_T_479=_id_ctrl_decoder_bit_T_27|_id_ctrl_decoder_bit_T_29; 
  assign _id_ctrl_decoder_bit_T_480=_id_ctrl_decoder_bit_T_479|_id_ctrl_decoder_bit_T_31; 
  assign _id_ctrl_decoder_bit_T_481=_id_ctrl_decoder_bit_T_480|_id_ctrl_decoder_bit_T_33; 
  assign _id_ctrl_decoder_bit_T_482=_id_ctrl_decoder_bit_T_481|_id_ctrl_decoder_bit_T_35; 
  assign _id_ctrl_decoder_bit_T_483=_id_ctrl_decoder_bit_T_482|_id_ctrl_decoder_bit_T_37; 
  assign _id_ctrl_decoder_bit_T_484=_id_ctrl_decoder_bit_T_483|_id_ctrl_decoder_bit_T_39; 
  assign _id_ctrl_decoder_bit_T_485=_id_ctrl_decoder_bit_T_484|_id_ctrl_decoder_bit_T_41; 
  assign _id_ctrl_decoder_bit_T_486=_id_ctrl_decoder_bit_T_485|_id_ctrl_decoder_bit_T_43; 
  assign _id_ctrl_decoder_bit_T_487=_id_ctrl_decoder_bit_T_486|_id_ctrl_decoder_bit_T_45; 
  assign _id_ctrl_decoder_bit_T_488=_id_ctrl_decoder_bit_T_487|_id_ctrl_decoder_bit_T_47; 
  assign _id_ctrl_decoder_bit_T_489=_id_ctrl_decoder_bit_T_488|_id_ctrl_decoder_bit_T_49; 
  assign _id_ctrl_decoder_bit_T_490=_id_ctrl_decoder_bit_T_489|_id_ctrl_decoder_bit_T_51; 
  assign _id_ctrl_decoder_bit_T_491=_id_ctrl_decoder_bit_T_490|_id_ctrl_decoder_bit_T_53; 
  assign _id_ctrl_decoder_bit_T_492=_id_ctrl_decoder_bit_T_491|_id_ctrl_decoder_bit_T_55; 
  assign _id_ctrl_decoder_bit_T_493=_id_ctrl_decoder_bit_T_492|_id_ctrl_decoder_bit_T_57; 
  assign _id_ctrl_decoder_bit_T_494=_id_ctrl_decoder_bit_T_493|_id_ctrl_decoder_bit_T_59; 
  assign _id_ctrl_decoder_bit_T_495=_id_ctrl_decoder_bit_T_494|_id_ctrl_decoder_bit_T_61; 
  assign _id_ctrl_decoder_bit_T_496=_id_ctrl_decoder_bit_T_495|_id_ctrl_decoder_bit_T_63; 
  assign _id_ctrl_decoder_bit_T_497=_id_ctrl_decoder_bit_T_496|_id_ctrl_decoder_bit_T_65; 
  assign _id_ctrl_decoder_bit_T_498=_id_ctrl_decoder_bit_T_497|_id_ctrl_decoder_bit_T_67; 
  assign _id_ctrl_decoder_bit_T_499=_id_ctrl_decoder_bit_T_498|_id_ctrl_decoder_bit_T_69; 
  assign _id_ctrl_decoder_bit_T_500=_id_ctrl_decoder_bit_T_499|_id_ctrl_decoder_bit_T_115; 
  assign _id_ctrl_decoder_bit_T_501=_id_ctrl_decoder_bit_T_500|_id_ctrl_decoder_bit_T_117; 
  assign _id_ctrl_decoder_bit_T_502=_id_ctrl_decoder_bit_T_501|_id_ctrl_decoder_bit_T_175; 
  assign _id_ctrl_decoder_bit_T_503=_id_ctrl_decoder_bit_T_502|_id_ctrl_decoder_bit_T_177; 
  assign _id_ctrl_decoder_bit_T_504=_id_ctrl_decoder_bit_T_503|_id_ctrl_decoder_bit_T_195; 
  assign _id_ctrl_decoder_bit_T_505=_id_ctrl_decoder_bit_T_504|_id_ctrl_decoder_bit_T_197; 
  assign _id_ctrl_decoder_bit_T_506=_id_ctrl_decoder_bit_T_505|_id_ctrl_decoder_bit_T_199; 
  assign _id_ctrl_decoder_bit_T_507=_id_ctrl_decoder_bit_T_506|_id_ctrl_decoder_bit_T_225; 
  assign _id_ctrl_decoder_bit_T_508=_id_ctrl_decoder_bit_T_507|_id_ctrl_decoder_bit_T_249; 
  assign _id_ctrl_decoder_bit_T_509=_id_ctrl_decoder_bit_T_508|_id_ctrl_decoder_bit_T_251; 
  assign _id_ctrl_decoder_bit_T_510=_id_ctrl_decoder_bit_T_509|_id_ctrl_decoder_bit_T_253; 
  assign _id_ctrl_decoder_bit_T_511=_id_ctrl_decoder_bit_T_510|_id_ctrl_decoder_bit_T_255; 
  assign _id_ctrl_decoder_bit_T_512=_id_ctrl_decoder_bit_T_511|_id_ctrl_decoder_bit_T_257; 
  assign _id_ctrl_decoder_bit_T_513=_id_ctrl_decoder_bit_T_512|_id_ctrl_decoder_bit_T_259; 
  assign _id_ctrl_decoder_bit_T_514=_id_ctrl_decoder_bit_T_513|_id_ctrl_decoder_bit_T_261; 
  assign id_ctrl_decoder_14=_id_ctrl_decoder_bit_T_514|_id_ctrl_decoder_bit_T_263; 
  assign _id_ctrl_decoder_T_149=_id_ctrl_decoder_T_7==32'h20; 
  assign _id_ctrl_decoder_T_150=ibuf_io_inst_0_bits_inst_bits&32'h18000020; 
  assign _id_ctrl_decoder_T_151=_id_ctrl_decoder_T_150==32'h18000020; 
  assign _id_ctrl_decoder_T_152=ibuf_io_inst_0_bits_inst_bits&32'h20000020; 
  assign _id_ctrl_decoder_T_153=_id_ctrl_decoder_T_152==32'h20000020; 
  assign _id_ctrl_decoder_T_155=_id_ctrl_decoder_T_149|_id_ctrl_decoder_T_151; 
  assign id_ctrl_decoder_lo_lo_1=_id_ctrl_decoder_T_155|_id_ctrl_decoder_T_153; 
  assign _id_ctrl_decoder_T_156=ibuf_io_inst_0_bits_inst_bits&32'h10000008; 
  assign _id_ctrl_decoder_T_157=_id_ctrl_decoder_T_156==32'h10000008; 
  assign _id_ctrl_decoder_T_158=ibuf_io_inst_0_bits_inst_bits&32'h40000008; 
  assign _id_ctrl_decoder_T_159=_id_ctrl_decoder_T_158==32'h40000008; 
  assign id_ctrl_decoder_lo_hi_1=_id_ctrl_decoder_T_157|_id_ctrl_decoder_T_159; 
  assign _id_ctrl_decoder_T_161=ibuf_io_inst_0_bits_inst_bits&32'h40; 
  assign id_ctrl_decoder_hi_hi_hi=_id_ctrl_decoder_T_161==32'h40; 
  assign _id_ctrl_decoder_T_163=ibuf_io_inst_0_bits_inst_bits&32'h8000008; 
  assign _id_ctrl_decoder_T_164=_id_ctrl_decoder_T_163==32'h8000008; 
  assign _id_ctrl_decoder_T_165=ibuf_io_inst_0_bits_inst_bits&32'h80000008; 
  assign _id_ctrl_decoder_T_166=_id_ctrl_decoder_T_165==32'h80000008; 
  assign _id_ctrl_decoder_T_168=id_ctrl_decoder_hi_hi_hi|_id_ctrl_decoder_T_164; 
  assign _id_ctrl_decoder_T_169=_id_ctrl_decoder_T_168|_id_ctrl_decoder_T_157; 
  assign id_ctrl_decoder_hi_lo_2=_id_ctrl_decoder_T_169|_id_ctrl_decoder_T_166; 
  assign _id_ctrl_decoder_T_170=ibuf_io_inst_0_bits_inst_bits&32'h18000008; 
  assign id_ctrl_decoder_hi_hi_lo=_id_ctrl_decoder_T_170==32'h8; 
  assign id_ctrl_decoder_15={id_ctrl_decoder_hi_hi_hi,id_ctrl_decoder_hi_hi_lo,id_ctrl_decoder_hi_lo_2,id_ctrl_decoder_lo_hi_1,id_ctrl_decoder_lo_lo_1}; 
  assign _id_ctrl_decoder_T_172=ibuf_io_inst_0_bits_inst_bits&32'h80000060; 
  assign _id_ctrl_decoder_T_173=_id_ctrl_decoder_T_172==32'h40; 
  assign _id_ctrl_decoder_T_174=ibuf_io_inst_0_bits_inst_bits&32'h10000060; 
  assign _id_ctrl_decoder_T_176=ibuf_io_inst_0_bits_inst_bits&32'h70; 
  assign id_ctrl_decoder_18=_id_ctrl_decoder_T_176==32'h40; 
  assign _id_ctrl_decoder_T_189=ibuf_io_inst_0_bits_inst_bits&32'h3c; 
  assign _id_ctrl_decoder_T_190=_id_ctrl_decoder_T_189==32'h4; 
  assign _id_ctrl_decoder_T_192=_id_ctrl_decoder_T_174==32'h10000040; 
  assign _id_ctrl_decoder_T_194=_id_ctrl_decoder_T_190|_id_ctrl_decoder_T_173; 
  assign _id_ctrl_decoder_T_195=_id_ctrl_decoder_T_194|id_ctrl_decoder_18; 
  assign id_ctrl_decoder_19=_id_ctrl_decoder_T_195|_id_ctrl_decoder_T_192; 
  assign _id_ctrl_decoder_T_196=ibuf_io_inst_0_bits_inst_bits&32'h2000074; 
  assign id_ctrl_decoder_21=_id_ctrl_decoder_T_196==32'h2000030; 
  assign _id_ctrl_decoder_T_199=_id_ctrl_decoder_T_11==32'h0; 
  assign _id_ctrl_decoder_T_201=_id_ctrl_decoder_T_61==32'h10; 
  assign _id_ctrl_decoder_T_202=ibuf_io_inst_0_bits_inst_bits&32'h2024; 
  assign _id_ctrl_decoder_T_203=_id_ctrl_decoder_T_202==32'h24; 
  assign _id_ctrl_decoder_T_204=ibuf_io_inst_0_bits_inst_bits&32'h28; 
  assign _id_ctrl_decoder_T_205=_id_ctrl_decoder_T_204==32'h28; 
  assign _id_ctrl_decoder_T_206=ibuf_io_inst_0_bits_inst_bits&32'h1030; 
  assign _id_ctrl_decoder_T_207=_id_ctrl_decoder_T_206==32'h1030; 
  assign _id_ctrl_decoder_T_208=ibuf_io_inst_0_bits_inst_bits&32'h2030; 
  assign _id_ctrl_decoder_T_209=_id_ctrl_decoder_T_208==32'h2030; 
  assign _id_ctrl_decoder_T_210=ibuf_io_inst_0_bits_inst_bits&32'h90000010; 
  assign _id_ctrl_decoder_T_211=_id_ctrl_decoder_T_210==32'h80000010; 
  assign _id_ctrl_decoder_T_213=_id_ctrl_decoder_T_199|_id_ctrl_decoder_T_201; 
  assign _id_ctrl_decoder_T_214=_id_ctrl_decoder_T_213|_id_ctrl_decoder_T_203; 
  assign _id_ctrl_decoder_T_215=_id_ctrl_decoder_T_214|_id_ctrl_decoder_T_205; 
  assign _id_ctrl_decoder_T_216=_id_ctrl_decoder_T_215|_id_ctrl_decoder_T_207; 
  assign _id_ctrl_decoder_T_217=_id_ctrl_decoder_T_216|_id_ctrl_decoder_T_209; 
  assign id_ctrl_decoder_22=_id_ctrl_decoder_T_217|_id_ctrl_decoder_T_211; 
  assign _id_ctrl_decoder_T_218=ibuf_io_inst_0_bits_inst_bits&32'h1070; 
  assign id_ctrl_decoder_lo_5=_id_ctrl_decoder_T_218==32'h1070; 
  assign _id_ctrl_decoder_T_220=ibuf_io_inst_0_bits_inst_bits&32'h2070; 
  assign id_ctrl_decoder_hi_lo_3=_id_ctrl_decoder_T_220==32'h2070; 
  assign _id_ctrl_decoder_T_222=ibuf_io_inst_0_bits_inst_bits&32'h10000070; 
  assign _id_ctrl_decoder_T_223=_id_ctrl_decoder_T_222==32'h70; 
  assign _id_ctrl_decoder_T_224=ibuf_io_inst_0_bits_inst_bits&32'h12000034; 
  assign _id_ctrl_decoder_T_225=_id_ctrl_decoder_T_224==32'h10000030; 
  assign _id_ctrl_decoder_T_226=ibuf_io_inst_0_bits_inst_bits&32'he0000050; 
  assign _id_ctrl_decoder_T_227=_id_ctrl_decoder_T_226==32'h60000050; 
  assign _id_ctrl_decoder_T_229=_id_ctrl_decoder_T_223|id_ctrl_decoder_lo_5; 
  assign _id_ctrl_decoder_T_230=_id_ctrl_decoder_T_229|id_ctrl_decoder_hi_lo_3; 
  assign _id_ctrl_decoder_T_231=_id_ctrl_decoder_T_230|_id_ctrl_decoder_T_225; 
  assign id_ctrl_decoder_hi_hi_3=_id_ctrl_decoder_T_231|_id_ctrl_decoder_T_227; 
  assign id_ctrl_decoder_23={id_ctrl_decoder_hi_hi_3,id_ctrl_decoder_hi_lo_3,id_ctrl_decoder_lo_5}; 
  assign _id_ctrl_decoder_T_232=ibuf_io_inst_0_bits_inst_bits&32'h3058; 
  assign id_ctrl_decoder_24=_id_ctrl_decoder_T_232==32'h1008; 
  assign id_ctrl_decoder_25=_id_ctrl_decoder_T_106==32'h8; 
  assign _id_ctrl_decoder_T_236=ibuf_io_inst_0_bits_inst_bits&32'h6048; 
  assign id_ctrl_decoder_26=_id_ctrl_decoder_T_236==32'h2008; 
  assign _id_ctrl_decoder_T_238=ibuf_io_inst_0_bits_inst_bits&32'h105c; 
  assign _id_ctrl_decoder_T_239=_id_ctrl_decoder_T_238==32'h1004; 
  assign _id_ctrl_decoder_T_240=ibuf_io_inst_0_bits_inst_bits&32'h2000060; 
  assign _id_ctrl_decoder_T_241=_id_ctrl_decoder_T_240==32'h2000040; 
  assign _id_ctrl_decoder_T_242=ibuf_io_inst_0_bits_inst_bits&32'hd0000070; 
  assign _id_ctrl_decoder_T_243=_id_ctrl_decoder_T_242==32'h40000050; 
  assign _id_ctrl_decoder_T_245=_id_ctrl_decoder_T_239|_id_ctrl_decoder_T_241; 
  assign id_ctrl_decoder_27=_id_ctrl_decoder_T_245|_id_ctrl_decoder_T_243; 
  assign id_raddr3=ibuf_io_inst_0_bits_inst_rs3; 
  assign id_raddr2=ibuf_io_inst_0_bits_inst_rs2; 
  assign id_raddr1=ibuf_io_inst_0_bits_inst_rs1; 
  assign id_waddr=ibuf_io_inst_0_bits_inst_rd; 
  assign _id_rs_T_4=rf_id_rs_MPORT_data; 
  assign _id_rs_T_9=rf_id_rs_MPORT_1_data; 
  assign _id_csr_en_T=id_ctrl_decoder_23==3'h6; 
  assign _id_csr_en_T_1=id_ctrl_decoder_23==3'h7; 
  assign _id_csr_en_T_2=id_ctrl_decoder_23==3'h5; 
  assign _id_csr_en_T_3=_id_csr_en_T|_id_csr_en_T_1; 
  assign id_csr_en=_id_csr_en_T_3|_id_csr_en_T_2; 
  assign id_system_insn=id_ctrl_decoder_23==3'h4; 
  assign _id_csr_ren_T_3=ibuf_io_inst_0_bits_inst_rs1==5'h0; 
  assign id_csr_ren=_id_csr_en_T_3&_id_csr_ren_T_3; 
  assign _id_sfence_T=id_ctrl_decoder_15==5'h14; 
  assign id_sfence=id_ctrl_decoder_14&_id_sfence_T; 
  assign _id_csr_flush_T=id_sfence|id_system_insn; 
  assign _id_csr_flush_T_2=id_csr_en&~id_csr_ren; 
  assign _id_csr_flush_T_3=_id_csr_flush_T_2&csr_io_decode_0_write_flush; 
  assign id_csr_flush=_id_csr_flush_T|_id_csr_flush_T_3; 
  assign _id_illegal_insn_T_4=id_ctrl_decoder_21&~csr_io_status_isa[12]; 
  assign _id_illegal_insn_T_5=~id_ctrl_decoder_0|_id_illegal_insn_T_4; 
  assign _id_illegal_insn_T_8=id_ctrl_decoder_26&~csr_io_status_isa[0]; 
  assign _id_illegal_insn_T_9=_id_illegal_insn_T_5|_id_illegal_insn_T_8; 
  assign _id_illegal_insn_T_10=csr_io_decode_0_fp_illegal|io_fpu_illegal_rm; 
  assign _id_illegal_insn_T_11=id_ctrl_decoder_1&_id_illegal_insn_T_10; 
  assign _id_illegal_insn_T_12=_id_illegal_insn_T_9|_id_illegal_insn_T_11; 
  assign _id_illegal_insn_T_15=id_ctrl_decoder_27&~csr_io_status_isa[3]; 
  assign _id_illegal_insn_T_16=_id_illegal_insn_T_12|_id_illegal_insn_T_15; 
  assign _id_illegal_insn_T_19=ibuf_io_inst_0_bits_rvc&~csr_io_status_isa[2]; 
  assign _id_illegal_insn_T_20=_id_illegal_insn_T_16|_id_illegal_insn_T_19; 
  assign _id_illegal_insn_T_40=~id_csr_ren&csr_io_decode_0_write_illegal; 
  assign _id_illegal_insn_T_41=csr_io_decode_0_read_illegal|_id_illegal_insn_T_40; 
  assign _id_illegal_insn_T_42=id_csr_en&_id_illegal_insn_T_41; 
  assign _id_illegal_insn_T_43=_id_illegal_insn_T_20|_id_illegal_insn_T_42; 
  assign _id_illegal_insn_T_46=_id_csr_flush_T&csr_io_decode_0_system_illegal; 
  assign _id_illegal_insn_T_47=~ibuf_io_inst_0_bits_rvc&_id_illegal_insn_T_46; 
  assign id_illegal_insn=_id_illegal_insn_T_43|_id_illegal_insn_T_47; 
  assign id_amo_aq=ibuf_io_inst_0_bits_inst_bits[26]; 
  assign id_amo_rl=ibuf_io_inst_0_bits_inst_bits[25]; 
  assign id_fence_succ=ibuf_io_inst_0_bits_inst_bits[23:20]; 
  assign _id_fence_next_T=id_ctrl_decoder_26&id_amo_aq; 
  assign id_fence_next=id_ctrl_decoder_25|_id_fence_next_T; 
  assign id_mem_busy=~io_dmem_ordered|io_dmem_req_valid; 
  assign _GEN_0=id_mem_busy ? id_reg_fence:1'h0; 
  assign _id_do_fence_x8_T_1=id_ctrl_decoder_26&id_amo_rl; 
  assign _id_do_fence_x8_T_2=_id_do_fence_x8_T_1|id_ctrl_decoder_24; 
  assign _id_do_fence_x8_T_4=id_reg_fence&id_ctrl_decoder_14; 
  assign _id_do_fence_x8_T_5=_id_do_fence_x8_T_2|_id_do_fence_x8_T_4; 
  assign id_do_fence_x8=id_mem_busy&_id_do_fence_x8_T_5; 
  assign _T_1=csr_io_interrupt|bpu_io_debug_if; 
  assign _T_2=_T_1|bpu_io_xcpt_if; 
  assign _T_3=_T_2|ibuf_io_inst_0_bits_xcpt0_pf_inst; 
  assign _T_4=_T_3|ibuf_io_inst_0_bits_xcpt0_ae_inst; 
  assign _T_5=_T_4|ibuf_io_inst_0_bits_xcpt1_pf_inst; 
  assign _T_6=_T_5|ibuf_io_inst_0_bits_xcpt1_ae_inst; 
  assign id_xcpt=_T_6|id_illegal_insn; 
  assign _T_7=ibuf_io_inst_0_bits_xcpt1_ae_inst ? 2'h1:2'h2; 
  assign _T_8=ibuf_io_inst_0_bits_xcpt1_pf_inst ? 4'hc:{2'b0,_T_7}; 
  assign _T_9=ibuf_io_inst_0_bits_xcpt0_ae_inst ? 4'h1:_T_8; 
  assign _T_10=ibuf_io_inst_0_bits_xcpt0_pf_inst ? 4'hc:_T_9; 
  assign _T_11=bpu_io_xcpt_if ? 4'h3:_T_10; 
  assign _T_12=bpu_io_debug_if ? 4'he:_T_11; 
  assign ex_waddr=ex_reg_inst[11:7]; 
  assign mem_waddr=mem_reg_inst[11:7]; 
  assign wb_waddr=wb_reg_inst[11:7]; 
  assign _T_23=ex_reg_valid&ex_ctrl_wxd; 
  assign _T_24=mem_reg_valid&mem_ctrl_wxd; 
  assign _T_26=_T_24&~mem_ctrl_mem; 
  assign id_bypass_src_0_0=5'h0==id_raddr1; 
  assign _id_bypass_src_T_1=ex_waddr==id_raddr1; 
  assign id_bypass_src_0_1=_T_23&_id_bypass_src_T_1; 
  assign _id_bypass_src_T_2=mem_waddr==id_raddr1; 
  assign id_bypass_src_0_2=_T_26&_id_bypass_src_T_2; 
  assign id_bypass_src_0_3=_T_24&_id_bypass_src_T_2; 
  assign id_bypass_src_1_0=5'h0==id_raddr2; 
  assign _id_bypass_src_T_5=ex_waddr==id_raddr2; 
  assign id_bypass_src_1_1=_T_23&_id_bypass_src_T_5; 
  assign _id_bypass_src_T_6=mem_waddr==id_raddr2; 
  assign id_bypass_src_1_2=_T_26&_id_bypass_src_T_6; 
  assign id_bypass_src_1_3=_T_24&_id_bypass_src_T_6; 
  assign _ex_rs_T=ex_reg_rs_lsb_0==2'h1; 
  assign _ex_rs_T_1=_ex_rs_T ? mem_reg_wdata:64'h0; 
  assign _ex_rs_T_2=ex_reg_rs_lsb_0==2'h2; 
  assign _ex_rs_T_3=_ex_rs_T_2 ? wb_reg_wdata:_ex_rs_T_1; 
  assign _ex_rs_T_4=ex_reg_rs_lsb_0==2'h3; 
  assign _ex_rs_T_5=_ex_rs_T_4 ? io_dmem_resp_bits_data_word_bypass:_ex_rs_T_3; 
  assign _ex_rs_T_6={ex_reg_rs_msb_0,ex_reg_rs_lsb_0}; 
  assign _ex_rs_T_7=ex_reg_rs_lsb_1==2'h1; 
  assign _ex_rs_T_8=_ex_rs_T_7 ? mem_reg_wdata:64'h0; 
  assign _ex_rs_T_9=ex_reg_rs_lsb_1==2'h2; 
  assign _ex_rs_T_10=_ex_rs_T_9 ? wb_reg_wdata:_ex_rs_T_8; 
  assign _ex_rs_T_11=ex_reg_rs_lsb_1==2'h3; 
  assign _ex_rs_T_12=_ex_rs_T_11 ? io_dmem_resp_bits_data_word_bypass:_ex_rs_T_10; 
  assign _ex_rs_T_13={ex_reg_rs_msb_1,ex_reg_rs_lsb_1}; 
  assign ex_rs_1=ex_reg_rs_bypass_1 ? _ex_rs_T_12:_ex_rs_T_13; 
  assign _ex_imm_sign_T=ex_ctrl_sel_imm==3'h5; 
  assign _ex_imm_sign_T_2=ex_reg_inst[31]; 
  assign ex_imm_sign=_ex_imm_sign_T ? $signed(1'sh0):$signed(_ex_imm_sign_T_2); 
  assign _ex_imm_b30_20_T=ex_ctrl_sel_imm==3'h2; 
  assign _ex_imm_b30_20_T_2=ex_reg_inst[30:20]; 
  assign _ex_imm_b19_12_T=ex_ctrl_sel_imm!=3'h2; 
  assign _ex_imm_b19_12_T_1=ex_ctrl_sel_imm!=3'h3; 
  assign _ex_imm_b19_12_T_2=_ex_imm_b19_12_T&_ex_imm_b19_12_T_1; 
  assign _ex_imm_b19_12_T_4=ex_reg_inst[19:12]; 
  assign _ex_imm_b11_T_2=_ex_imm_b30_20_T|_ex_imm_sign_T; 
  assign _ex_imm_b11_T_3=ex_ctrl_sel_imm==3'h3; 
  assign _ex_imm_b11_T_5=ex_reg_inst[20]; 
  assign _ex_imm_b11_T_6=ex_ctrl_sel_imm==3'h1; 
  assign _ex_imm_b11_T_8=ex_reg_inst[7]; 
  assign _ex_imm_b11_T_9=_ex_imm_b11_T_6 ? $signed(_ex_imm_b11_T_8):$signed(ex_imm_sign); 
  assign _ex_imm_b11_T_10=_ex_imm_b11_T_3 ? $signed(_ex_imm_b11_T_5):$signed(_ex_imm_b11_T_9); 
  assign ex_imm_lo_hi_hi=_ex_imm_b11_T_2 ? 6'h0:ex_reg_inst[30:25]; 
  assign _ex_imm_b4_1_T_1=ex_ctrl_sel_imm==3'h0; 
  assign _ex_imm_b4_1_T_3=_ex_imm_b4_1_T_1|_ex_imm_b11_T_6; 
  assign _ex_imm_b4_1_T_8=_ex_imm_sign_T ? ex_reg_inst[19:16]:ex_reg_inst[24:21]; 
  assign _ex_imm_b4_1_T_9=_ex_imm_b4_1_T_3 ? ex_reg_inst[11:8]:_ex_imm_b4_1_T_8; 
  assign ex_imm_lo_hi_lo=_ex_imm_b30_20_T ? 4'h0:_ex_imm_b4_1_T_9; 
  assign _ex_imm_b0_T_2=ex_ctrl_sel_imm==3'h4; 
  assign _ex_imm_b0_T_6=_ex_imm_sign_T&ex_reg_inst[15]; 
  assign _ex_imm_b0_T_7=_ex_imm_b0_T_2 ? ex_reg_inst[20]:_ex_imm_b0_T_6; 
  assign ex_imm_lo_lo=_ex_imm_b4_1_T_1 ? ex_reg_inst[7]:_ex_imm_b0_T_7; 
  assign ex_imm_hi_lo_lo=_ex_imm_b11_T_2 ? $signed(1'sh0):$signed(_ex_imm_b11_T_10); 
  assign ex_imm_hi_lo_hi=_ex_imm_b19_12_T_2 ? $signed({8{ex_imm_sign}}):$signed(_ex_imm_b19_12_T_4); 
  assign ex_imm_hi_hi_lo=_ex_imm_b30_20_T ? $signed(_ex_imm_b30_20_T_2):$signed({11{ex_imm_sign}}); 
  assign ex_imm_hi_hi_hi=_ex_imm_sign_T ? $signed(1'sh0):$signed(_ex_imm_sign_T_2); 
  assign ex_imm={ex_imm_hi_hi_hi,ex_imm_hi_hi_lo,ex_imm_hi_lo_hi,ex_imm_hi_lo_lo,ex_imm_lo_hi_hi,ex_imm_lo_hi_lo,ex_imm_lo_lo}; 
  assign _ex_op1_T=ex_reg_rs_bypass_0 ? _ex_rs_T_5:_ex_rs_T_6; 
  assign _ex_op1_T_2=2'h1==ex_ctrl_sel_alu1; 
  assign _ex_op1_T_3=_ex_op1_T_2 ? $signed(_ex_op1_T):$signed(64'sh0); 
  assign _ex_op1_T_4=2'h2==ex_ctrl_sel_alu1; 
  assign _ex_op2_T=ex_reg_rs_bypass_1 ? _ex_rs_T_12:_ex_rs_T_13; 
  assign _ex_op2_T_1=ex_reg_rvc ? $signed(4'sh2):$signed(4'sh4); 
  assign _ex_op2_T_2=2'h2==ex_ctrl_sel_alu2; 
  assign _ex_op2_T_3=_ex_op2_T_2 ? $signed(_ex_op2_T):$signed(64'sh0); 
  assign _ex_op2_T_4=2'h3==ex_ctrl_sel_alu2; 
  assign _ex_op2_T_5=_ex_op2_T_4 ? $signed({{32{ex_imm[31]}},ex_imm}):$signed(_ex_op2_T_3); 
  assign _ex_op2_T_6=2'h1==ex_ctrl_sel_alu2; 
  assign _ctrl_killd_T_1=~ibuf_io_inst_0_valid|ibuf_io_inst_0_bits_replay; 
  assign _ctrl_killd_T_2=_ctrl_killd_T_1|take_pc_mem_wb; 
  assign _T_123=id_raddr1!=5'h0; 
  assign _T_124=id_ctrl_decoder_7&_T_123; 
  assign _data_hazard_ex_T=id_raddr1==ex_waddr; 
  assign _data_hazard_ex_T_1=_T_124&_data_hazard_ex_T; 
  assign _T_125=id_raddr2!=5'h0; 
  assign _T_126=id_ctrl_decoder_6&_T_125; 
  assign _data_hazard_ex_T_2=id_raddr2==ex_waddr; 
  assign _data_hazard_ex_T_3=_T_126&_data_hazard_ex_T_2; 
  assign _data_hazard_ex_T_6=_data_hazard_ex_T_1|_data_hazard_ex_T_3; 
  assign _T_127=id_waddr!=5'h0; 
  assign _T_128=id_ctrl_decoder_22&_T_127; 
  assign _data_hazard_ex_T_4=id_waddr==ex_waddr; 
  assign _data_hazard_ex_T_5=_T_128&_data_hazard_ex_T_4; 
  assign _data_hazard_ex_T_7=_data_hazard_ex_T_6|_data_hazard_ex_T_5; 
  assign data_hazard_ex=ex_ctrl_wxd&_data_hazard_ex_T_7; 
  assign _ex_cannot_bypass_T=ex_ctrl_csr!=3'h0; 
  assign _ex_cannot_bypass_T_1=_ex_cannot_bypass_T|ex_ctrl_jalr; 
  assign _ex_cannot_bypass_T_2=_ex_cannot_bypass_T_1|ex_ctrl_mem; 
  assign _ex_cannot_bypass_T_4=_ex_cannot_bypass_T_2|ex_ctrl_div; 
  assign ex_cannot_bypass=_ex_cannot_bypass_T_4|ex_ctrl_fp; 
  assign _id_ex_hazard_T=data_hazard_ex&ex_cannot_bypass; 
  assign _fp_data_hazard_ex_T_1=io_fpu_dec_ren1&_data_hazard_ex_T; 
  assign _fp_data_hazard_ex_T_3=io_fpu_dec_ren2&_data_hazard_ex_T_2; 
  assign _fp_data_hazard_ex_T_8=_fp_data_hazard_ex_T_1|_fp_data_hazard_ex_T_3; 
  assign _fp_data_hazard_ex_T_4=id_raddr3==ex_waddr; 
  assign _fp_data_hazard_ex_T_5=io_fpu_dec_ren3&_fp_data_hazard_ex_T_4; 
  assign _fp_data_hazard_ex_T_9=_fp_data_hazard_ex_T_8|_fp_data_hazard_ex_T_5; 
  assign _fp_data_hazard_ex_T_7=io_fpu_dec_wen&_data_hazard_ex_T_4; 
  assign _fp_data_hazard_ex_T_10=_fp_data_hazard_ex_T_9|_fp_data_hazard_ex_T_7; 
  assign fp_data_hazard_ex=ex_ctrl_wfd&_fp_data_hazard_ex_T_10; 
  assign _id_ex_hazard_T_1=_id_ex_hazard_T|fp_data_hazard_ex; 
  assign id_ex_hazard=ex_reg_valid&_id_ex_hazard_T_1; 
  assign _data_hazard_mem_T=id_raddr1==mem_waddr; 
  assign _data_hazard_mem_T_1=_T_124&_data_hazard_mem_T; 
  assign _data_hazard_mem_T_2=id_raddr2==mem_waddr; 
  assign _data_hazard_mem_T_3=_T_126&_data_hazard_mem_T_2; 
  assign _data_hazard_mem_T_6=_data_hazard_mem_T_1|_data_hazard_mem_T_3; 
  assign _data_hazard_mem_T_4=id_waddr==mem_waddr; 
  assign _data_hazard_mem_T_5=_T_128&_data_hazard_mem_T_4; 
  assign _data_hazard_mem_T_7=_data_hazard_mem_T_6|_data_hazard_mem_T_5; 
  assign data_hazard_mem=mem_ctrl_wxd&_data_hazard_mem_T_7; 
  assign _mem_cannot_bypass_T=mem_ctrl_csr!=3'h0; 
  assign _mem_cannot_bypass_T_1=mem_ctrl_mem&mem_reg_slow_bypass; 
  assign _mem_cannot_bypass_T_2=_mem_cannot_bypass_T|_mem_cannot_bypass_T_1; 
  assign _mem_cannot_bypass_T_4=_mem_cannot_bypass_T_2|mem_ctrl_div; 
  assign mem_cannot_bypass=_mem_cannot_bypass_T_4|mem_ctrl_fp; 
  assign _id_mem_hazard_T=data_hazard_mem&mem_cannot_bypass; 
  assign _fp_data_hazard_mem_T_1=io_fpu_dec_ren1&_data_hazard_mem_T; 
  assign _fp_data_hazard_mem_T_3=io_fpu_dec_ren2&_data_hazard_mem_T_2; 
  assign _fp_data_hazard_mem_T_8=_fp_data_hazard_mem_T_1|_fp_data_hazard_mem_T_3; 
  assign _fp_data_hazard_mem_T_4=id_raddr3==mem_waddr; 
  assign _fp_data_hazard_mem_T_5=io_fpu_dec_ren3&_fp_data_hazard_mem_T_4; 
  assign _fp_data_hazard_mem_T_9=_fp_data_hazard_mem_T_8|_fp_data_hazard_mem_T_5; 
  assign _fp_data_hazard_mem_T_7=io_fpu_dec_wen&_data_hazard_mem_T_4; 
  assign _fp_data_hazard_mem_T_10=_fp_data_hazard_mem_T_9|_fp_data_hazard_mem_T_7; 
  assign fp_data_hazard_mem=mem_ctrl_wfd&_fp_data_hazard_mem_T_10; 
  assign _id_mem_hazard_T_1=_id_mem_hazard_T|fp_data_hazard_mem; 
  assign id_mem_hazard=mem_reg_valid&_id_mem_hazard_T_1; 
  assign _ctrl_stalld_T=id_ex_hazard|id_mem_hazard; 
  assign _data_hazard_wb_T=id_raddr1==wb_waddr; 
  assign _data_hazard_wb_T_1=_T_124&_data_hazard_wb_T; 
  assign _data_hazard_wb_T_2=id_raddr2==wb_waddr; 
  assign _data_hazard_wb_T_3=_T_126&_data_hazard_wb_T_2; 
  assign _data_hazard_wb_T_6=_data_hazard_wb_T_1|_data_hazard_wb_T_3; 
  assign _data_hazard_wb_T_4=id_waddr==wb_waddr; 
  assign _data_hazard_wb_T_5=_T_128&_data_hazard_wb_T_4; 
  assign _data_hazard_wb_T_7=_data_hazard_wb_T_6|_data_hazard_wb_T_5; 
  assign data_hazard_wb=wb_ctrl_wxd&_data_hazard_wb_T_7; 
  assign wb_dcache_miss=wb_ctrl_mem&~io_dmem_resp_valid; 
  assign wb_set_sboard=wb_ctrl_div|wb_dcache_miss; 
  assign _id_wb_hazard_T=data_hazard_wb&wb_set_sboard; 
  assign _fp_data_hazard_wb_T_1=io_fpu_dec_ren1&_data_hazard_wb_T; 
  assign _fp_data_hazard_wb_T_3=io_fpu_dec_ren2&_data_hazard_wb_T_2; 
  assign _fp_data_hazard_wb_T_8=_fp_data_hazard_wb_T_1|_fp_data_hazard_wb_T_3; 
  assign _fp_data_hazard_wb_T_4=id_raddr3==wb_waddr; 
  assign _fp_data_hazard_wb_T_5=io_fpu_dec_ren3&_fp_data_hazard_wb_T_4; 
  assign _fp_data_hazard_wb_T_9=_fp_data_hazard_wb_T_8|_fp_data_hazard_wb_T_5; 
  assign _fp_data_hazard_wb_T_7=io_fpu_dec_wen&_data_hazard_wb_T_4; 
  assign _fp_data_hazard_wb_T_10=_fp_data_hazard_wb_T_9|_fp_data_hazard_wb_T_7; 
  assign fp_data_hazard_wb=wb_ctrl_wfd&_fp_data_hazard_wb_T_10; 
  assign _id_wb_hazard_T_1=_id_wb_hazard_T|fp_data_hazard_wb; 
  assign id_wb_hazard=wb_reg_valid&_id_wb_hazard_T_1; 
  assign _ctrl_stalld_T_1=_ctrl_stalld_T|id_wb_hazard; 
  assign r={_r[31:1],1'h0}; 
  assign _id_sboard_hazard_T=r>>id_raddr1; 
  assign dmem_resp_valid=io_dmem_resp_valid&io_dmem_resp_bits_has_data; 
  assign dmem_resp_replay=dmem_resp_valid&io_dmem_resp_bits_replay; 
  assign dmem_resp_xpu=~io_dmem_resp_bits_tag[0]; 
  assign _T_117=dmem_resp_replay&dmem_resp_xpu; 
  assign ll_wen_x1=div_io_resp_ready&div_io_resp_valid; 
  assign ll_wen=_T_117|ll_wen_x1; 
  assign dmem_resp_waddr=io_dmem_resp_bits_tag[5:1]; 
  assign ll_waddr=_T_117 ? dmem_resp_waddr:div_io_resp_bits_tag; 
  assign _id_sboard_hazard_T_2=ll_waddr==id_raddr1; 
  assign _id_sboard_hazard_T_3=ll_wen&_id_sboard_hazard_T_2; 
  assign _id_sboard_hazard_T_5=_id_sboard_hazard_T[0]&~_id_sboard_hazard_T_3; 
  assign _id_sboard_hazard_T_6=_T_124&_id_sboard_hazard_T_5; 
  assign _id_sboard_hazard_T_7=r>>id_raddr2; 
  assign _id_sboard_hazard_T_9=ll_waddr==id_raddr2; 
  assign _id_sboard_hazard_T_10=ll_wen&_id_sboard_hazard_T_9; 
  assign _id_sboard_hazard_T_12=_id_sboard_hazard_T_7[0]&~_id_sboard_hazard_T_10; 
  assign _id_sboard_hazard_T_13=_T_126&_id_sboard_hazard_T_12; 
  assign _id_sboard_hazard_T_21=_id_sboard_hazard_T_6|_id_sboard_hazard_T_13; 
  assign _id_sboard_hazard_T_14=r>>id_waddr; 
  assign _id_sboard_hazard_T_16=ll_waddr==id_waddr; 
  assign _id_sboard_hazard_T_17=ll_wen&_id_sboard_hazard_T_16; 
  assign _id_sboard_hazard_T_19=_id_sboard_hazard_T_14[0]&~_id_sboard_hazard_T_17; 
  assign _id_sboard_hazard_T_20=_T_128&_id_sboard_hazard_T_19; 
  assign id_sboard_hazard=_id_sboard_hazard_T_21|_id_sboard_hazard_T_20; 
  assign _ctrl_stalld_T_2=_ctrl_stalld_T_1|id_sboard_hazard; 
  assign _ctrl_stalld_T_3=ex_reg_valid|mem_reg_valid; 
  assign _ctrl_stalld_T_4=_ctrl_stalld_T_3|wb_reg_valid; 
  assign _ctrl_stalld_T_5=csr_io_singleStep&_ctrl_stalld_T_4; 
  assign _ctrl_stalld_T_6=_ctrl_stalld_T_2|_ctrl_stalld_T_5; 
  assign _ctrl_stalld_T_7=id_csr_en&csr_io_decode_0_fp_csr; 
  assign _ctrl_stalld_T_9=_ctrl_stalld_T_7&~io_fpu_fcsr_rdy; 
  assign _ctrl_stalld_T_10=_ctrl_stalld_T_6|_ctrl_stalld_T_9; 
  assign _id_stall_fpu_T_18=id_stall_fpu__r>>id_raddr1; 
  assign _id_stall_fpu_T_20=io_fpu_dec_ren1&_id_stall_fpu_T_18[0]; 
  assign _id_stall_fpu_T_21=id_stall_fpu__r>>id_raddr2; 
  assign _id_stall_fpu_T_23=io_fpu_dec_ren2&_id_stall_fpu_T_21[0]; 
  assign _id_stall_fpu_T_30=_id_stall_fpu_T_20|_id_stall_fpu_T_23; 
  assign _id_stall_fpu_T_24=id_stall_fpu__r>>id_raddr3; 
  assign _id_stall_fpu_T_26=io_fpu_dec_ren3&_id_stall_fpu_T_24[0]; 
  assign _id_stall_fpu_T_31=_id_stall_fpu_T_30|_id_stall_fpu_T_26; 
  assign _id_stall_fpu_T_27=id_stall_fpu__r>>id_waddr; 
  assign _id_stall_fpu_T_29=io_fpu_dec_wen&_id_stall_fpu_T_27[0]; 
  assign id_stall_fpu=_id_stall_fpu_T_31|_id_stall_fpu_T_29; 
  assign _ctrl_stalld_T_11=id_ctrl_decoder_1&id_stall_fpu; 
  assign _ctrl_stalld_T_12=_ctrl_stalld_T_10|_ctrl_stalld_T_11; 
  assign dcache_blocked=blocked&~io_dmem_perf_grant; 
  assign _ctrl_stalld_T_13=id_ctrl_decoder_14&dcache_blocked; 
  assign _ctrl_stalld_T_14=_ctrl_stalld_T_12|_ctrl_stalld_T_13; 
  assign wb_wxd=wb_reg_valid&wb_ctrl_wxd; 
  assign _ctrl_stalld_T_18=div_io_resp_valid&~wb_wxd; 
  assign _ctrl_stalld_T_19=div_io_req_ready|_ctrl_stalld_T_18; 
  assign _ctrl_stalld_T_21=~_ctrl_stalld_T_19|div_io_req_valid; 
  assign _ctrl_stalld_T_22=id_ctrl_decoder_21&_ctrl_stalld_T_21; 
  assign _ctrl_stalld_T_23=_ctrl_stalld_T_14|_ctrl_stalld_T_22; 
  assign _ctrl_stalld_T_26=_ctrl_stalld_T_23|id_do_fence_x8; 
  assign _ctrl_stalld_T_27=_ctrl_stalld_T_26|csr_io_csr_stall; 
  assign ctrl_stalld=_ctrl_stalld_T_27|id_reg_pause; 
  assign _ctrl_killd_T_3=_ctrl_killd_T_2|ctrl_stalld; 
  assign ctrl_killd=_ctrl_killd_T_3|csr_io_interrupt; 
  assign _ex_reg_replay_T_1=~take_pc_mem_wb&ibuf_io_inst_0_valid; 
  assign _T_29=id_fence_succ==4'h0; 
  assign _T_30=id_ctrl_decoder_25&_T_29; 
  assign _GEN_1=_T_30|id_reg_pause; 
  assign _GEN_2=id_fence_next|_GEN_0; 
  assign _T_31={ibuf_io_inst_0_bits_xcpt1_pf_inst,ibuf_io_inst_0_bits_xcpt1_ae_inst}; 
  assign _T_32=|_T_31; 
  assign _GEN_5=_T_32|ibuf_io_inst_0_bits_rvc; 
  assign _T_33={ibuf_io_inst_0_bits_xcpt0_pf_inst,ibuf_io_inst_0_bits_xcpt0_ae_inst}; 
  assign _T_34=|_T_33; 
  assign _T_35=bpu_io_xcpt_if|_T_34; 
  assign _GEN_9=id_xcpt|id_ctrl_decoder_12; 
  assign _ex_reg_flush_pipe_T=id_ctrl_decoder_24|id_csr_flush; 
  assign _T_37=id_ctrl_decoder_15==5'h5; 
  assign _T_38=_id_sfence_T|_T_37; 
  assign _ex_reg_mem_size_T_1={_T_125,_T_123}; 
  assign _do_bypass_T=id_bypass_src_0_0|id_bypass_src_0_1; 
  assign _do_bypass_T_1=_do_bypass_T|id_bypass_src_0_2; 
  assign do_bypass=_do_bypass_T_1|id_bypass_src_0_3; 
  assign _T_40=id_ctrl_decoder_7&~do_bypass; 
  assign _wb_valid_T_1=wb_reg_valid&~replay_wb_common; 
  assign wb_valid=_wb_valid_T_1&~wb_xcpt; 
  assign wb_wen=wb_valid&wb_ctrl_wxd; 
  assign rf_wen=wb_wen|ll_wen; 
  assign rf_waddr=ll_wen ? ll_waddr:wb_waddr; 
  assign _T_118=rf_waddr!=5'h0; 
  assign _T_121=rf_waddr==id_raddr1; 
  assign _rf_wdata_T=dmem_resp_valid&dmem_resp_xpu; 
  assign ll_wdata=div_io_resp_bits_data; 
  assign _rf_wdata_T_2=wb_ctrl_csr!=3'h0; 
  assign _rf_wdata_T_4=_rf_wdata_T_2 ? csr_io_rw_rdata:wb_reg_wdata; 
  assign _rf_wdata_T_5=ll_wen ? ll_wdata:_rf_wdata_T_4; 
  assign rf_wdata=_rf_wdata_T ? io_dmem_resp_bits_data:_rf_wdata_T_5; 
  assign _GEN_226=_T_121 ? rf_wdata:_id_rs_T_4; 
  assign _GEN_233=_T_118 ? _GEN_226:_id_rs_T_4; 
  assign id_rs_0=rf_wen ? _GEN_233:_id_rs_T_4; 
  assign _do_bypass_T_2=id_bypass_src_1_0|id_bypass_src_1_1; 
  assign _do_bypass_T_3=_do_bypass_T_2|id_bypass_src_1_2; 
  assign do_bypass_1=_do_bypass_T_3|id_bypass_src_1_3; 
  assign _T_42=id_ctrl_decoder_6&~do_bypass_1; 
  assign _T_122=rf_waddr==id_raddr2; 
  assign _GEN_227=_T_122 ? rf_wdata:_id_rs_T_9; 
  assign _GEN_234=_T_118 ? _GEN_227:_id_rs_T_9; 
  assign id_rs_1=rf_wen ? _GEN_234:_id_rs_T_9; 
  assign inst=ibuf_io_inst_0_bits_rvc ? {16'b0,ibuf_io_inst_0_bits_raw[15:0]}:ibuf_io_inst_0_bits_raw; 
  assign _id_load_use_T=mem_reg_valid&data_hazard_mem; 
  assign id_load_use=_id_load_use_T&mem_ctrl_mem; 
  assign _T_44=~ctrl_killd|csr_io_interrupt; 
  assign _T_45=_T_44|ibuf_io_inst_0_bits_replay; 
  assign _replay_ex_structural_T_1=ex_ctrl_mem&~io_dmem_req_ready; 
  assign _replay_ex_structural_T_3=ex_ctrl_div&~div_io_req_ready; 
  assign replay_ex_structural=_replay_ex_structural_T_1|_replay_ex_structural_T_3; 
  assign replay_ex_load_use=wb_dcache_miss&ex_reg_load_use; 
  assign _replay_ex_T=replay_ex_structural|replay_ex_load_use; 
  assign _replay_ex_T_1=ex_reg_valid&_replay_ex_T; 
  assign replay_ex=ex_reg_replay|_replay_ex_T_1; 
  assign _ctrl_killx_T=take_pc_mem_wb|replay_ex; 
  assign ctrl_killx=_ctrl_killx_T|~ex_reg_valid; 
  assign _ex_slow_bypass_T=ex_ctrl_mem_cmd==5'h7; 
  assign _ex_slow_bypass_T_1=ex_reg_mem_size<2'h2; 
  assign ex_slow_bypass=_ex_slow_bypass_T|_ex_slow_bypass_T_1; 
  assign _ex_sfence_T_1=ex_ctrl_mem_cmd==5'h14; 
  assign ex_sfence=ex_ctrl_mem&_ex_sfence_T_1; 
  assign ex_xcpt=ex_reg_xcpt_interrupt|ex_reg_xcpt; 
  assign _mem_pc_valid_T=mem_reg_valid|mem_reg_replay; 
  assign mem_pc_valid=_mem_pc_valid_T|mem_reg_xcpt_interrupt; 
  assign _mem_npc_misaligned_T_3=~csr_io_status_isa[2]&mem_npc[1]; 
  assign mem_npc_misaligned=_mem_npc_misaligned_T_3&~mem_reg_sfence; 
  assign _mem_int_wdata_T_1=mem_ctrl_jalr^mem_npc_misaligned; 
  assign _mem_int_wdata_T_2=~mem_reg_xcpt&_mem_int_wdata_T_1; 
  assign mem_int_wdata=_mem_int_wdata_T_2 ? $signed({{24{mem_br_target[39]}},mem_br_target}):$signed(mem_reg_wdata); 
  assign _mem_cfi_T=mem_ctrl_branch|mem_ctrl_jalr; 
  assign mem_cfi=_mem_cfi_T|mem_ctrl_jal; 
  assign _mem_cfi_taken_T_1=_mem_br_target_T_1|mem_ctrl_jalr; 
  assign mem_cfi_taken=_mem_cfi_taken_T_1|mem_ctrl_jal; 
  assign _T_56=mem_reg_valid&mem_reg_flush_pipe; 
  assign _mem_reg_load_T=ex_ctrl_mem_cmd==5'h0; 
  assign _mem_reg_load_T_1=ex_ctrl_mem_cmd==5'h6; 
  assign _mem_reg_load_T_2=_mem_reg_load_T|_mem_reg_load_T_1; 
  assign _mem_reg_load_T_4=_mem_reg_load_T_2|_ex_slow_bypass_T; 
  assign _mem_reg_load_T_5=ex_ctrl_mem_cmd==5'h4; 
  assign _mem_reg_load_T_6=ex_ctrl_mem_cmd==5'h9; 
  assign _mem_reg_load_T_7=ex_ctrl_mem_cmd==5'ha; 
  assign _mem_reg_load_T_8=ex_ctrl_mem_cmd==5'hb; 
  assign _mem_reg_load_T_9=_mem_reg_load_T_5|_mem_reg_load_T_6; 
  assign _mem_reg_load_T_10=_mem_reg_load_T_9|_mem_reg_load_T_7; 
  assign _mem_reg_load_T_11=_mem_reg_load_T_10|_mem_reg_load_T_8; 
  assign _mem_reg_load_T_12=ex_ctrl_mem_cmd==5'h8; 
  assign _mem_reg_load_T_13=ex_ctrl_mem_cmd==5'hc; 
  assign _mem_reg_load_T_14=ex_ctrl_mem_cmd==5'hd; 
  assign _mem_reg_load_T_15=ex_ctrl_mem_cmd==5'he; 
  assign _mem_reg_load_T_16=ex_ctrl_mem_cmd==5'hf; 
  assign _mem_reg_load_T_17=_mem_reg_load_T_12|_mem_reg_load_T_13; 
  assign _mem_reg_load_T_18=_mem_reg_load_T_17|_mem_reg_load_T_14; 
  assign _mem_reg_load_T_19=_mem_reg_load_T_18|_mem_reg_load_T_15; 
  assign _mem_reg_load_T_20=_mem_reg_load_T_19|_mem_reg_load_T_16; 
  assign _mem_reg_load_T_21=_mem_reg_load_T_11|_mem_reg_load_T_20; 
  assign _mem_reg_load_T_22=_mem_reg_load_T_4|_mem_reg_load_T_21; 
  assign _mem_reg_load_T_23=ex_ctrl_mem&_mem_reg_load_T_22; 
  assign _mem_reg_store_T=ex_ctrl_mem_cmd==5'h1; 
  assign _mem_reg_store_T_1=ex_ctrl_mem_cmd==5'h11; 
  assign _mem_reg_store_T_2=_mem_reg_store_T|_mem_reg_store_T_1; 
  assign _mem_reg_store_T_4=_mem_reg_store_T_2|_ex_slow_bypass_T; 
  assign _mem_reg_store_T_22=_mem_reg_store_T_4|_mem_reg_load_T_21; 
  assign _mem_reg_store_T_23=ex_ctrl_mem&_mem_reg_store_T_22; 
  assign _mem_reg_wdata_T=alu_io_out; 
  assign _T_58=ex_ctrl_mem|ex_sfence; 
  assign _T_59=ex_ctrl_rxs2&_T_58; 
  assign _mem_reg_rs2_T=ex_reg_mem_size==2'h0; 
  assign mem_reg_rs2_hi=ex_rs_1[7:0]; 
  assign _mem_reg_rs2_T_1={mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi,mem_reg_rs2_hi}; 
  assign _mem_reg_rs2_T_2=ex_reg_mem_size==2'h1; 
  assign mem_reg_rs2_hi_3=ex_rs_1[15:0]; 
  assign _mem_reg_rs2_T_3={mem_reg_rs2_hi_3,mem_reg_rs2_hi_3,mem_reg_rs2_hi_3,mem_reg_rs2_hi_3}; 
  assign _mem_reg_rs2_T_4=ex_reg_mem_size==2'h2; 
  assign mem_reg_rs2_hi_5=ex_rs_1[31:0]; 
  assign _mem_reg_rs2_T_5={mem_reg_rs2_hi_5,mem_reg_rs2_hi_5}; 
  assign _T_60=ex_ctrl_jalr&csr_io_status_debug; 
  assign _GEN_77=_T_60|ex_ctrl_fence_i; 
  assign _GEN_78=_T_60|ex_reg_flush_pipe; 
  assign _mem_breakpoint_T=mem_reg_load&bpu_io_xcpt_ld; 
  assign _mem_breakpoint_T_1=mem_reg_store&bpu_io_xcpt_st; 
  assign mem_breakpoint=_mem_breakpoint_T|_mem_breakpoint_T_1; 
  assign _mem_debug_breakpoint_T=mem_reg_load&bpu_io_debug_ld; 
  assign _mem_debug_breakpoint_T_1=mem_reg_store&bpu_io_debug_st; 
  assign mem_debug_breakpoint=_mem_debug_breakpoint_T|_mem_debug_breakpoint_T_1; 
  assign mem_ldst_xcpt=mem_debug_breakpoint|mem_breakpoint; 
  assign mem_ldst_cause=mem_debug_breakpoint ? 4'he:4'h3; 
  assign _T_61=mem_reg_xcpt_interrupt|mem_reg_xcpt; 
  assign _T_62=mem_reg_valid&mem_npc_misaligned; 
  assign _T_63=mem_reg_valid&mem_ldst_xcpt; 
  assign _T_64=_T_61|_T_62; 
  assign mem_xcpt=_T_64|_T_63; 
  assign _T_65=_T_62 ? 4'h0:mem_ldst_cause; 
  assign dcache_kill_mem=_T_24&io_dmem_replay_next; 
  assign _fpu_kill_mem_T=mem_reg_valid&mem_ctrl_fp; 
  assign fpu_kill_mem=_fpu_kill_mem_T&io_fpu_nack_mem; 
  assign _replay_mem_T=dcache_kill_mem|mem_reg_replay; 
  assign replay_mem=_replay_mem_T|fpu_kill_mem; 
  assign _killm_common_T=dcache_kill_mem|take_pc_wb; 
  assign _killm_common_T_1=_killm_common_T|mem_reg_xcpt; 
  assign killm_common=_killm_common_T_1|~mem_reg_valid; 
  assign _ctrl_killm_T=killm_common|mem_xcpt; 
  assign ctrl_killm=_ctrl_killm_T|fpu_kill_mem; 
  assign _wb_reg_wdata_T_1=~mem_reg_xcpt&mem_ctrl_fp; 
  assign _wb_reg_wdata_T_2=_wb_reg_wdata_T_1&mem_ctrl_wxd; 
  assign _T_100=_T_92 ? 3'h7:3'h5; 
  assign _T_101=_T_90 ? 4'hd:{1'b0,_T_100}; 
  assign _T_102=_T_88 ? 4'hf:_T_101; 
  assign _T_103=_T_86 ? 4'h4:_T_102; 
  assign _T_104=_T_84 ? 4'h6:_T_103; 
  assign wb_cause=wb_reg_xcpt ? wb_reg_cause:{60'b0,_T_104}; 
  assign _T_105=wb_cause==64'h6; 
  assign _T_107=wb_cause==64'h4; 
  assign _T_109=wb_cause==64'h7; 
  assign _T_111=wb_cause==64'h5; 
  assign _T_113=wb_cause==64'hf; 
  assign _T_115=wb_cause==64'hd; 
  assign _csr_io_inst_0_T_1=&wb_reg_raw_inst[1:0]; 
  assign csr_io_inst_0_hi=_csr_io_inst_0_T_1 ? wb_reg_inst[31:16]:16'h0; 
  assign csr_io_inst_0_lo=wb_reg_raw_inst[15:0]; 
  assign _tval_valid_T=wb_cause==64'h2; 
  assign _tval_valid_T_1=wb_cause==64'h3; 
  assign _tval_valid_T_6=wb_cause==64'h1; 
  assign _tval_valid_T_9=wb_cause==64'hc; 
  assign _tval_valid_T_10=_tval_valid_T|_tval_valid_T_1; 
  assign _tval_valid_T_11=_tval_valid_T_10|_T_107; 
  assign _tval_valid_T_12=_tval_valid_T_11|_T_105; 
  assign _tval_valid_T_13=_tval_valid_T_12|_T_111; 
  assign _tval_valid_T_14=_tval_valid_T_13|_T_109; 
  assign _tval_valid_T_15=_tval_valid_T_14|_tval_valid_T_6; 
  assign _tval_valid_T_16=_tval_valid_T_15|_T_115; 
  assign _tval_valid_T_17=_tval_valid_T_16|_T_113; 
  assign _tval_valid_T_18=_tval_valid_T_17|_tval_valid_T_9; 
  assign tval_valid=wb_xcpt&_tval_valid_T_18; 
  assign a_1=wb_reg_wdata[63:39]; 
  assign _csr_io_tval_msb_T=$signed(a_1)==25'sh0; 
  assign _csr_io_tval_msb_T_1=$signed(a_1)==-25'sh1; 
  assign _csr_io_tval_msb_T_2=_csr_io_tval_msb_T|_csr_io_tval_msb_T_1; 
  assign msb_1=_csr_io_tval_msb_T_2 ? wb_reg_wdata[39]:~wb_reg_wdata[38]; 
  assign csr_io_tval_lo=wb_reg_wdata[38:0]; 
  assign _csr_io_tval_T={msb_1,csr_io_tval_lo}; 
  assign _csr_io_rw_cmd_T=wb_reg_valid ? 3'h0:3'h4; 
  assign _T_129=32'h1<<ll_waddr; 
  assign _T_130=ll_wen ? _T_129:32'h0; 
  assign _T_132=r&~_T_130; 
  assign _T_134=wb_set_sboard&wb_wen; 
  assign _T_135=32'h1<<wb_waddr; 
  assign _T_136=_T_134 ? _T_135:32'h0; 
  assign _T_137=_T_132|_T_136; 
  assign _T_138=ll_wen|_T_134; 
  assign _id_stall_fpu_T=wb_dcache_miss&wb_ctrl_wfd; 
  assign _id_stall_fpu_T_1=_id_stall_fpu_T|io_fpu_sboard_set; 
  assign _id_stall_fpu_T_2=_id_stall_fpu_T_1&wb_valid; 
  assign _id_stall_fpu_T_4=_id_stall_fpu_T_2 ? _T_135:32'h0; 
  assign _id_stall_fpu_T_5=id_stall_fpu__r|_id_stall_fpu_T_4; 
  assign _id_stall_fpu_T_7=dmem_resp_replay&io_dmem_resp_bits_tag[0]; 
  assign _id_stall_fpu_T_8=32'h1<<dmem_resp_waddr; 
  assign _id_stall_fpu_T_9=_id_stall_fpu_T_7 ? _id_stall_fpu_T_8:32'h0; 
  assign _id_stall_fpu_T_11=_id_stall_fpu_T_5&~_id_stall_fpu_T_9; 
  assign _id_stall_fpu_T_12=_id_stall_fpu_T_2|_id_stall_fpu_T_7; 
  assign _id_stall_fpu_T_13=32'h1<<io_fpu_sboard_clra; 
  assign _id_stall_fpu_T_14=io_fpu_sboard_clr ? _id_stall_fpu_T_13:32'h0; 
  assign _id_stall_fpu_T_16=_id_stall_fpu_T_11&~_id_stall_fpu_T_14; 
  assign _id_stall_fpu_T_17=_id_stall_fpu_T_12|io_fpu_sboard_clr; 
  assign _dcache_blocked_blocked_T_3=~io_dmem_req_ready&~io_dmem_perf_grant; 
  assign _dcache_blocked_blocked_T_4=blocked|io_dmem_req_valid; 
  assign _dcache_blocked_blocked_T_5=_dcache_blocked_blocked_T_4|io_dmem_s2_nack; 
  assign _io_imem_req_bits_pc_T=wb_xcpt|csr_io_eret; 
  assign _io_imem_req_bits_pc_T_1=replay_wb_common ? wb_reg_pc:mem_npc; 
  assign _io_imem_flush_icache_T=wb_reg_valid&wb_ctrl_fence_i; 
  assign _io_imem_might_request_imem_might_request_reg_T=ex_pc_valid|mem_pc_valid; 
  assign _io_imem_btb_update_valid_T_1=mem_reg_valid&~take_pc_wb; 
  assign _io_imem_btb_update_valid_T_2=_io_imem_btb_update_valid_T_1&mem_wrong_npc; 
  assign _io_imem_btb_update_valid_T_4=~mem_cfi|mem_cfi_taken; 
  assign _io_imem_btb_update_bits_cfiType_T=mem_ctrl_jal|mem_ctrl_jalr; 
  assign _io_imem_btb_update_bits_cfiType_T_2=_io_imem_btb_update_bits_cfiType_T&mem_waddr[0]; 
  assign _io_imem_btb_update_bits_cfiType_T_5=mem_reg_inst[19:15]&5'h1b; 
  assign _io_imem_btb_update_bits_cfiType_T_6=5'h1==_io_imem_btb_update_bits_cfiType_T_5; 
  assign _io_imem_btb_update_bits_cfiType_T_7=mem_ctrl_jalr&_io_imem_btb_update_bits_cfiType_T_6; 
  assign _io_imem_btb_update_bits_cfiType_T_10=_io_imem_btb_update_bits_cfiType_T_7 ? 2'h3:{1'b0,_io_imem_btb_update_bits_cfiType_T}; 
  assign _io_imem_btb_update_bits_br_pc_T=mem_reg_rvc ? 2'h0:2'h2; 
  assign _GEN_250={38'b0,_io_imem_btb_update_bits_br_pc_T}; 
  assign _io_imem_btb_update_bits_br_pc_T_2=mem_reg_pc+_GEN_250; 
  assign _io_imem_btb_update_bits_pc_T_1=~io_imem_btb_update_bits_br_pc|39'h3; 
  assign ex_dcache_tag={ex_waddr,ex_ctrl_fp}; 
  assign a_2=_ex_op1_T[63:39]; 
  assign _io_dmem_req_bits_addr_msb_T=$signed(a_2)==25'sh0; 
  assign _io_dmem_req_bits_addr_msb_T_1=$signed(a_2)==-25'sh1; 
  assign _io_dmem_req_bits_addr_msb_T_2=_io_dmem_req_bits_addr_msb_T|_io_dmem_req_bits_addr_msb_T_1; 
  assign msb_2=_io_dmem_req_bits_addr_msb_T_2 ? alu_io_adder_out[39]:~alu_io_adder_out[38]; 
  assign io_dmem_req_bits_addr_lo=alu_io_adder_out[38:0]; 
  assign _io_dmem_s1_kill_T=killm_common|mem_ldst_xcpt; 
  assign _unpause_T_1=csr_io_time[4:0]==5'h0; 
  assign _unpause_T_2=_unpause_T_1|csr_io_inhibit_cycle; 
  assign _unpause_T_3=_unpause_T_2|io_dmem_perf_release; 
  assign unpause=_unpause_T_3|take_pc_mem_wb; 
   reg reg_coreMonitorBundle_valid ;  
  assign reg_coreMonitorBundle_valid=coreMonitorBundle_valid; 
  assign coreMonitorBundle_valid=csr_io_trace_0_valid&~csr_io_trace_0_exception; 
  assign coreMonitorBundle_wrenx=wb_wen&~wb_set_sboard; 
  assign _GEN_251={1'b0,wb_waddr}; 
  assign _T_142=_GEN_251+6'h20; 
  assign _T_145=wb_waddr!=5'h0; 
  assign _T_146=wb_ctrl_wxd&_T_145; 
  assign _T_147=_T_146&coreMonitorBundle_wrenx; 
  assign _T_153=_T_146&~coreMonitorBundle_wrenx; 
  assign _T_159=ll_wen&_T_118; 
  assign io_imem_might_request=imem_might_request_reg; 
  assign io_imem_req_valid=take_pc_wb|take_pc_mem; 
  assign io_imem_req_bits_pc=_io_imem_req_bits_pc_T ? csr_io_evec:_io_imem_req_bits_pc_T_1; 
  assign io_imem_req_bits_speculative=~take_pc_wb; 
  assign io_imem_sfence_valid=wb_reg_valid&wb_reg_sfence; 
  assign io_imem_sfence_bits_rs1=wb_reg_mem_size[0]; 
  assign io_imem_sfence_bits_rs2=wb_reg_mem_size[1]; 
  assign io_imem_sfence_bits_addr=wb_reg_wdata[38:0]; 
  assign io_imem_resp_ready=ibuf_io_imem_ready; 
  assign io_imem_btb_update_valid=_io_imem_btb_update_valid_T_2&_io_imem_btb_update_valid_T_4; 
  assign io_imem_btb_update_bits_prediction_entry=mem_reg_btb_resp_entry; 
  assign io_imem_btb_update_bits_pc=~_io_imem_btb_update_bits_pc_T_1; 
  assign io_imem_btb_update_bits_isValid=_mem_cfi_T|mem_ctrl_jal; 
  assign io_imem_btb_update_bits_br_pc=_io_imem_btb_update_bits_br_pc_T_2[38:0]; 
  assign io_imem_btb_update_bits_cfiType=_io_imem_btb_update_bits_cfiType_T_2 ? 2'h2:_io_imem_btb_update_bits_cfiType_T_10; 
  assign io_imem_bht_update_valid=mem_reg_valid&~take_pc_wb; 
  assign io_imem_bht_update_bits_prediction_history=mem_reg_btb_resp_bht_history; 
  assign io_imem_bht_update_bits_pc=io_imem_btb_update_bits_pc; 
  assign io_imem_bht_update_bits_branch=mem_ctrl_branch; 
  assign io_imem_bht_update_bits_taken=mem_br_taken; 
  assign io_imem_bht_update_bits_mispredict=ex_pc_valid ? _mem_wrong_npc_T:_mem_wrong_npc_T_3; 
  assign io_imem_flush_icache=_io_imem_flush_icache_T&~io_dmem_s2_nack; 
  assign io_dmem_req_valid=ex_reg_valid&ex_ctrl_mem; 
  assign io_dmem_req_bits_addr={msb_2,io_dmem_req_bits_addr_lo}; 
  assign io_dmem_req_bits_tag={1'b0,ex_dcache_tag}; 
  assign io_dmem_req_bits_cmd=ex_ctrl_mem_cmd; 
  assign io_dmem_req_bits_size=ex_reg_mem_size; 
  assign io_dmem_req_bits_signed=~ex_reg_inst[14]; 
  assign io_dmem_s1_kill=_io_dmem_s1_kill_T|fpu_kill_mem; 
  assign io_dmem_s1_data_data=mem_ctrl_fp ? io_fpu_store_data:mem_reg_rs2; 
  assign io_ptw_ptbr_mode=csr_io_ptbr_mode; 
  assign io_ptw_ptbr_ppn=csr_io_ptbr_ppn; 
  assign io_ptw_sfence_valid=io_imem_sfence_valid; 
  assign io_ptw_sfence_bits_rs1=io_imem_sfence_bits_rs1; 
  assign io_ptw_status_debug=csr_io_status_debug; 
  assign io_ptw_status_dprv=csr_io_status_dprv; 
  assign io_ptw_status_prv=csr_io_status_prv; 
  assign io_ptw_status_mxr=csr_io_status_mxr; 
  assign io_ptw_status_sum=csr_io_status_sum; 
  assign io_ptw_pmp_0_cfg_l=csr_io_pmp_0_cfg_l; 
  assign io_ptw_pmp_0_cfg_a=csr_io_pmp_0_cfg_a; 
  assign io_ptw_pmp_0_cfg_x=csr_io_pmp_0_cfg_x; 
  assign io_ptw_pmp_0_cfg_w=csr_io_pmp_0_cfg_w; 
  assign io_ptw_pmp_0_cfg_r=csr_io_pmp_0_cfg_r; 
  assign io_ptw_pmp_0_addr=csr_io_pmp_0_addr; 
  assign io_ptw_pmp_0_mask=csr_io_pmp_0_mask; 
  assign io_ptw_pmp_1_cfg_l=csr_io_pmp_1_cfg_l; 
  assign io_ptw_pmp_1_cfg_a=csr_io_pmp_1_cfg_a; 
  assign io_ptw_pmp_1_cfg_x=csr_io_pmp_1_cfg_x; 
  assign io_ptw_pmp_1_cfg_w=csr_io_pmp_1_cfg_w; 
  assign io_ptw_pmp_1_cfg_r=csr_io_pmp_1_cfg_r; 
  assign io_ptw_pmp_1_addr=csr_io_pmp_1_addr; 
  assign io_ptw_pmp_1_mask=csr_io_pmp_1_mask; 
  assign io_ptw_pmp_2_cfg_l=csr_io_pmp_2_cfg_l; 
  assign io_ptw_pmp_2_cfg_a=csr_io_pmp_2_cfg_a; 
  assign io_ptw_pmp_2_cfg_x=csr_io_pmp_2_cfg_x; 
  assign io_ptw_pmp_2_cfg_w=csr_io_pmp_2_cfg_w; 
  assign io_ptw_pmp_2_cfg_r=csr_io_pmp_2_cfg_r; 
  assign io_ptw_pmp_2_addr=csr_io_pmp_2_addr; 
  assign io_ptw_pmp_2_mask=csr_io_pmp_2_mask; 
  assign io_ptw_pmp_3_cfg_l=csr_io_pmp_3_cfg_l; 
  assign io_ptw_pmp_3_cfg_a=csr_io_pmp_3_cfg_a; 
  assign io_ptw_pmp_3_cfg_x=csr_io_pmp_3_cfg_x; 
  assign io_ptw_pmp_3_cfg_w=csr_io_pmp_3_cfg_w; 
  assign io_ptw_pmp_3_cfg_r=csr_io_pmp_3_cfg_r; 
  assign io_ptw_pmp_3_addr=csr_io_pmp_3_addr; 
  assign io_ptw_pmp_3_mask=csr_io_pmp_3_mask; 
  assign io_ptw_pmp_4_cfg_l=csr_io_pmp_4_cfg_l; 
  assign io_ptw_pmp_4_cfg_a=csr_io_pmp_4_cfg_a; 
  assign io_ptw_pmp_4_cfg_x=csr_io_pmp_4_cfg_x; 
  assign io_ptw_pmp_4_cfg_w=csr_io_pmp_4_cfg_w; 
  assign io_ptw_pmp_4_cfg_r=csr_io_pmp_4_cfg_r; 
  assign io_ptw_pmp_4_addr=csr_io_pmp_4_addr; 
  assign io_ptw_pmp_4_mask=csr_io_pmp_4_mask; 
  assign io_ptw_pmp_5_cfg_l=csr_io_pmp_5_cfg_l; 
  assign io_ptw_pmp_5_cfg_a=csr_io_pmp_5_cfg_a; 
  assign io_ptw_pmp_5_cfg_x=csr_io_pmp_5_cfg_x; 
  assign io_ptw_pmp_5_cfg_w=csr_io_pmp_5_cfg_w; 
  assign io_ptw_pmp_5_cfg_r=csr_io_pmp_5_cfg_r; 
  assign io_ptw_pmp_5_addr=csr_io_pmp_5_addr; 
  assign io_ptw_pmp_5_mask=csr_io_pmp_5_mask; 
  assign io_ptw_pmp_6_cfg_l=csr_io_pmp_6_cfg_l; 
  assign io_ptw_pmp_6_cfg_a=csr_io_pmp_6_cfg_a; 
  assign io_ptw_pmp_6_cfg_x=csr_io_pmp_6_cfg_x; 
  assign io_ptw_pmp_6_cfg_w=csr_io_pmp_6_cfg_w; 
  assign io_ptw_pmp_6_cfg_r=csr_io_pmp_6_cfg_r; 
  assign io_ptw_pmp_6_addr=csr_io_pmp_6_addr; 
  assign io_ptw_pmp_6_mask=csr_io_pmp_6_mask; 
  assign io_ptw_pmp_7_cfg_l=csr_io_pmp_7_cfg_l; 
  assign io_ptw_pmp_7_cfg_a=csr_io_pmp_7_cfg_a; 
  assign io_ptw_pmp_7_cfg_x=csr_io_pmp_7_cfg_x; 
  assign io_ptw_pmp_7_cfg_w=csr_io_pmp_7_cfg_w; 
  assign io_ptw_pmp_7_cfg_r=csr_io_pmp_7_cfg_r; 
  assign io_ptw_pmp_7_addr=csr_io_pmp_7_addr; 
  assign io_ptw_pmp_7_mask=csr_io_pmp_7_mask; 
  assign io_ptw_customCSRs_csrs_0_value=csr_io_customCSRs_0_value; 
  assign io_fpu_inst=ibuf_io_inst_0_bits_inst_bits; 
  assign io_fpu_fromint_data=ex_reg_rs_bypass_0 ? _ex_rs_T_5:_ex_rs_T_6; 
  assign io_fpu_fcsr_rm=csr_io_fcsr_rm; 
  assign io_fpu_dmem_resp_val=dmem_resp_valid&io_dmem_resp_bits_tag[0]; 
  assign io_fpu_dmem_resp_type={1'b0,io_dmem_resp_bits_size}; 
  assign io_fpu_dmem_resp_tag=io_dmem_resp_bits_tag[5:1]; 
  assign io_fpu_dmem_resp_data=io_dmem_resp_bits_data_word_bypass; 
  assign io_fpu_valid=~ctrl_killd&id_ctrl_decoder_1; 
  assign io_fpu_killx=_ctrl_killx_T|~ex_reg_valid; 
  assign io_fpu_killm=_killm_common_T_1|~mem_reg_valid; 
  assign io_trace_0_valid=csr_io_trace_0_valid; 
  assign io_trace_0_iaddr=csr_io_trace_0_iaddr; 
  assign io_trace_0_insn=csr_io_trace_0_insn; 
  assign io_trace_0_priv=csr_io_trace_0_priv; 
  assign io_trace_0_exception=csr_io_trace_0_exception; 
  assign io_trace_0_interrupt=csr_io_trace_0_interrupt; 
  assign io_trace_0_cause=csr_io_trace_0_cause; 
  assign io_trace_0_tval=csr_io_trace_0_tval; 
  assign io_wfi=csr_io_status_wfi; 
  assign ibuf_clock=clock; 
  assign ibuf_reset=reset; 
  assign ibuf_io_imem_valid=io_imem_resp_valid; 
  assign ibuf_io_imem_bits_btb_taken=io_imem_resp_bits_btb_taken; 
  assign ibuf_io_imem_bits_btb_bridx=io_imem_resp_bits_btb_bridx; 
  assign ibuf_io_imem_bits_btb_entry=io_imem_resp_bits_btb_entry; 
  assign ibuf_io_imem_bits_btb_bht_history=io_imem_resp_bits_btb_bht_history; 
  assign ibuf_io_imem_bits_pc=io_imem_resp_bits_pc; 
  assign ibuf_io_imem_bits_data=io_imem_resp_bits_data; 
  assign ibuf_io_imem_bits_xcpt_pf_inst=io_imem_resp_bits_xcpt_pf_inst; 
  assign ibuf_io_imem_bits_xcpt_ae_inst=io_imem_resp_bits_xcpt_ae_inst; 
  assign ibuf_io_imem_bits_replay=io_imem_resp_bits_replay; 
  assign ibuf_io_kill=take_pc_wb|take_pc_mem; 
  assign ibuf_io_inst_0_ready=~ctrl_stalld; 
  assign csr_clock=clock; 
  assign csr_reset=reset; 
  assign csr_io_ungated_clock=clock; 
  assign csr_io_interrupts_debug=io_interrupts_debug; 
  assign csr_io_interrupts_mtip=io_interrupts_mtip; 
  assign csr_io_interrupts_msip=io_interrupts_msip; 
  assign csr_io_interrupts_meip=io_interrupts_meip; 
  assign csr_io_interrupts_seip=io_interrupts_seip; 
  assign csr_io_hartid=io_hartid; 
  assign csr_io_rw_addr=wb_reg_inst[31:20]; 
  assign csr_io_rw_cmd=wb_ctrl_csr&~_csr_io_rw_cmd_T; 
  assign csr_io_rw_wdata=wb_reg_wdata; 
  assign csr_io_decode_0_csr=ibuf_io_inst_0_bits_raw[31:20]; 
  assign csr_io_exception=_T_99|_T_94; 
  assign csr_io_retire=_wb_valid_T_1&~wb_xcpt; 
  assign csr_io_cause=wb_reg_xcpt ? wb_reg_cause:{60'b0,_T_104}; 
  assign csr_io_pc=wb_reg_pc; 
  assign csr_io_tval=tval_valid ? _csr_io_tval_T:40'h0; 
  assign csr_io_fcsr_flags_valid=io_fpu_fcsr_flags_valid; 
  assign csr_io_fcsr_flags_bits=io_fpu_fcsr_flags_bits; 
  assign csr_io_inst_0={csr_io_inst_0_hi,csr_io_inst_0_lo}; 
  assign bpu_io_status_debug=csr_io_status_debug; 
  assign bpu_io_status_prv=csr_io_status_prv; 
  assign bpu_io_bp_0_control_action=csr_io_bp_0_control_action; 
  assign bpu_io_bp_0_control_tmatch=csr_io_bp_0_control_tmatch; 
  assign bpu_io_bp_0_control_m=csr_io_bp_0_control_m; 
  assign bpu_io_bp_0_control_s=csr_io_bp_0_control_s; 
  assign bpu_io_bp_0_control_u=csr_io_bp_0_control_u; 
  assign bpu_io_bp_0_control_x=csr_io_bp_0_control_x; 
  assign bpu_io_bp_0_control_w=csr_io_bp_0_control_w; 
  assign bpu_io_bp_0_control_r=csr_io_bp_0_control_r; 
  assign bpu_io_bp_0_address=csr_io_bp_0_address; 
  assign bpu_io_pc=ibuf_io_pc[38:0]; 
  assign bpu_io_ea=mem_reg_wdata[38:0]; 
  assign alu_io_dw=ex_ctrl_alu_dw; 
  assign alu_io_fn=ex_ctrl_alu_fn; 
  assign alu_io_in2=_ex_op2_T_6 ? $signed({{60{_ex_op2_T_1[3]}},_ex_op2_T_1}):$signed(_ex_op2_T_5); 
  assign alu_io_in1=_ex_op1_T_4 ? $signed({{24{ex_reg_pc[39]}},ex_reg_pc}):$signed(_ex_op1_T_3); 
  assign div_clock=clock; 
  assign div_reset=reset; 
  assign div_io_req_valid=ex_reg_valid&ex_ctrl_div; 
  assign div_io_req_bits_fn=ex_ctrl_alu_fn; 
  assign div_io_req_bits_dw=ex_ctrl_alu_dw; 
  assign div_io_req_bits_in1=ex_reg_rs_bypass_0 ? _ex_rs_T_5:_ex_rs_T_6; 
  assign div_io_req_bits_in2=ex_reg_rs_bypass_1 ? _ex_rs_T_12:_ex_rs_T_13; 
  assign div_io_req_bits_tag=ex_reg_inst[11:7]; 
  assign div_io_kill=killm_common&div_io_kill_REG; 
  assign div_io_resp_ready=_T_117 ? 1'h0:~wb_wxd; 
  assign PlusArgTimeout_clock=clock; 
  assign PlusArgTimeout_reset=reset; 
  assign PlusArgTimeout_io_count=csr_io_time[31:0]; 
  assign _GEN_254=coreMonitorBundle_valid&wb_ctrl_wfd; 
  assign _GEN_256=coreMonitorBundle_valid&~wb_ctrl_wfd; 
  assign _GEN_257=_GEN_256&_T_147; 
  assign _GEN_261=_GEN_256&~_T_147; 
  assign _GEN_262=_GEN_261&_T_153; 
  assign _GEN_268=_GEN_261&~_T_153; 
  assign Rocket_cov_read_addr=Rocket_state; 
  assign Rocket_cov_read_data=Rocket_cov[Rocket_cov_read_addr]; 
  assign Rocket_cov_write_data=1'h1; 
  assign Rocket_cov_write_addr=Rocket_state; 
  assign Rocket_cov_write_mask=1'h1; 
  assign Rocket_cov_write_en=1'h1; 
  assign mux_cond_0=_T_122; 
  assign mux_cond_1=_csr_io_tval_msb_T_2; 
  assign mux_cond_2=_mem_npc_msb_T_2; 
  assign mux_cond_3=_csr_io_inst_0_T_1; 
  assign mux_cond_4=_T_118; 
  assign mux_cond_5=_T_121; 
  assign ex_ctrl_wfd_shl={ex_ctrl_wfd,10'h0}; 
  assign ex_ctrl_wfd_pad={9'h0,ex_ctrl_wfd_shl}; 
  assign ex_ctrl_fp_shl={ex_ctrl_fp,15'h0}; 
  assign ex_ctrl_fp_pad={4'h0,ex_ctrl_fp_shl}; 
  assign mem_ctrl_jalr_shl={mem_ctrl_jalr,15'h0}; 
  assign mem_ctrl_jalr_pad={4'h0,mem_ctrl_jalr_shl}; 
  assign wb_ctrl_mem_shl={wb_ctrl_mem,11'h0}; 
  assign wb_ctrl_mem_pad={8'h0,wb_ctrl_mem_shl}; 
  assign ex_ctrl_wxd_shl={ex_ctrl_wxd,6'h0}; 
  assign ex_ctrl_wxd_pad={13'h0,ex_ctrl_wxd_shl}; 
  assign ex_ctrl_mem_shl={ex_ctrl_mem,19'h0}; 
  assign ex_ctrl_mem_pad=ex_ctrl_mem_shl; 
  assign ex_ctrl_sel_alu1_shl={ex_ctrl_sel_alu1,18'h0}; 
  assign ex_ctrl_sel_alu1_pad=ex_ctrl_sel_alu1_shl; 
  assign mem_reg_replay_shl={mem_reg_replay,11'h0}; 
  assign mem_reg_replay_pad={8'h0,mem_reg_replay_shl}; 
  assign blocked_shl={blocked,16'h0}; 
  assign blocked_pad={3'h0,blocked_shl}; 
  assign wb_ctrl_div_shl={wb_ctrl_div,2'h0}; 
  assign wb_ctrl_div_pad={17'h0,wb_ctrl_div_shl}; 
  assign wb_reg_flush_pipe_shl={wb_reg_flush_pipe,15'h0}; 
  assign wb_reg_flush_pipe_pad={4'h0,wb_reg_flush_pipe_shl}; 
  assign mem_ctrl_jal_shl={mem_ctrl_jal,11'h0}; 
  assign mem_ctrl_jal_pad={8'h0,mem_ctrl_jal_shl}; 
  assign ex_ctrl_sel_imm_shl={ex_ctrl_sel_imm,7'h0}; 
  assign ex_ctrl_sel_imm_pad={10'h0,ex_ctrl_sel_imm_shl}; 
  assign wb_ctrl_wfd_shl={wb_ctrl_wfd,8'h0}; 
  assign wb_ctrl_wfd_pad={11'h0,wb_ctrl_wfd_shl}; 
  assign mem_reg_slow_bypass_shl={mem_reg_slow_bypass,19'h0}; 
  assign mem_reg_slow_bypass_pad=mem_reg_slow_bypass_shl; 
  assign mem_reg_sfence_shl={mem_reg_sfence,16'h0}; 
  assign mem_reg_sfence_pad={3'h0,mem_reg_sfence_shl}; 
  assign wb_reg_xcpt_shl={wb_reg_xcpt,2'h0}; 
  assign wb_reg_xcpt_pad={17'h0,wb_reg_xcpt_shl}; 
  assign id_reg_pause_shl={id_reg_pause,15'h0}; 
  assign id_reg_pause_pad={4'h0,id_reg_pause_shl}; 
  assign ex_reg_rvc_shl={ex_reg_rvc,8'h0}; 
  assign ex_reg_rvc_pad={11'h0,ex_reg_rvc_shl}; 
  assign wb_reg_valid_shl={wb_reg_valid,3'h0}; 
  assign wb_reg_valid_pad={16'h0,wb_reg_valid_shl}; 
  assign mem_br_taken_shl={mem_br_taken,13'h0}; 
  assign mem_br_taken_pad={6'h0,mem_br_taken_shl}; 
  assign mem_reg_flush_pipe_shl={mem_reg_flush_pipe,18'h0}; 
  assign mem_reg_flush_pipe_pad={1'h0,mem_reg_flush_pipe_shl}; 
  assign ex_ctrl_div_shl={ex_ctrl_div,17'h0}; 
  assign ex_ctrl_div_pad={2'h0,ex_ctrl_div_shl}; 
  assign mem_ctrl_fp_shl={mem_ctrl_fp,15'h0}; 
  assign mem_ctrl_fp_pad={4'h0,mem_ctrl_fp_shl}; 
  assign mem_reg_xcpt_shl={mem_reg_xcpt,5'h0}; 
  assign mem_reg_xcpt_pad={14'h0,mem_reg_xcpt_shl}; 
  assign mem_ctrl_wxd_shl={mem_ctrl_wxd,14'h0}; 
  assign mem_ctrl_wxd_pad={5'h0,mem_ctrl_wxd_shl}; 
  assign mem_ctrl_mem_shl={mem_ctrl_mem,8'h0}; 
  assign mem_ctrl_mem_pad={11'h0,mem_ctrl_mem_shl}; 
  assign ex_reg_mem_size_shl={ex_reg_mem_size,15'h0}; 
  assign ex_reg_mem_size_pad={3'h0,ex_reg_mem_size_shl}; 
  assign ex_ctrl_sel_alu2_shl={ex_ctrl_sel_alu2,7'h0}; 
  assign ex_ctrl_sel_alu2_pad={11'h0,ex_ctrl_sel_alu2_shl}; 
  assign ex_ctrl_rxs2_shl={ex_ctrl_rxs2,2'h0}; 
  assign ex_ctrl_rxs2_pad={17'h0,ex_ctrl_rxs2_shl}; 
  assign ex_ctrl_jalr_shl={ex_ctrl_jalr,3'h0}; 
  assign ex_ctrl_jalr_pad={16'h0,ex_ctrl_jalr_shl}; 
  assign ex_reg_replay_shl={ex_reg_replay,4'h0}; 
  assign ex_reg_replay_pad={15'h0,ex_reg_replay_shl}; 
  assign ex_reg_valid_shl={ex_reg_valid,3'h0}; 
  assign ex_reg_valid_pad={16'h0,ex_reg_valid_shl}; 
  assign mem_reg_valid_shl={mem_reg_valid,6'h0}; 
  assign mem_reg_valid_pad={13'h0,mem_reg_valid_shl}; 
  assign mem_reg_rvc_shl=mem_reg_rvc; 
  assign mem_reg_rvc_pad={19'h0,mem_reg_rvc_shl}; 
  assign mem_ctrl_wfd_shl=mem_ctrl_wfd; 
  assign mem_ctrl_wfd_pad={19'h0,mem_ctrl_wfd_shl}; 
  assign id_reg_fence_shl={id_reg_fence,11'h0}; 
  assign id_reg_fence_pad={8'h0,id_reg_fence_shl}; 
  assign mem_reg_load_shl={mem_reg_load,8'h0}; 
  assign mem_reg_load_pad={11'h0,mem_reg_load_shl}; 
  assign wb_ctrl_wxd_shl={wb_ctrl_wxd,18'h0}; 
  assign wb_ctrl_wxd_pad={1'h0,wb_ctrl_wxd_shl}; 
  assign wb_reg_replay_shl={wb_reg_replay,1'h0}; 
  assign wb_reg_replay_pad={18'h0,wb_reg_replay_shl}; 
  assign ex_reg_xcpt_interrupt_shl={ex_reg_xcpt_interrupt,10'h0}; 
  assign ex_reg_xcpt_interrupt_pad={9'h0,ex_reg_xcpt_interrupt_shl}; 
  assign mem_ctrl_branch_shl={mem_ctrl_branch,6'h0}; 
  assign mem_ctrl_branch_pad={13'h0,mem_ctrl_branch_shl}; 
  assign mem_reg_xcpt_interrupt_shl={mem_reg_xcpt_interrupt,1'h0}; 
  assign mem_reg_xcpt_interrupt_pad={18'h0,mem_reg_xcpt_interrupt_shl}; 
  assign mem_reg_store_shl={mem_reg_store,4'h0}; 
  assign mem_reg_store_pad={15'h0,mem_reg_store_shl}; 
  assign mem_ctrl_div_shl={mem_ctrl_div,5'h0}; 
  assign mem_ctrl_div_pad={14'h0,mem_ctrl_div_shl}; 
  assign mux_cond_0_shl={mux_cond_0,17'h0}; 
  assign mux_cond_0_pad={2'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,8'h0}; 
  assign mux_cond_1_pad={11'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl={mux_cond_2,15'h0}; 
  assign mux_cond_2_pad={4'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,4'h0}; 
  assign mux_cond_3_pad={15'h0,mux_cond_3_shl}; 
  assign mux_cond_4_shl={mux_cond_4,9'h0}; 
  assign mux_cond_4_pad={10'h0,mux_cond_4_shl}; 
  assign mux_cond_5_shl={mux_cond_5,17'h0}; 
  assign mux_cond_5_pad={2'h0,mux_cond_5_shl}; 
  assign ex_reg_rs_lsb_0_shl={ex_reg_rs_lsb_0,11'h0}; 
  assign ex_reg_rs_lsb_0_pad={7'h0,ex_reg_rs_lsb_0_shl}; 
  assign ex_reg_rs_lsb_1_shl={ex_reg_rs_lsb_1,11'h0}; 
  assign ex_reg_rs_lsb_1_pad={7'h0,ex_reg_rs_lsb_1_shl}; 
  assign ex_reg_rs_bypass_0_shl={ex_reg_rs_bypass_0,10'h0}; 
  assign ex_reg_rs_bypass_0_pad={9'h0,ex_reg_rs_bypass_0_shl}; 
  assign ex_reg_rs_bypass_1_shl={ex_reg_rs_bypass_1,10'h0}; 
  assign ex_reg_rs_bypass_1_pad={9'h0,ex_reg_rs_bypass_1_shl}; 
  assign Rocket_xor32=ex_ctrl_fp_pad^mem_ctrl_jalr_pad; 
  assign Rocket_xor15=ex_ctrl_wfd_pad^Rocket_xor32; 
  assign Rocket_xor34=ex_ctrl_wxd_pad^ex_ctrl_mem_pad; 
  assign Rocket_xor16=wb_ctrl_mem_pad^Rocket_xor34; 
  assign Rocket_xor7=Rocket_xor15^Rocket_xor16; 
  assign Rocket_xor36=mem_reg_replay_pad^blocked_pad; 
  assign Rocket_xor17=ex_ctrl_sel_alu1_pad^Rocket_xor36; 
  assign Rocket_xor37=wb_ctrl_div_pad^wb_reg_flush_pipe_pad; 
  assign Rocket_xor38=mem_ctrl_jal_pad^ex_ctrl_sel_imm_pad; 
  assign Rocket_xor18=Rocket_xor37^Rocket_xor38; 
  assign Rocket_xor8=Rocket_xor17^Rocket_xor18; 
  assign Rocket_xor3=Rocket_xor7^Rocket_xor8; 
  assign Rocket_xor40=mem_reg_slow_bypass_pad^mem_reg_sfence_pad; 
  assign Rocket_xor19=wb_ctrl_wfd_pad^Rocket_xor40; 
  assign Rocket_xor41=wb_reg_xcpt_pad^id_reg_pause_pad; 
  assign Rocket_xor42=ex_reg_rvc_pad^wb_reg_valid_pad; 
  assign Rocket_xor20=Rocket_xor41^Rocket_xor42; 
  assign Rocket_xor9=Rocket_xor19^Rocket_xor20; 
  assign Rocket_xor44=mem_reg_flush_pipe_pad^ex_ctrl_div_pad; 
  assign Rocket_xor21=mem_br_taken_pad^Rocket_xor44; 
  assign Rocket_xor45=mem_ctrl_fp_pad^mem_reg_xcpt_pad; 
  assign Rocket_xor46=mem_ctrl_wxd_pad^mem_ctrl_mem_pad; 
  assign Rocket_xor22=Rocket_xor45^Rocket_xor46; 
  assign Rocket_xor10=Rocket_xor21^Rocket_xor22; 
  assign Rocket_xor4=Rocket_xor9^Rocket_xor10; 
  assign Rocket_xor1=Rocket_xor3^Rocket_xor4; 
  assign Rocket_xor48=ex_ctrl_sel_alu2_pad^ex_ctrl_rxs2_pad; 
  assign Rocket_xor23=ex_reg_mem_size_pad^Rocket_xor48; 
  assign Rocket_xor49=ex_ctrl_jalr_pad^ex_reg_replay_pad; 
  assign Rocket_xor50=ex_reg_valid_pad^mem_reg_valid_pad; 
  assign Rocket_xor24=Rocket_xor49^Rocket_xor50; 
  assign Rocket_xor11=Rocket_xor23^Rocket_xor24; 
  assign Rocket_xor52=mem_ctrl_wfd_pad^id_reg_fence_pad; 
  assign Rocket_xor25=mem_reg_rvc_pad^Rocket_xor52; 
  assign Rocket_xor53=mem_reg_load_pad^wb_ctrl_wxd_pad; 
  assign Rocket_xor54=wb_reg_replay_pad^ex_reg_xcpt_interrupt_pad; 
  assign Rocket_xor26=Rocket_xor53^Rocket_xor54; 
  assign Rocket_xor12=Rocket_xor25^Rocket_xor26; 
  assign Rocket_xor5=Rocket_xor11^Rocket_xor12; 
  assign Rocket_xor56=mem_reg_xcpt_interrupt_pad^mem_reg_store_pad; 
  assign Rocket_xor27=mem_ctrl_branch_pad^Rocket_xor56; 
  assign Rocket_xor57=mem_ctrl_div_pad^mux_cond_0_pad; 
  assign Rocket_xor58=mux_cond_1_pad^mux_cond_2_pad; 
  assign Rocket_xor28=Rocket_xor57^Rocket_xor58; 
  assign Rocket_xor13=Rocket_xor27^Rocket_xor28; 
  assign Rocket_xor60=mux_cond_4_pad^mux_cond_5_pad; 
  assign Rocket_xor29=mux_cond_3_pad^Rocket_xor60; 
  assign Rocket_xor61=ex_reg_rs_lsb_0_pad^ex_reg_rs_lsb_1_pad; 
  assign Rocket_xor62=ex_reg_rs_bypass_0_pad^ex_reg_rs_bypass_1_pad; 
  assign Rocket_xor30=Rocket_xor61^Rocket_xor62; 
  assign Rocket_xor14=Rocket_xor29^Rocket_xor30; 
  assign Rocket_xor6=Rocket_xor13^Rocket_xor14; 
  assign Rocket_xor2=Rocket_xor5^Rocket_xor6; 
  assign Rocket_xor0=Rocket_xor1^Rocket_xor2; 
  assign PlusArgTimeout_sum=Rocket_covSum+PlusArgTimeout_io_covSum; 
  assign csr_sum=PlusArgTimeout_sum+csr_io_covSum; 
  assign bpu_sum=csr_sum+bpu_io_covSum; 
  assign ibuf_sum=bpu_sum+ibuf_io_covSum; 
  assign div_sum=ibuf_sum+div_io_covSum; 
  assign alu_sum=div_sum+alu_io_covSum; 
  assign io_covSum=alu_sum; 
  assign alu_metaAssert_wire=alu_metaAssert; 
  assign bpu_metaAssert_wire=bpu_metaAssert; 
  assign PlusArgTimeout_metaAssert_wire=PlusArgTimeout_metaAssert; 
  assign csr_metaAssert_wire=csr_metaAssert; 
  assign ibuf_metaAssert_wire=ibuf_metaAssert; 
  assign div_metaAssert_wire=div_metaAssert; 
  assign Rocket_or4=alu_metaAssert_wire|PlusArgTimeout_metaAssert_wire; 
  assign Rocket_or1=ibuf_metaAssert_wire|Rocket_or4; 
  assign Rocket_or6=div_metaAssert_wire|csr_metaAssert_wire; 
  assign Rocket_or2=bpu_metaAssert_wire|Rocket_or6; 
  assign Rocket_or0=Rocket_or1|Rocket_or2; 
  assign metaAssert=Rocket_metaAssert; 
  assign PlusArgTimeout_metaReset=metaReset|PlusArgTimeout_halt; 
  assign csr_metaReset=metaReset|csr_halt; 
  assign ibuf_metaReset=metaReset|ibuf_halt; 
  assign div_metaReset=metaReset|div_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (rf_MPORT_en&rf_MPORT_mask)
            begin 
              rf [rf_MPORT_addr]<=rf_MPORT_data;
            end 
         if (metaReset)
            begin 
              id_reg_pause <=1'h0;
            end 
          else 
            if (unpause)
               begin 
                 id_reg_pause <=1'h0;
               end 
             else 
               if (~ctrl_killd)
                  begin 
                    id_reg_pause <=_GEN_1;
                  end 
         if (metaReset)
            begin 
              imem_might_request_reg <=1'h0;
            end 
          else 
            begin 
              imem_might_request_reg <=_io_imem_might_request_imem_might_request_reg_T|io_ptw_customCSRs_csrs_0_value[1];
            end 
         if (metaReset)
            begin 
              ex_ctrl_fp <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_fp <=id_ctrl_decoder_1;
               end 
         if (metaReset)
            begin 
              ex_ctrl_branch <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_branch <=id_ctrl_decoder_3;
               end 
         if (metaReset)
            begin 
              ex_ctrl_jal <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_jal <=id_ctrl_decoder_4;
               end 
         if (metaReset)
            begin 
              ex_ctrl_jalr <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_jalr <=id_ctrl_decoder_5;
               end 
         if (metaReset)
            begin 
              ex_ctrl_rxs2 <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_rxs2 <=id_ctrl_decoder_6;
               end 
         if (metaReset)
            begin 
              ex_ctrl_sel_alu2 <=2'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_xcpt)
                    begin 
                      if (_T_35)
                         begin 
                           ex_ctrl_sel_alu2 <=2'h0;
                         end 
                       else 
                         if (_T_32)
                            begin 
                              ex_ctrl_sel_alu2 <=2'h1;
                            end 
                          else 
                            begin 
                              ex_ctrl_sel_alu2 <=2'h0;
                            end 
                    end 
                  else 
                    begin 
                      ex_ctrl_sel_alu2 <=id_ctrl_decoder_9;
                    end 
               end 
         if (metaReset)
            begin 
              ex_ctrl_sel_alu1 <=2'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_xcpt)
                    begin 
                      if (_T_35)
                         begin 
                           ex_ctrl_sel_alu1 <=2'h2;
                         end 
                       else 
                         if (_T_32)
                            begin 
                              ex_ctrl_sel_alu1 <=2'h2;
                            end 
                          else 
                            begin 
                              ex_ctrl_sel_alu1 <=2'h1;
                            end 
                    end 
                  else 
                    begin 
                      ex_ctrl_sel_alu1 <=id_ctrl_decoder_10;
                    end 
               end 
         if (metaReset)
            begin 
              ex_ctrl_sel_imm <=3'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_sel_imm <=id_ctrl_decoder_11;
               end 
         if (metaReset)
            begin 
              ex_ctrl_alu_dw <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_alu_dw <=_GEN_9;
               end 
         if (metaReset)
            begin 
              ex_ctrl_alu_fn <=4'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_xcpt)
                    begin 
                      ex_ctrl_alu_fn <=4'h0;
                    end 
                  else 
                    begin 
                      ex_ctrl_alu_fn <=id_ctrl_decoder_13;
                    end 
               end 
         if (metaReset)
            begin 
              ex_ctrl_mem <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_mem <=id_ctrl_decoder_14;
               end 
         if (metaReset)
            begin 
              ex_ctrl_mem_cmd <=5'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_mem_cmd <=id_ctrl_decoder_15;
               end 
         if (metaReset)
            begin 
              ex_ctrl_wfd <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_wfd <=id_ctrl_decoder_19;
               end 
         if (metaReset)
            begin 
              ex_ctrl_div <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_div <=id_ctrl_decoder_21;
               end 
         if (metaReset)
            begin 
              ex_ctrl_wxd <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_wxd <=id_ctrl_decoder_22;
               end 
         if (metaReset)
            begin 
              ex_ctrl_csr <=3'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_csr_ren)
                    begin 
                      ex_ctrl_csr <=3'h2;
                    end 
                  else 
                    begin 
                      ex_ctrl_csr <=id_ctrl_decoder_23;
                    end 
               end 
         if (metaReset)
            begin 
              ex_ctrl_fence_i <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_ctrl_fence_i <=id_ctrl_decoder_24;
               end 
         if (metaReset)
            begin 
              mem_ctrl_fp <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_fp <=ex_ctrl_fp;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_branch <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_branch <=ex_ctrl_branch;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_jal <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_jal <=ex_ctrl_jal;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_jalr <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_jalr <=ex_ctrl_jalr;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_mem <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_mem <=ex_ctrl_mem;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_wfd <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_wfd <=ex_ctrl_wfd;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_div <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_div <=ex_ctrl_div;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_wxd <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_wxd <=ex_ctrl_wxd;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_csr <=3'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_csr <=ex_ctrl_csr;
                    end 
               end 
         if (metaReset)
            begin 
              mem_ctrl_fence_i <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_ctrl_fence_i <=_GEN_77;
                    end 
               end 
         if (metaReset)
            begin 
              wb_ctrl_mem <=1'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_ctrl_mem <=mem_ctrl_mem;
               end 
         if (metaReset)
            begin 
              wb_ctrl_wfd <=1'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_ctrl_wfd <=mem_ctrl_wfd;
               end 
         if (metaReset)
            begin 
              wb_ctrl_div <=1'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_ctrl_div <=mem_ctrl_div;
               end 
         if (metaReset)
            begin 
              wb_ctrl_wxd <=1'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_ctrl_wxd <=mem_ctrl_wxd;
               end 
         if (metaReset)
            begin 
              wb_ctrl_csr <=3'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_ctrl_csr <=mem_ctrl_csr;
               end 
         if (metaReset)
            begin 
              wb_ctrl_fence_i <=1'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_ctrl_fence_i <=mem_ctrl_fence_i;
               end 
         if (metaReset)
            begin 
              ex_reg_xcpt_interrupt <=1'h0;
            end 
          else 
            begin 
              ex_reg_xcpt_interrupt <=_ex_reg_replay_T_1&csr_io_interrupt;
            end 
         if (metaReset)
            begin 
              ex_reg_valid <=1'h0;
            end 
          else 
            begin 
              ex_reg_valid <=~ctrl_killd;
            end 
         if (metaReset)
            begin 
              ex_reg_rvc <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_xcpt)
                    begin 
                      ex_reg_rvc <=_GEN_5;
                    end 
                  else 
                    begin 
                      ex_reg_rvc <=ibuf_io_inst_0_bits_rvc;
                    end 
               end 
         if (metaReset)
            begin 
              ex_reg_btb_resp_entry <=5'h0;
            end 
          else 
            if (_T_45)
               begin 
                 ex_reg_btb_resp_entry <=ibuf_io_btb_resp_entry;
               end 
         if (metaReset)
            begin 
              ex_reg_btb_resp_bht_history <=8'h0;
            end 
          else 
            if (_T_45)
               begin 
                 ex_reg_btb_resp_bht_history <=ibuf_io_btb_resp_bht_history;
               end 
         if (metaReset)
            begin 
              ex_reg_xcpt <=1'h0;
            end 
          else 
            begin 
              ex_reg_xcpt <=~ctrl_killd&id_xcpt;
            end 
         if (metaReset)
            begin 
              ex_reg_flush_pipe <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_reg_flush_pipe <=_ex_reg_flush_pipe_T;
               end 
         if (metaReset)
            begin 
              ex_reg_load_use <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_reg_load_use <=id_load_use;
               end 
         if (metaReset)
            begin 
              ex_reg_cause <=64'h0;
            end 
          else 
            if (_T_45)
               begin 
                 if (csr_io_interrupt)
                    begin 
                      ex_reg_cause <=csr_io_interrupt_cause;
                    end 
                  else 
                    begin 
                      ex_reg_cause <={60'b0,_T_12};
                    end 
               end 
         if (metaReset)
            begin 
              ex_reg_replay <=1'h0;
            end 
          else 
            begin 
              ex_reg_replay <=_ex_reg_replay_T_1&ibuf_io_inst_0_bits_replay;
            end 
         if (metaReset)
            begin 
              ex_reg_pc <=40'h0;
            end 
          else 
            if (_T_45)
               begin 
                 ex_reg_pc <=ibuf_io_pc;
               end 
         if (metaReset)
            begin 
              ex_reg_mem_size <=2'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (_T_38)
                    begin 
                      ex_reg_mem_size <=_ex_reg_mem_size_T_1;
                    end 
                  else 
                    begin 
                      ex_reg_mem_size <=ibuf_io_inst_0_bits_inst_bits[13:12];
                    end 
               end 
         if (metaReset)
            begin 
              ex_reg_inst <=32'h0;
            end 
          else 
            if (_T_45)
               begin 
                 ex_reg_inst <=ibuf_io_inst_0_bits_inst_bits;
               end 
         if (metaReset)
            begin 
              ex_reg_raw_inst <=32'h0;
            end 
          else 
            if (_T_45)
               begin 
                 ex_reg_raw_inst <=ibuf_io_inst_0_bits_raw;
               end 
         if (metaReset)
            begin 
              mem_reg_xcpt_interrupt <=1'h0;
            end 
          else 
            begin 
              mem_reg_xcpt_interrupt <=~take_pc_mem_wb&ex_reg_xcpt_interrupt;
            end 
         if (metaReset)
            begin 
              mem_reg_valid <=1'h0;
            end 
          else 
            begin 
              mem_reg_valid <=~ctrl_killx;
            end 
         if (metaReset)
            begin 
              mem_reg_rvc <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_rvc <=ex_reg_rvc;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_btb_resp_entry <=5'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_btb_resp_entry <=ex_reg_btb_resp_entry;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_btb_resp_bht_history <=8'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_btb_resp_bht_history <=ex_reg_btb_resp_bht_history;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_xcpt <=1'h0;
            end 
          else 
            begin 
              mem_reg_xcpt <=~ctrl_killx&ex_xcpt;
            end 
         if (metaReset)
            begin 
              mem_reg_replay <=1'h0;
            end 
          else 
            begin 
              mem_reg_replay <=~take_pc_mem_wb&replay_ex;
            end 
         if (metaReset)
            begin 
              mem_reg_flush_pipe <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_flush_pipe <=_GEN_78;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_cause <=64'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_cause <=ex_reg_cause;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_slow_bypass <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_slow_bypass <=ex_slow_bypass;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_load <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_load <=_mem_reg_load_T_23;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_store <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_store <=_mem_reg_store_T_23;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_sfence <=1'h0;
            end 
          else 
            if (_T_56)
               begin 
                 mem_reg_sfence <=1'h0;
               end 
             else 
               if (ex_pc_valid)
                  begin 
                    mem_reg_sfence <=ex_sfence;
                  end 
         if (metaReset)
            begin 
              mem_reg_pc <=40'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_pc <=ex_reg_pc;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_inst <=32'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_inst <=ex_reg_inst;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_mem_size <=2'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_mem_size <=ex_reg_mem_size;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_raw_inst <=32'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_raw_inst <=ex_reg_raw_inst;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_wdata <=64'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_reg_wdata <=_mem_reg_wdata_T;
                    end 
               end 
         if (metaReset)
            begin 
              mem_reg_rs2 <=64'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      if (_T_59)
                         begin 
                           if (_mem_reg_rs2_T)
                              begin 
                                mem_reg_rs2 <=_mem_reg_rs2_T_1;
                              end 
                            else 
                              if (_mem_reg_rs2_T_2)
                                 begin 
                                   mem_reg_rs2 <=_mem_reg_rs2_T_3;
                                 end 
                               else 
                                 if (_mem_reg_rs2_T_4)
                                    begin 
                                      mem_reg_rs2 <=_mem_reg_rs2_T_5;
                                    end 
                                  else 
                                    if (ex_reg_rs_bypass_1)
                                       begin 
                                         if (_ex_rs_T_11)
                                            begin 
                                              mem_reg_rs2 <=io_dmem_resp_bits_data_word_bypass;
                                            end 
                                          else 
                                            if (_ex_rs_T_9)
                                               begin 
                                                 mem_reg_rs2 <=wb_reg_wdata;
                                               end 
                                             else 
                                               if (_ex_rs_T_7)
                                                  begin 
                                                    mem_reg_rs2 <=mem_reg_wdata;
                                                  end 
                                                else 
                                                  begin 
                                                    mem_reg_rs2 <=64'h0;
                                                  end 
                                       end 
                                     else 
                                       begin 
                                         mem_reg_rs2 <=_ex_rs_T_13;
                                       end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              mem_br_taken <=1'h0;
            end 
          else 
            if (!(_T_56))
               begin 
                 if (ex_pc_valid)
                    begin 
                      mem_br_taken <=alu_io_cmp_out;
                    end 
               end 
         if (metaReset)
            begin 
              wb_reg_valid <=1'h0;
            end 
          else 
            begin 
              wb_reg_valid <=~ctrl_killm;
            end 
         if (metaReset)
            begin 
              wb_reg_xcpt <=1'h0;
            end 
          else 
            begin 
              wb_reg_xcpt <=mem_xcpt&~take_pc_wb;
            end 
         if (metaReset)
            begin 
              wb_reg_replay <=1'h0;
            end 
          else 
            begin 
              wb_reg_replay <=replay_mem&~take_pc_wb;
            end 
         if (metaReset)
            begin 
              wb_reg_flush_pipe <=1'h0;
            end 
          else 
            begin 
              wb_reg_flush_pipe <=~ctrl_killm&mem_reg_flush_pipe;
            end 
         if (metaReset)
            begin 
              wb_reg_cause <=64'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 if (_T_61)
                    begin 
                      wb_reg_cause <=mem_reg_cause;
                    end 
                  else 
                    begin 
                      wb_reg_cause <={60'b0,_T_65};
                    end 
               end 
         if (metaReset)
            begin 
              wb_reg_sfence <=1'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_reg_sfence <=mem_reg_sfence;
               end 
         if (metaReset)
            begin 
              wb_reg_pc <=40'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_reg_pc <=mem_reg_pc;
               end 
         if (metaReset)
            begin 
              wb_reg_mem_size <=2'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_reg_mem_size <=mem_reg_mem_size;
               end 
         if (metaReset)
            begin 
              wb_reg_inst <=32'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_reg_inst <=mem_reg_inst;
               end 
         if (metaReset)
            begin 
              wb_reg_raw_inst <=32'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 wb_reg_raw_inst <=mem_reg_raw_inst;
               end 
         if (metaReset)
            begin 
              wb_reg_wdata <=64'h0;
            end 
          else 
            if (mem_pc_valid)
               begin 
                 if (_wb_reg_wdata_T_2)
                    begin 
                      wb_reg_wdata <=io_fpu_toint_data;
                    end 
                  else 
                    begin 
                      wb_reg_wdata <=mem_int_wdata;
                    end 
               end 
         if (metaReset)
            begin 
              id_reg_fence <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 id_reg_fence <=1'h0;
               end 
             else 
               if (~ctrl_killd)
                  begin 
                    id_reg_fence <=_GEN_2;
                  end 
                else 
                  if (~id_mem_busy)
                     begin 
                       id_reg_fence <=1'h0;
                     end 
         if (metaReset)
            begin 
              ex_reg_rs_bypass_0 <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_illegal_insn)
                    begin 
                      ex_reg_rs_bypass_0 <=1'h0;
                    end 
                  else 
                    begin 
                      ex_reg_rs_bypass_0 <=do_bypass;
                    end 
               end 
         if (metaReset)
            begin 
              ex_reg_rs_bypass_1 <=1'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 ex_reg_rs_bypass_1 <=do_bypass_1;
               end 
         if (metaReset)
            begin 
              ex_reg_rs_lsb_0 <=2'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_illegal_insn)
                    begin 
                      ex_reg_rs_lsb_0 <=inst[1:0];
                    end 
                  else 
                    if (_T_40)
                       begin 
                         ex_reg_rs_lsb_0 <=id_rs_0[1:0];
                       end 
                     else 
                       if (id_bypass_src_0_0)
                          begin 
                            ex_reg_rs_lsb_0 <=2'h0;
                          end 
                        else 
                          if (id_bypass_src_0_1)
                             begin 
                               ex_reg_rs_lsb_0 <=2'h1;
                             end 
                           else 
                             if (id_bypass_src_0_2)
                                begin 
                                  ex_reg_rs_lsb_0 <=2'h2;
                                end 
                              else 
                                begin 
                                  ex_reg_rs_lsb_0 <=2'h3;
                                end 
               end 
         if (metaReset)
            begin 
              ex_reg_rs_lsb_1 <=2'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (_T_42)
                    begin 
                      ex_reg_rs_lsb_1 <=id_rs_1[1:0];
                    end 
                  else 
                    if (id_bypass_src_1_0)
                       begin 
                         ex_reg_rs_lsb_1 <=2'h0;
                       end 
                     else 
                       if (id_bypass_src_1_1)
                          begin 
                            ex_reg_rs_lsb_1 <=2'h1;
                          end 
                        else 
                          if (id_bypass_src_1_2)
                             begin 
                               ex_reg_rs_lsb_1 <=2'h2;
                             end 
                           else 
                             begin 
                               ex_reg_rs_lsb_1 <=2'h3;
                             end 
               end 
         if (metaReset)
            begin 
              ex_reg_rs_msb_0 <=62'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (id_illegal_insn)
                    begin 
                      ex_reg_rs_msb_0 <={32'b0,inst[31:2]};
                    end 
                  else 
                    if (_T_40)
                       begin 
                         ex_reg_rs_msb_0 <=id_rs_0[63:2];
                       end 
               end 
         if (metaReset)
            begin 
              ex_reg_rs_msb_1 <=62'h0;
            end 
          else 
            if (~ctrl_killd)
               begin 
                 if (_T_42)
                    begin 
                      ex_reg_rs_msb_1 <=id_rs_1[63:2];
                    end 
               end 
         if (metaReset)
            begin 
              _r <=32'h0;
            end 
          else 
            if (reset)
               begin 
                 _r <=32'h0;
               end 
             else 
               if (_T_138)
                  begin 
                    _r <=_T_137;
                  end 
                else 
                  if (ll_wen)
                     begin 
                       _r <=_T_132;
                     end 
         if (metaReset)
            begin 
              id_stall_fpu__r <=32'h0;
            end 
          else 
            if (reset)
               begin 
                 id_stall_fpu__r <=32'h0;
               end 
             else 
               if (_id_stall_fpu_T_17)
                  begin 
                    id_stall_fpu__r <=_id_stall_fpu_T_16;
                  end 
                else 
                  if (_id_stall_fpu_T_12)
                     begin 
                       id_stall_fpu__r <=_id_stall_fpu_T_11;
                     end 
                   else 
                     if (_id_stall_fpu_T_2)
                        begin 
                          id_stall_fpu__r <=_id_stall_fpu_T_5;
                        end 
         if (metaReset)
            begin 
              blocked <=1'h0;
            end 
          else 
            begin 
              blocked <=_dcache_blocked_blocked_T_3&_dcache_blocked_blocked_T_5;
            end 
         if (metaReset)
            begin 
              div_io_kill_REG <=1'h0;
            end 
          else 
            begin 
              div_io_kill_REG <=div_io_req_ready&div_io_req_valid;
            end 
         if (_GEN_254&~reset)
            begin $display("%d 0x%x (0x%x) f%d p%d 0xXXXXXXXXXXXXXXXX\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn,wb_waddr,_T_142);
            end 
         if (_GEN_257&~reset)
            begin $display("%d 0x%x (0x%x) x%d 0x%x\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn,wb_waddr,rf_wdata);
            end 
         if (_GEN_262&~reset)
            begin $display("%d 0x%x (0x%x) x%d p%d 0xXXXXXXXXXXXXXXXX\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn,wb_waddr,wb_waddr);
            end 
         if (_GEN_268&~reset)
            begin $display("%d 0x%x (0x%x)\n",csr_io_trace_0_priv,csr_io_trace_0_iaddr,csr_io_trace_0_insn);
            end 
         if (_T_159&~reset)
            begin $display("x%d p%d 0x%x\n",rf_waddr,rf_waddr,rf_wdata);
            end 
         Rocket_state <=Rocket_xor0;
         if (!(Rocket_cov_read_data))
            begin 
              Rocket_covSum <=Rocket_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              Rocket_metaAssert <=1'h0;
            end 
          else 
            begin 
              Rocket_metaAssert <=Rocket_metaAssert|Rocket_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (Rocket_cov_write_en&Rocket_cov_write_mask)
            begin 
              Rocket_cov [Rocket_cov_write_addr]<=Rocket_cov_write_data;
            end 
       end
  
endmodule
 
module TLMonitor_23 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_b_ready,
  input io_in_b_valid,
  input [2:0] io_in_b_bits_opcode,
  input [1:0] io_in_b_bits_param,
  input [3:0] io_in_b_bits_size,
  input io_in_b_bits_source,
  input [31:0] io_in_b_bits_address,
  input [7:0] io_in_b_bits_mask,
  input io_in_b_bits_corrupt,
  input io_in_c_ready,
  input io_in_c_valid,
  input [2:0] io_in_c_bits_opcode,
  input [2:0] io_in_c_bits_param,
  input [3:0] io_in_c_bits_size,
  input io_in_c_bits_source,
  input [31:0] io_in_c_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt,
  input io_in_e_ready,
  input io_in_e_valid,
  input [1:0] io_in_e_bits_sink,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [31:0] plusarg_reader_out ;  
   wire [31:0] plusarg_reader_1_out ;  
   wire source_ok ;  
   wire [26:0] _is_aligned_mask_T_1 ;  
   wire [11:0] is_aligned_mask ;  
   wire [31:0] _GEN_86 ;  
   wire [31:0] _is_aligned_T ;  
   wire is_aligned ;  
   wire [1:0] mask_sizeOH_shiftAmount ;  
   wire [3:0] _mask_sizeOH_T_1 ;  
   wire [2:0] mask_sizeOH ;  
   wire _mask_T ;  
   wire mask_size ;  
   wire mask_bit ;  
   wire mask_nbit ;  
   wire _mask_acc_T ;  
   wire mask_acc ;  
   wire _mask_acc_T_1 ;  
   wire mask_acc_1 ;  
   wire mask_size_1 ;  
   wire mask_bit_1 ;  
   wire mask_nbit_1 ;  
   wire mask_eq_2 ;  
   wire _mask_acc_T_2 ;  
   wire mask_acc_2 ;  
   wire mask_eq_3 ;  
   wire _mask_acc_T_3 ;  
   wire mask_acc_3 ;  
   wire mask_eq_4 ;  
   wire _mask_acc_T_4 ;  
   wire mask_acc_4 ;  
   wire mask_eq_5 ;  
   wire _mask_acc_T_5 ;  
   wire mask_acc_5 ;  
   wire mask_size_2 ;  
   wire mask_bit_2 ;  
   wire mask_nbit_2 ;  
   wire mask_eq_6 ;  
   wire _mask_acc_T_6 ;  
   wire mask_lo_lo_lo ;  
   wire mask_eq_7 ;  
   wire _mask_acc_T_7 ;  
   wire mask_lo_lo_hi ;  
   wire mask_eq_8 ;  
   wire _mask_acc_T_8 ;  
   wire mask_lo_hi_lo ;  
   wire mask_eq_9 ;  
   wire _mask_acc_T_9 ;  
   wire mask_lo_hi_hi ;  
   wire mask_eq_10 ;  
   wire _mask_acc_T_10 ;  
   wire mask_hi_lo_lo ;  
   wire mask_eq_11 ;  
   wire _mask_acc_T_11 ;  
   wire mask_hi_lo_hi ;  
   wire mask_eq_12 ;  
   wire _mask_acc_T_12 ;  
   wire mask_hi_hi_lo ;  
   wire mask_eq_13 ;  
   wire _mask_acc_T_13 ;  
   wire mask_hi_hi_hi ;  
   wire [7:0] mask ;  
   wire [32:0] _T_7 ;  
   wire _T_24 ;  
   wire _T_26 ;  
   wire _T_31 ;  
   wire [32:0] _T_37 ;  
   wire _T_38 ;  
   wire [31:0] _T_39 ;  
   wire [32:0] _T_40 ;  
   wire [32:0] _T_42 ;  
   wire _T_43 ;  
   wire [31:0] _T_44 ;  
   wire [32:0] _T_45 ;  
   wire [32:0] _T_47 ;  
   wire _T_48 ;  
   wire [31:0] _T_49 ;  
   wire [32:0] _T_50 ;  
   wire [32:0] _T_52 ;  
   wire _T_53 ;  
   wire [31:0] _T_54 ;  
   wire [32:0] _T_55 ;  
   wire [32:0] _T_57 ;  
   wire _T_58 ;  
   wire [31:0] _T_59 ;  
   wire [32:0] _T_60 ;  
   wire [32:0] _T_62 ;  
   wire _T_63 ;  
   wire _T_64 ;  
   wire _T_65 ;  
   wire _T_66 ;  
   wire _T_67 ;  
   wire _T_68 ;  
   wire _T_71 ;  
   wire [31:0] _T_74 ;  
   wire [32:0] _T_75 ;  
   wire [32:0] _T_77 ;  
   wire _T_78 ;  
   wire _T_79 ;  
   wire _T_82 ;  
   wire _T_84 ;  
   wire _T_88 ;  
   wire _T_89 ;  
   wire _T_136 ;  
   wire _T_137 ;  
   wire _T_139 ;  
   wire _T_141 ;  
   wire _T_144 ;  
   wire _T_148 ;  
   wire _T_151 ;  
   wire _T_153 ;  
   wire _T_155 ;  
   wire _T_158 ;  
   wire _T_160 ;  
   wire _T_166 ;  
   wire _T_299 ;  
   wire _T_301 ;  
   wire _T_312 ;  
   wire _T_322 ;  
   wire _T_333 ;  
   wire _T_368 ;  
   wire _T_369 ;  
   wire _T_370 ;  
   wire _T_371 ;  
   wire _T_372 ;  
   wire _T_373 ;  
   wire _T_375 ;  
   wire _T_377 ;  
   wire _T_385 ;  
   wire _T_387 ;  
   wire _T_389 ;  
   wire _T_391 ;  
   wire _T_397 ;  
   wire _T_440 ;  
   wire _T_441 ;  
   wire _T_442 ;  
   wire _T_443 ;  
   wire _T_452 ;  
   wire _T_460 ;  
   wire _T_462 ;  
   wire _T_464 ;  
   wire _T_465 ;  
   wire _T_467 ;  
   wire _T_483 ;  
   wire [7:0] _T_566 ;  
   wire _T_567 ;  
   wire _T_569 ;  
   wire _T_571 ;  
   wire _T_581 ;  
   wire _T_605 ;  
   wire _T_606 ;  
   wire _T_607 ;  
   wire _T_629 ;  
   wire _T_631 ;  
   wire _T_639 ;  
   wire _T_641 ;  
   wire _T_647 ;  
   wire _T_715 ;  
   wire _T_717 ;  
   wire _T_723 ;  
   wire _T_781 ;  
   wire _T_783 ;  
   wire _T_791 ;  
   wire _T_793 ;  
   wire _T_803 ;  
   wire _T_805 ;  
   wire source_ok_1 ;  
   wire _T_807 ;  
   wire _T_809 ;  
   wire _T_811 ;  
   wire _T_813 ;  
   wire _T_815 ;  
   wire _T_817 ;  
   wire _T_821 ;  
   wire _T_825 ;  
   wire _T_827 ;  
   wire _T_838 ;  
   wire _T_840 ;  
   wire _T_842 ;  
   wire _T_844 ;  
   wire _T_855 ;  
   wire _T_875 ;  
   wire _T_877 ;  
   wire _T_884 ;  
   wire _T_901 ;  
   wire _T_919 ;  
   wire _T_936 ;  
   wire _T_938 ;  
   wire [32:0] _T_943 ;  
   wire [31:0] _address_ok_T ;  
   wire [32:0] _address_ok_T_1 ;  
   wire [32:0] _address_ok_T_3 ;  
   wire _address_ok_T_4 ;  
   wire [31:0] _address_ok_T_5 ;  
   wire [32:0] _address_ok_T_6 ;  
   wire [32:0] _address_ok_T_8 ;  
   wire _address_ok_T_9 ;  
   wire [31:0] _address_ok_T_10 ;  
   wire [32:0] _address_ok_T_11 ;  
   wire [32:0] _address_ok_T_13 ;  
   wire _address_ok_T_14 ;  
   wire [32:0] _address_ok_T_18 ;  
   wire _address_ok_T_19 ;  
   wire [31:0] _address_ok_T_20 ;  
   wire [32:0] _address_ok_T_21 ;  
   wire [32:0] _address_ok_T_23 ;  
   wire _address_ok_T_24 ;  
   wire [31:0] _address_ok_T_25 ;  
   wire [32:0] _address_ok_T_26 ;  
   wire [32:0] _address_ok_T_28 ;  
   wire _address_ok_T_29 ;  
   wire [31:0] _address_ok_T_30 ;  
   wire [32:0] _address_ok_T_31 ;  
   wire [32:0] _address_ok_T_33 ;  
   wire _address_ok_T_34 ;  
   wire _address_ok_T_35 ;  
   wire _address_ok_T_36 ;  
   wire _address_ok_T_37 ;  
   wire _address_ok_T_38 ;  
   wire _address_ok_T_39 ;  
   wire address_ok ;  
   wire [26:0] _is_aligned_mask_T_4 ;  
   wire [11:0] is_aligned_mask_1 ;  
   wire [31:0] _GEN_87 ;  
   wire [31:0] _is_aligned_T_1 ;  
   wire is_aligned_1 ;  
   wire [1:0] mask_sizeOH_shiftAmount_1 ;  
   wire [3:0] _mask_sizeOH_T_4 ;  
   wire [2:0] mask_sizeOH_1 ;  
   wire _mask_T_1 ;  
   wire mask_size_3 ;  
   wire mask_bit_3 ;  
   wire mask_nbit_3 ;  
   wire _mask_acc_T_14 ;  
   wire mask_acc_6 ;  
   wire _mask_acc_T_15 ;  
   wire mask_acc_7 ;  
   wire mask_size_4 ;  
   wire mask_bit_4 ;  
   wire mask_nbit_4 ;  
   wire mask_eq_16 ;  
   wire _mask_acc_T_16 ;  
   wire mask_acc_8 ;  
   wire mask_eq_17 ;  
   wire _mask_acc_T_17 ;  
   wire mask_acc_9 ;  
   wire mask_eq_18 ;  
   wire _mask_acc_T_18 ;  
   wire mask_acc_10 ;  
   wire mask_eq_19 ;  
   wire _mask_acc_T_19 ;  
   wire mask_acc_11 ;  
   wire mask_size_5 ;  
   wire mask_bit_5 ;  
   wire mask_nbit_5 ;  
   wire mask_eq_20 ;  
   wire _mask_acc_T_20 ;  
   wire mask_lo_lo_lo_1 ;  
   wire mask_eq_21 ;  
   wire _mask_acc_T_21 ;  
   wire mask_lo_lo_hi_1 ;  
   wire mask_eq_22 ;  
   wire _mask_acc_T_22 ;  
   wire mask_lo_hi_lo_1 ;  
   wire mask_eq_23 ;  
   wire _mask_acc_T_23 ;  
   wire mask_lo_hi_hi_1 ;  
   wire mask_eq_24 ;  
   wire _mask_acc_T_24 ;  
   wire mask_hi_lo_lo_1 ;  
   wire mask_eq_25 ;  
   wire _mask_acc_T_25 ;  
   wire mask_hi_lo_hi_1 ;  
   wire mask_eq_26 ;  
   wire _mask_acc_T_26 ;  
   wire mask_hi_hi_lo_1 ;  
   wire mask_eq_27 ;  
   wire _mask_acc_T_27 ;  
   wire mask_hi_hi_hi_1 ;  
   wire [7:0] mask_1 ;  
   wire legal_source ;  
   wire _T_960 ;  
   wire _T_963 ;  
   wire _T_964 ;  
   wire _T_968 ;  
   wire _T_1006 ;  
   wire _T_1007 ;  
   wire _T_1008 ;  
   wire _T_1009 ;  
   wire _T_1010 ;  
   wire _T_1011 ;  
   wire _T_1012 ;  
   wire _T_1014 ;  
   wire _T_1016 ;  
   wire _T_1019 ;  
   wire _T_1022 ;  
   wire _T_1025 ;  
   wire _T_1027 ;  
   wire _T_1029 ;  
   wire _T_1031 ;  
   wire _T_1033 ;  
   wire _T_1037 ;  
   wire _T_1039 ;  
   wire _T_1100 ;  
   wire _T_1102 ;  
   wire _T_1112 ;  
   wire _T_1181 ;  
   wire [7:0] _T_1247 ;  
   wire _T_1248 ;  
   wire _T_1250 ;  
   wire _T_1252 ;  
   wire _T_1321 ;  
   wire _T_1390 ;  
   wire source_ok_2 ;  
   wire [26:0] _is_aligned_mask_T_7 ;  
   wire [11:0] is_aligned_mask_2 ;  
   wire [31:0] _GEN_88 ;  
   wire [31:0] _is_aligned_T_2 ;  
   wire is_aligned_2 ;  
   wire [31:0] _address_ok_T_40 ;  
   wire [32:0] _address_ok_T_41 ;  
   wire [32:0] _address_ok_T_43 ;  
   wire _address_ok_T_44 ;  
   wire [31:0] _address_ok_T_45 ;  
   wire [32:0] _address_ok_T_46 ;  
   wire [32:0] _address_ok_T_48 ;  
   wire _address_ok_T_49 ;  
   wire [31:0] _address_ok_T_50 ;  
   wire [32:0] _address_ok_T_51 ;  
   wire [32:0] _address_ok_T_53 ;  
   wire _address_ok_T_54 ;  
   wire [32:0] _address_ok_T_56 ;  
   wire [32:0] _address_ok_T_58 ;  
   wire _address_ok_T_59 ;  
   wire [31:0] _address_ok_T_60 ;  
   wire [32:0] _address_ok_T_61 ;  
   wire [32:0] _address_ok_T_63 ;  
   wire _address_ok_T_64 ;  
   wire [31:0] _address_ok_T_65 ;  
   wire [32:0] _address_ok_T_66 ;  
   wire [32:0] _address_ok_T_68 ;  
   wire _address_ok_T_69 ;  
   wire [31:0] _address_ok_T_70 ;  
   wire [32:0] _address_ok_T_71 ;  
   wire [32:0] _address_ok_T_73 ;  
   wire _address_ok_T_74 ;  
   wire _address_ok_T_75 ;  
   wire _address_ok_T_76 ;  
   wire _address_ok_T_77 ;  
   wire _address_ok_T_78 ;  
   wire _address_ok_T_79 ;  
   wire address_ok_1 ;  
   wire _T_1483 ;  
   wire _T_1485 ;  
   wire _T_1488 ;  
   wire _T_1490 ;  
   wire _T_1492 ;  
   wire _T_1495 ;  
   wire _T_1497 ;  
   wire _T_1499 ;  
   wire _T_1505 ;  
   wire _T_1523 ;  
   wire _T_1525 ;  
   wire _T_1530 ;  
   wire _T_1563 ;  
   wire _T_1564 ;  
   wire _T_1565 ;  
   wire _T_1566 ;  
   wire _T_1567 ;  
   wire _T_1570 ;  
   wire _T_1578 ;  
   wire _T_1581 ;  
   wire _T_1583 ;  
   wire _T_1587 ;  
   wire _T_1588 ;  
   wire _T_1635 ;  
   wire _T_1636 ;  
   wire _T_1638 ;  
   wire _T_1640 ;  
   wire _T_1660 ;  
   wire _T_1793 ;  
   wire _T_1803 ;  
   wire _T_1805 ;  
   wire _T_1811 ;  
   wire _T_1825 ;  
   wire _a_first_T ;  
   wire [8:0] a_first_beats1_decode ;  
   wire a_first_beats1_opdata ;  
   reg [8:0] a_first_counter ;  
   reg [31:0] _RAND_0 ;  
   wire [8:0] a_first_counter1 ;  
   wire a_first ;  
   reg [2:0] opcode ;  
   reg [31:0] _RAND_1 ;  
   reg [2:0] param ;  
   reg [31:0] _RAND_2 ;  
   reg [3:0] size ;  
   reg [31:0] _RAND_3 ;  
   reg source ;  
   reg [31:0] _RAND_4 ;  
   reg [31:0] address ;  
   reg [31:0] _RAND_5 ;  
   wire _T_1847 ;  
   wire _T_1848 ;  
   wire _T_1850 ;  
   wire _T_1852 ;  
   wire _T_1854 ;  
   wire _T_1856 ;  
   wire _T_1858 ;  
   wire _T_1860 ;  
   wire _T_1862 ;  
   wire _T_1864 ;  
   wire _T_1866 ;  
   wire _T_1869 ;  
   wire _d_first_T ;  
   wire [26:0] _d_first_beats1_decode_T_1 ;  
   wire [8:0] d_first_beats1_decode ;  
   wire d_first_beats1_opdata ;  
   reg [8:0] d_first_counter ;  
   reg [31:0] _RAND_6 ;  
   wire [8:0] d_first_counter1 ;  
   wire d_first ;  
   reg [2:0] opcode_1 ;  
   reg [31:0] _RAND_7 ;  
   reg [1:0] param_1 ;  
   reg [31:0] _RAND_8 ;  
   reg [3:0] size_1 ;  
   reg [31:0] _RAND_9 ;  
   reg source_1 ;  
   reg [31:0] _RAND_10 ;  
   reg [1:0] sink ;  
   reg [31:0] _RAND_11 ;  
   reg denied ;  
   reg [31:0] _RAND_12 ;  
   wire _T_1871 ;  
   wire _T_1872 ;  
   wire _T_1874 ;  
   wire _T_1876 ;  
   wire _T_1878 ;  
   wire _T_1880 ;  
   wire _T_1882 ;  
   wire _T_1884 ;  
   wire _T_1886 ;  
   wire _T_1888 ;  
   wire _T_1890 ;  
   wire _T_1892 ;  
   wire _T_1894 ;  
   wire _T_1897 ;  
   wire b_first_done ;  
   reg [8:0] b_first_counter ;  
   reg [31:0] _RAND_13 ;  
   wire [8:0] b_first_counter1 ;  
   wire b_first ;  
   reg [2:0] opcode_2 ;  
   reg [31:0] _RAND_14 ;  
   reg [1:0] param_2 ;  
   reg [31:0] _RAND_15 ;  
   reg [3:0] size_2 ;  
   reg [31:0] _RAND_16 ;  
   reg source_2 ;  
   reg [31:0] _RAND_17 ;  
   reg [31:0] address_1 ;  
   reg [31:0] _RAND_18 ;  
   wire _T_1899 ;  
   wire _T_1900 ;  
   wire _T_1902 ;  
   wire _T_1904 ;  
   wire _T_1906 ;  
   wire _T_1908 ;  
   wire _T_1910 ;  
   wire _T_1912 ;  
   wire _T_1914 ;  
   wire _T_1916 ;  
   wire _T_1918 ;  
   wire _T_1921 ;  
   wire _c_first_T ;  
   wire [8:0] c_first_beats1_decode ;  
   wire c_first_beats1_opdata ;  
   reg [8:0] c_first_counter ;  
   reg [31:0] _RAND_19 ;  
   wire [8:0] c_first_counter1 ;  
   wire c_first ;  
   reg [2:0] opcode_3 ;  
   reg [31:0] _RAND_20 ;  
   reg [2:0] param_3 ;  
   reg [31:0] _RAND_21 ;  
   reg [3:0] size_3 ;  
   reg [31:0] _RAND_22 ;  
   reg source_3 ;  
   reg [31:0] _RAND_23 ;  
   reg [31:0] address_2 ;  
   reg [31:0] _RAND_24 ;  
   wire _T_1923 ;  
   wire _T_1924 ;  
   wire _T_1926 ;  
   wire _T_1928 ;  
   wire _T_1930 ;  
   wire _T_1932 ;  
   wire _T_1934 ;  
   wire _T_1936 ;  
   wire _T_1938 ;  
   wire _T_1940 ;  
   wire _T_1942 ;  
   wire _T_1945 ;  
   reg [1:0] inflight ;  
   reg [31:0] _RAND_25 ;  
   reg [7:0] inflight_opcodes ;  
   reg [31:0] _RAND_26 ;  
   reg [15:0] inflight_sizes ;  
   reg [31:0] _RAND_27 ;  
   reg [8:0] a_first_counter_1 ;  
   reg [31:0] _RAND_28 ;  
   wire [8:0] a_first_counter1_1 ;  
   wire a_first_1 ;  
   reg [8:0] d_first_counter_1 ;  
   reg [31:0] _RAND_29 ;  
   wire [8:0] d_first_counter1_1 ;  
   wire d_first_1 ;  
   wire [2:0] _GEN_89 ;  
   wire [3:0] _a_opcode_lookup_T ;  
   wire [7:0] _a_opcode_lookup_T_1 ;  
   wire [15:0] _a_opcode_lookup_T_5 ;  
   wire [15:0] _GEN_90 ;  
   wire [15:0] _a_opcode_lookup_T_6 ;  
   wire [15:0] _a_opcode_lookup_T_7 ;  
   wire [3:0] _a_size_lookup_T ;  
   wire [15:0] _a_size_lookup_T_1 ;  
   wire [15:0] _a_size_lookup_T_5 ;  
   wire [15:0] _a_size_lookup_T_6 ;  
   wire [15:0] _a_size_lookup_T_7 ;  
   wire _T_1946 ;  
   wire [1:0] _a_set_wo_ready_T ;  
   wire [1:0] a_set_wo_ready ;  
   wire _T_1949 ;  
   wire [3:0] _a_opcodes_set_interm_T ;  
   wire [3:0] _a_opcodes_set_interm_T_1 ;  
   wire [4:0] _a_sizes_set_interm_T ;  
   wire [4:0] _a_sizes_set_interm_T_1 ;  
   wire [2:0] _GEN_93 ;  
   wire [3:0] _a_opcodes_set_T ;  
   wire [3:0] a_opcodes_set_interm ;  
   wire [18:0] _GEN_94 ;  
   wire [18:0] _a_opcodes_set_T_1 ;  
   wire [3:0] _a_sizes_set_T ;  
   wire [4:0] a_sizes_set_interm ;  
   wire [19:0] _GEN_95 ;  
   wire [19:0] _a_sizes_set_T_1 ;  
   wire [1:0] _T_1951 ;  
   wire _T_1955 ;  
   wire [1:0] a_set ;  
   wire [18:0] _GEN_31 ;  
   wire [19:0] _GEN_32 ;  
   wire _T_1957 ;  
   wire _T_1960 ;  
   wire [1:0] _d_clr_wo_ready_T ;  
   wire [1:0] d_clr_wo_ready ;  
   wire _T_1962 ;  
   wire _T_1965 ;  
   wire [30:0] _GEN_97 ;  
   wire [30:0] _d_opcodes_clr_T_5 ;  
   wire [30:0] _GEN_98 ;  
   wire [30:0] _d_sizes_clr_T_5 ;  
   wire [1:0] d_clr ;  
   wire [30:0] _GEN_35 ;  
   wire [30:0] _GEN_36 ;  
   wire _same_cycle_resp_T_2 ;  
   wire same_cycle_resp ;  
   wire [1:0] _T_1970 ;  
   wire _T_1972 ;  
   wire _T_1974 ;  
   wire [2:0] _GEN_39 ;  
   wire [2:0] _GEN_40 ;  
   wire [2:0] _GEN_41 ;  
   wire [2:0] _GEN_42 ;  
   wire [2:0] _GEN_43 ;  
   wire [2:0] _GEN_44 ;  
   wire _T_1976 ;  
   wire [2:0] _GEN_51 ;  
   wire [2:0] _GEN_52 ;  
   wire _T_1977 ;  
   wire _T_1978 ;  
   wire _T_1980 ;  
   wire _T_1982 ;  
   wire _T_1984 ;  
   wire [3:0] a_opcode_lookup ;  
   wire [2:0] _GEN_55 ;  
   wire [2:0] _GEN_56 ;  
   wire [2:0] _GEN_57 ;  
   wire [2:0] _GEN_58 ;  
   wire [2:0] _GEN_59 ;  
   wire [2:0] _GEN_60 ;  
   wire _T_1987 ;  
   wire [2:0] _GEN_67 ;  
   wire [2:0] _GEN_68 ;  
   wire _T_1989 ;  
   wire _T_1990 ;  
   wire _T_1992 ;  
   wire [7:0] a_size_lookup ;  
   wire [7:0] _GEN_99 ;  
   wire _T_1994 ;  
   wire _T_1996 ;  
   wire _T_1999 ;  
   wire _T_2000 ;  
   wire _T_2002 ;  
   wire _T_2004 ;  
   wire _T_2006 ;  
   wire _T_2008 ;  
   wire _T_2010 ;  
   wire _T_2011 ;  
   wire _T_2013 ;  
   wire _T_2015 ;  
   wire [1:0] _inflight_T ;  
   wire [1:0] _inflight_T_2 ;  
   wire [7:0] a_opcodes_set ;  
   wire [7:0] _inflight_opcodes_T ;  
   wire [7:0] d_opcodes_clr ;  
   wire [7:0] _inflight_opcodes_T_2 ;  
   wire [15:0] a_sizes_set ;  
   wire [15:0] _inflight_sizes_T ;  
   wire [15:0] d_sizes_clr ;  
   wire [15:0] _inflight_sizes_T_2 ;  
   reg [31:0] watchdog ;  
   reg [31:0] _RAND_30 ;  
   wire _T_2017 ;  
   wire _T_2019 ;  
   wire _T_2020 ;  
   wire _T_2021 ;  
   wire _T_2022 ;  
   wire _T_2024 ;  
   wire [31:0] _watchdog_T_1 ;  
   wire _T_2028 ;  
   reg [1:0] inflight_1 ;  
   reg [31:0] _RAND_31 ;  
   reg [15:0] inflight_sizes_1 ;  
   reg [31:0] _RAND_32 ;  
   reg [8:0] c_first_counter_1 ;  
   reg [31:0] _RAND_33 ;  
   wire [8:0] c_first_counter1_1 ;  
   wire c_first_1 ;  
   reg [8:0] d_first_counter_2 ;  
   reg [31:0] _RAND_34 ;  
   wire [8:0] d_first_counter1_2 ;  
   wire d_first_2 ;  
   wire [15:0] _c_size_lookup_T_1 ;  
   wire [15:0] _c_size_lookup_T_6 ;  
   wire [15:0] _c_size_lookup_T_7 ;  
   wire _T_2029 ;  
   wire _T_2032 ;  
   wire _T_2033 ;  
   wire [1:0] _c_set_wo_ready_T ;  
   wire [1:0] c_set_wo_ready ;  
   wire _T_2035 ;  
   wire _T_2039 ;  
   wire [4:0] _c_sizes_set_interm_T ;  
   wire [4:0] _c_sizes_set_interm_T_1 ;  
   wire [3:0] _c_sizes_set_T ;  
   wire [4:0] c_sizes_set_interm ;  
   wire [19:0] _GEN_106 ;  
   wire [19:0] _c_sizes_set_T_1 ;  
   wire [1:0] _T_2040 ;  
   wire _T_2044 ;  
   wire [1:0] c_set ;  
   wire [19:0] _GEN_77 ;  
   wire _T_2046 ;  
   wire _T_2048 ;  
   wire [1:0] d_clr_wo_ready_1 ;  
   wire _T_2050 ;  
   wire _T_2052 ;  
   wire [1:0] d_clr_1 ;  
   wire [30:0] _GEN_81 ;  
   wire _same_cycle_resp_T_8 ;  
   wire same_cycle_resp_1 ;  
   wire [1:0] _T_2056 ;  
   wire _T_2058 ;  
   wire _T_2060 ;  
   wire _T_2062 ;  
   wire _T_2064 ;  
   wire [7:0] c_size_lookup ;  
   wire _T_2066 ;  
   wire _T_2068 ;  
   wire _T_2071 ;  
   wire _T_2072 ;  
   wire _T_2074 ;  
   wire _T_2075 ;  
   wire _T_2077 ;  
   wire _T_2079 ;  
   wire _T_2081 ;  
   wire _T_2082 ;  
   wire _T_2084 ;  
   wire [1:0] _inflight_T_3 ;  
   wire [1:0] _inflight_T_5 ;  
   wire [15:0] c_sizes_set ;  
   wire [15:0] _inflight_sizes_T_3 ;  
   wire [15:0] d_sizes_clr_1 ;  
   wire [15:0] _inflight_sizes_T_5 ;  
   reg [31:0] watchdog_1 ;  
   reg [31:0] _RAND_35 ;  
   wire _T_2086 ;  
   wire _T_2088 ;  
   wire _T_2089 ;  
   wire _T_2090 ;  
   wire _T_2091 ;  
   wire _T_2093 ;  
   wire [31:0] _watchdog_T_3 ;  
   wire _T_2097 ;  
   reg [3:0] inflight_2 ;  
   reg [31:0] _RAND_36 ;  
   reg [8:0] d_first_counter_3 ;  
   reg [31:0] _RAND_37 ;  
   wire [8:0] d_first_counter1_3 ;  
   wire d_first_3 ;  
   wire _T_2099 ;  
   wire _T_2103 ;  
   wire _T_2104 ;  
   wire [3:0] _d_set_T ;  
   wire [3:0] _T_2105 ;  
   wire _T_2109 ;  
   wire [3:0] d_set ;  
   wire _T_2111 ;  
   wire [3:0] _e_clr_T ;  
   wire [3:0] _T_2114 ;  
   wire [3:0] _T_2115 ;  
   wire _T_2118 ;  
   wire [3:0] e_clr ;  
   wire [3:0] _inflight_T_6 ;  
   wire [3:0] _inflight_T_8 ;  
   wire _GEN_111 ;  
   wire _GEN_125 ;  
   wire _GEN_141 ;  
   wire _GEN_153 ;  
   wire _GEN_163 ;  
   wire _GEN_173 ;  
   wire _GEN_183 ;  
   wire _GEN_193 ;  
   wire _GEN_203 ;  
   wire _GEN_213 ;  
   wire _GEN_223 ;  
   wire _GEN_233 ;  
   wire _GEN_239 ;  
   wire _GEN_245 ;  
   wire _GEN_251 ;  
   wire _GEN_265 ;  
   wire _GEN_279 ;  
   wire _GEN_291 ;  
   wire _GEN_303 ;  
   wire _GEN_313 ;  
   wire _GEN_323 ;  
   wire _GEN_335 ;  
   wire _GEN_345 ;  
   wire _GEN_355 ;  
   wire _GEN_367 ;  
   wire _GEN_379 ;  
   wire _GEN_387 ;  
   wire _GEN_395 ;  
   wire _GEN_403 ;  
   wire _GEN_408 ;  
   wire _GEN_415 ;  
   wire _GEN_418 ;  
   wire [29:0] TLMonitor_23_covSum ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire stopEn2 ;  
   wire stopEn3 ;  
   wire stopEn4 ;  
   wire stopEn5 ;  
   wire stopEn6 ;  
   wire stopEn7 ;  
   wire stopEn8 ;  
   wire stopEn9 ;  
   wire stopEn10 ;  
   wire stopEn11 ;  
   wire stopEn12 ;  
   wire stopEn13 ;  
   wire stopEn14 ;  
   wire stopEn15 ;  
   wire stopEn16 ;  
   wire stopEn17 ;  
   wire stopEn18 ;  
   wire stopEn19 ;  
   wire stopEn20 ;  
   wire stopEn21 ;  
   wire stopEn22 ;  
   wire stopEn23 ;  
   wire stopEn24 ;  
   wire stopEn25 ;  
   wire stopEn26 ;  
   wire stopEn27 ;  
   wire stopEn28 ;  
   wire stopEn29 ;  
   wire stopEn30 ;  
   wire stopEn31 ;  
   wire stopEn32 ;  
   wire stopEn33 ;  
   wire stopEn34 ;  
   wire stopEn35 ;  
   wire stopEn36 ;  
   wire stopEn37 ;  
   wire stopEn38 ;  
   wire stopEn39 ;  
   wire stopEn40 ;  
   wire stopEn41 ;  
   wire stopEn42 ;  
   wire stopEn43 ;  
   wire stopEn44 ;  
   wire stopEn45 ;  
   wire stopEn46 ;  
   wire stopEn47 ;  
   wire stopEn48 ;  
   wire stopEn49 ;  
   wire stopEn50 ;  
   wire stopEn51 ;  
   wire stopEn52 ;  
   wire stopEn53 ;  
   wire stopEn54 ;  
   wire stopEn55 ;  
   wire stopEn56 ;  
   wire stopEn57 ;  
   wire stopEn58 ;  
   wire stopEn59 ;  
   wire stopEn60 ;  
   wire stopEn61 ;  
   wire stopEn62 ;  
   wire stopEn63 ;  
   wire stopEn64 ;  
   wire stopEn65 ;  
   wire stopEn66 ;  
   wire stopEn67 ;  
   wire stopEn68 ;  
   wire stopEn69 ;  
   wire stopEn70 ;  
   wire stopEn71 ;  
   wire stopEn72 ;  
   wire stopEn73 ;  
   wire stopEn74 ;  
   wire stopEn75 ;  
   wire stopEn76 ;  
   wire stopEn77 ;  
   wire stopEn78 ;  
   wire stopEn79 ;  
   wire stopEn80 ;  
   wire stopEn81 ;  
   wire stopEn82 ;  
   wire stopEn83 ;  
   wire stopEn84 ;  
   wire stopEn85 ;  
   wire stopEn86 ;  
   wire stopEn87 ;  
   wire stopEn88 ;  
   wire stopEn89 ;  
   wire stopEn90 ;  
   wire stopEn91 ;  
   wire stopEn92 ;  
   wire stopEn93 ;  
   wire stopEn94 ;  
   wire stopEn95 ;  
   wire stopEn96 ;  
   wire stopEn97 ;  
   wire stopEn98 ;  
   wire stopEn99 ;  
   wire stopEn100 ;  
   wire stopEn101 ;  
   wire stopEn102 ;  
   wire stopEn103 ;  
   wire stopEn104 ;  
   wire stopEn105 ;  
   wire stopEn106 ;  
   wire stopEn107 ;  
   wire stopEn108 ;  
   wire stopEn109 ;  
   wire stopEn110 ;  
   wire stopEn111 ;  
   wire stopEn112 ;  
   wire stopEn113 ;  
   wire stopEn114 ;  
   wire stopEn115 ;  
   wire stopEn116 ;  
   wire stopEn117 ;  
   wire stopEn118 ;  
   wire stopEn119 ;  
   wire stopEn120 ;  
   wire stopEn121 ;  
   wire stopEn122 ;  
   wire stopEn123 ;  
   wire stopEn124 ;  
   wire stopEn125 ;  
   wire stopEn126 ;  
   wire stopEn127 ;  
   wire stopEn128 ;  
   wire stopEn129 ;  
   wire stopEn130 ;  
   wire stopEn131 ;  
   wire stopEn132 ;  
   wire stopEn133 ;  
   wire stopEn134 ;  
   wire stopEn135 ;  
   wire stopEn136 ;  
   wire stopEn137 ;  
   wire stopEn138 ;  
   wire stopEn139 ;  
   wire stopEn140 ;  
   wire stopEn141 ;  
   wire stopEn142 ;  
   wire stopEn143 ;  
   wire stopEn144 ;  
   wire stopEn145 ;  
   wire stopEn146 ;  
   wire stopEn147 ;  
   wire stopEn148 ;  
   wire stopEn149 ;  
   wire stopEn150 ;  
   wire stopEn151 ;  
   wire stopEn152 ;  
   wire stopEn153 ;  
   wire stopEn154 ;  
   wire stopEn155 ;  
   wire stopEn156 ;  
   wire stopEn157 ;  
   wire stopEn158 ;  
   wire stopEn159 ;  
   wire stopEn160 ;  
   wire stopEn161 ;  
   wire stopEn162 ;  
   wire stopEn163 ;  
   wire stopEn164 ;  
   wire stopEn165 ;  
   wire stopEn166 ;  
   wire stopEn167 ;  
   wire stopEn168 ;  
   wire stopEn169 ;  
   wire stopEn170 ;  
   wire stopEn171 ;  
   wire stopEn172 ;  
   wire stopEn173 ;  
   wire stopEn174 ;  
   wire stopEn175 ;  
   wire stopEn176 ;  
   wire stopEn177 ;  
   wire stopEn178 ;  
   wire stopEn179 ;  
   wire stopEn180 ;  
   wire stopEn181 ;  
   wire stopEn182 ;  
   wire stopEn183 ;  
   wire stopEn184 ;  
   wire stopEn185 ;  
   wire stopEn186 ;  
   wire plusarg_reader_metaAssert_wire ;  
   wire plusarg_reader_1_metaAssert_wire ;  
   wire TLMonitor_23_or63 ;  
   wire TLMonitor_23_or130 ;  
   wire TLMonitor_23_or64 ;  
   wire TLMonitor_23_or31 ;  
   wire TLMonitor_23_or132 ;  
   wire TLMonitor_23_or65 ;  
   wire TLMonitor_23_or134 ;  
   wire TLMonitor_23_or66 ;  
   wire TLMonitor_23_or32 ;  
   wire TLMonitor_23_or15 ;  
   wire TLMonitor_23_or136 ;  
   wire TLMonitor_23_or67 ;  
   wire TLMonitor_23_or138 ;  
   wire TLMonitor_23_or68 ;  
   wire TLMonitor_23_or33 ;  
   wire TLMonitor_23_or140 ;  
   wire TLMonitor_23_or69 ;  
   wire TLMonitor_23_or142 ;  
   wire TLMonitor_23_or70 ;  
   wire TLMonitor_23_or34 ;  
   wire TLMonitor_23_or16 ;  
   wire TLMonitor_23_or7 ;  
   wire TLMonitor_23_or144 ;  
   wire TLMonitor_23_or71 ;  
   wire TLMonitor_23_or146 ;  
   wire TLMonitor_23_or72 ;  
   wire TLMonitor_23_or35 ;  
   wire TLMonitor_23_or148 ;  
   wire TLMonitor_23_or73 ;  
   wire TLMonitor_23_or150 ;  
   wire TLMonitor_23_or74 ;  
   wire TLMonitor_23_or36 ;  
   wire TLMonitor_23_or17 ;  
   wire TLMonitor_23_or152 ;  
   wire TLMonitor_23_or75 ;  
   wire TLMonitor_23_or154 ;  
   wire TLMonitor_23_or76 ;  
   wire TLMonitor_23_or37 ;  
   wire TLMonitor_23_or156 ;  
   wire TLMonitor_23_or77 ;  
   wire TLMonitor_23_or158 ;  
   wire TLMonitor_23_or78 ;  
   wire TLMonitor_23_or38 ;  
   wire TLMonitor_23_or18 ;  
   wire TLMonitor_23_or8 ;  
   wire TLMonitor_23_or3 ;  
   wire TLMonitor_23_or79 ;  
   wire TLMonitor_23_or162 ;  
   wire TLMonitor_23_or80 ;  
   wire TLMonitor_23_or39 ;  
   wire TLMonitor_23_or164 ;  
   wire TLMonitor_23_or81 ;  
   wire TLMonitor_23_or166 ;  
   wire TLMonitor_23_or82 ;  
   wire TLMonitor_23_or40 ;  
   wire TLMonitor_23_or19 ;  
   wire TLMonitor_23_or168 ;  
   wire TLMonitor_23_or83 ;  
   wire TLMonitor_23_or170 ;  
   wire TLMonitor_23_or84 ;  
   wire TLMonitor_23_or41 ;  
   wire TLMonitor_23_or172 ;  
   wire TLMonitor_23_or85 ;  
   wire TLMonitor_23_or174 ;  
   wire TLMonitor_23_or86 ;  
   wire TLMonitor_23_or42 ;  
   wire TLMonitor_23_or20 ;  
   wire TLMonitor_23_or9 ;  
   wire TLMonitor_23_or176 ;  
   wire TLMonitor_23_or87 ;  
   wire TLMonitor_23_or178 ;  
   wire TLMonitor_23_or88 ;  
   wire TLMonitor_23_or43 ;  
   wire TLMonitor_23_or180 ;  
   wire TLMonitor_23_or89 ;  
   wire TLMonitor_23_or182 ;  
   wire TLMonitor_23_or90 ;  
   wire TLMonitor_23_or44 ;  
   wire TLMonitor_23_or21 ;  
   wire TLMonitor_23_or184 ;  
   wire TLMonitor_23_or91 ;  
   wire TLMonitor_23_or186 ;  
   wire TLMonitor_23_or92 ;  
   wire TLMonitor_23_or45 ;  
   wire TLMonitor_23_or188 ;  
   wire TLMonitor_23_or93 ;  
   wire TLMonitor_23_or190 ;  
   wire TLMonitor_23_or94 ;  
   wire TLMonitor_23_or46 ;  
   wire TLMonitor_23_or22 ;  
   wire TLMonitor_23_or10 ;  
   wire TLMonitor_23_or4 ;  
   wire TLMonitor_23_or1 ;  
   wire TLMonitor_23_or95 ;  
   wire TLMonitor_23_or194 ;  
   wire TLMonitor_23_or96 ;  
   wire TLMonitor_23_or47 ;  
   wire TLMonitor_23_or196 ;  
   wire TLMonitor_23_or97 ;  
   wire TLMonitor_23_or198 ;  
   wire TLMonitor_23_or98 ;  
   wire TLMonitor_23_or48 ;  
   wire TLMonitor_23_or23 ;  
   wire TLMonitor_23_or200 ;  
   wire TLMonitor_23_or99 ;  
   wire TLMonitor_23_or202 ;  
   wire TLMonitor_23_or100 ;  
   wire TLMonitor_23_or49 ;  
   wire TLMonitor_23_or204 ;  
   wire TLMonitor_23_or101 ;  
   wire TLMonitor_23_or206 ;  
   wire TLMonitor_23_or102 ;  
   wire TLMonitor_23_or50 ;  
   wire TLMonitor_23_or24 ;  
   wire TLMonitor_23_or11 ;  
   wire TLMonitor_23_or208 ;  
   wire TLMonitor_23_or103 ;  
   wire TLMonitor_23_or210 ;  
   wire TLMonitor_23_or104 ;  
   wire TLMonitor_23_or51 ;  
   wire TLMonitor_23_or212 ;  
   wire TLMonitor_23_or105 ;  
   wire TLMonitor_23_or214 ;  
   wire TLMonitor_23_or106 ;  
   wire TLMonitor_23_or52 ;  
   wire TLMonitor_23_or25 ;  
   wire TLMonitor_23_or216 ;  
   wire TLMonitor_23_or107 ;  
   wire TLMonitor_23_or218 ;  
   wire TLMonitor_23_or108 ;  
   wire TLMonitor_23_or53 ;  
   wire TLMonitor_23_or220 ;  
   wire TLMonitor_23_or109 ;  
   wire TLMonitor_23_or222 ;  
   wire TLMonitor_23_or110 ;  
   wire TLMonitor_23_or54 ;  
   wire TLMonitor_23_or26 ;  
   wire TLMonitor_23_or12 ;  
   wire TLMonitor_23_or5 ;  
   wire TLMonitor_23_or224 ;  
   wire TLMonitor_23_or111 ;  
   wire TLMonitor_23_or226 ;  
   wire TLMonitor_23_or112 ;  
   wire TLMonitor_23_or55 ;  
   wire TLMonitor_23_or228 ;  
   wire TLMonitor_23_or113 ;  
   wire TLMonitor_23_or230 ;  
   wire TLMonitor_23_or114 ;  
   wire TLMonitor_23_or56 ;  
   wire TLMonitor_23_or27 ;  
   wire TLMonitor_23_or232 ;  
   wire TLMonitor_23_or115 ;  
   wire TLMonitor_23_or234 ;  
   wire TLMonitor_23_or116 ;  
   wire TLMonitor_23_or57 ;  
   wire TLMonitor_23_or236 ;  
   wire TLMonitor_23_or117 ;  
   wire TLMonitor_23_or238 ;  
   wire TLMonitor_23_or118 ;  
   wire TLMonitor_23_or58 ;  
   wire TLMonitor_23_or28 ;  
   wire TLMonitor_23_or13 ;  
   wire TLMonitor_23_or240 ;  
   wire TLMonitor_23_or119 ;  
   wire TLMonitor_23_or242 ;  
   wire TLMonitor_23_or120 ;  
   wire TLMonitor_23_or59 ;  
   wire TLMonitor_23_or244 ;  
   wire TLMonitor_23_or121 ;  
   wire TLMonitor_23_or246 ;  
   wire TLMonitor_23_or122 ;  
   wire TLMonitor_23_or60 ;  
   wire TLMonitor_23_or29 ;  
   wire TLMonitor_23_or248 ;  
   wire TLMonitor_23_or123 ;  
   wire TLMonitor_23_or250 ;  
   wire TLMonitor_23_or124 ;  
   wire TLMonitor_23_or61 ;  
   wire TLMonitor_23_or252 ;  
   wire TLMonitor_23_or125 ;  
   wire TLMonitor_23_or254 ;  
   wire TLMonitor_23_or126 ;  
   wire TLMonitor_23_or62 ;  
   wire TLMonitor_23_or30 ;  
   wire TLMonitor_23_or14 ;  
   wire TLMonitor_23_or6 ;  
   wire TLMonitor_23_or2 ;  
   wire TLMonitor_23_or0 ;  
   reg TLMonitor_23_metaAssert ;  
   reg [31:0] _RAND_38 ;  
  assign source_ok=~io_in_a_bits_source|io_in_a_bits_source; 
  assign _is_aligned_mask_T_1=27'hfff<<io_in_a_bits_size; 
  assign is_aligned_mask=~_is_aligned_mask_T_1[11:0]; 
  assign _GEN_86={20'b0,is_aligned_mask}; 
  assign _is_aligned_T=io_in_a_bits_address&_GEN_86; 
  assign is_aligned=_is_aligned_T==32'h0; 
  assign mask_sizeOH_shiftAmount=io_in_a_bits_size[1:0]; 
  assign _mask_sizeOH_T_1=4'h1<<mask_sizeOH_shiftAmount; 
  assign mask_sizeOH=_mask_sizeOH_T_1[2:0]|3'h1; 
  assign _mask_T=io_in_a_bits_size>=4'h3; 
  assign mask_size=mask_sizeOH[2]; 
  assign mask_bit=io_in_a_bits_address[2]; 
  assign mask_nbit=~mask_bit; 
  assign _mask_acc_T=mask_size&mask_nbit; 
  assign mask_acc=_mask_T|_mask_acc_T; 
  assign _mask_acc_T_1=mask_size&mask_bit; 
  assign mask_acc_1=_mask_T|_mask_acc_T_1; 
  assign mask_size_1=mask_sizeOH[1]; 
  assign mask_bit_1=io_in_a_bits_address[1]; 
  assign mask_nbit_1=~mask_bit_1; 
  assign mask_eq_2=mask_nbit&mask_nbit_1; 
  assign _mask_acc_T_2=mask_size_1&mask_eq_2; 
  assign mask_acc_2=mask_acc|_mask_acc_T_2; 
  assign mask_eq_3=mask_nbit&mask_bit_1; 
  assign _mask_acc_T_3=mask_size_1&mask_eq_3; 
  assign mask_acc_3=mask_acc|_mask_acc_T_3; 
  assign mask_eq_4=mask_bit&mask_nbit_1; 
  assign _mask_acc_T_4=mask_size_1&mask_eq_4; 
  assign mask_acc_4=mask_acc_1|_mask_acc_T_4; 
  assign mask_eq_5=mask_bit&mask_bit_1; 
  assign _mask_acc_T_5=mask_size_1&mask_eq_5; 
  assign mask_acc_5=mask_acc_1|_mask_acc_T_5; 
  assign mask_size_2=mask_sizeOH[0]; 
  assign mask_bit_2=io_in_a_bits_address[0]; 
  assign mask_nbit_2=~mask_bit_2; 
  assign mask_eq_6=mask_eq_2&mask_nbit_2; 
  assign _mask_acc_T_6=mask_size_2&mask_eq_6; 
  assign mask_lo_lo_lo=mask_acc_2|_mask_acc_T_6; 
  assign mask_eq_7=mask_eq_2&mask_bit_2; 
  assign _mask_acc_T_7=mask_size_2&mask_eq_7; 
  assign mask_lo_lo_hi=mask_acc_2|_mask_acc_T_7; 
  assign mask_eq_8=mask_eq_3&mask_nbit_2; 
  assign _mask_acc_T_8=mask_size_2&mask_eq_8; 
  assign mask_lo_hi_lo=mask_acc_3|_mask_acc_T_8; 
  assign mask_eq_9=mask_eq_3&mask_bit_2; 
  assign _mask_acc_T_9=mask_size_2&mask_eq_9; 
  assign mask_lo_hi_hi=mask_acc_3|_mask_acc_T_9; 
  assign mask_eq_10=mask_eq_4&mask_nbit_2; 
  assign _mask_acc_T_10=mask_size_2&mask_eq_10; 
  assign mask_hi_lo_lo=mask_acc_4|_mask_acc_T_10; 
  assign mask_eq_11=mask_eq_4&mask_bit_2; 
  assign _mask_acc_T_11=mask_size_2&mask_eq_11; 
  assign mask_hi_lo_hi=mask_acc_4|_mask_acc_T_11; 
  assign mask_eq_12=mask_eq_5&mask_nbit_2; 
  assign _mask_acc_T_12=mask_size_2&mask_eq_12; 
  assign mask_hi_hi_lo=mask_acc_5|_mask_acc_T_12; 
  assign mask_eq_13=mask_eq_5&mask_bit_2; 
  assign _mask_acc_T_13=mask_size_2&mask_eq_13; 
  assign mask_hi_hi_hi=mask_acc_5|_mask_acc_T_13; 
  assign mask={mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,mask_lo_lo_lo}; 
  assign _T_7={1'b0,$signed(io_in_a_bits_address)}; 
  assign _T_24=io_in_a_bits_opcode==3'h6; 
  assign _T_26=io_in_a_bits_size<=4'hc; 
  assign _T_31=_T_26&source_ok; 
  assign _T_37=$signed(_T_7)&-33'sh1000; 
  assign _T_38=$signed(_T_37)==33'sh0; 
  assign _T_39=io_in_a_bits_address^32'h3000; 
  assign _T_40={1'b0,$signed(_T_39)}; 
  assign _T_42=$signed(_T_40)&-33'sh1000; 
  assign _T_43=$signed(_T_42)==33'sh0; 
  assign _T_44=io_in_a_bits_address^32'h10000; 
  assign _T_45={1'b0,$signed(_T_44)}; 
  assign _T_47=$signed(_T_45)&-33'sh10000; 
  assign _T_48=$signed(_T_47)==33'sh0; 
  assign _T_49=io_in_a_bits_address^32'h2000000; 
  assign _T_50={1'b0,$signed(_T_49)}; 
  assign _T_52=$signed(_T_50)&-33'sh10000; 
  assign _T_53=$signed(_T_52)==33'sh0; 
  assign _T_54=io_in_a_bits_address^32'hc000000; 
  assign _T_55={1'b0,$signed(_T_54)}; 
  assign _T_57=$signed(_T_55)&-33'sh4000000; 
  assign _T_58=$signed(_T_57)==33'sh0; 
  assign _T_59=io_in_a_bits_address^32'h60000000; 
  assign _T_60={1'b0,$signed(_T_59)}; 
  assign _T_62=$signed(_T_60)&-33'sh20000000; 
  assign _T_63=$signed(_T_62)==33'sh0; 
  assign _T_64=_T_38|_T_43; 
  assign _T_65=_T_64|_T_48; 
  assign _T_66=_T_65|_T_53; 
  assign _T_67=_T_66|_T_58; 
  assign _T_68=_T_67|_T_63; 
  assign _T_71=io_in_a_bits_size<=4'h6; 
  assign _T_74=io_in_a_bits_address^32'h80000000; 
  assign _T_75={1'b0,$signed(_T_74)}; 
  assign _T_77=$signed(_T_75)&-33'sh10000000; 
  assign _T_78=$signed(_T_77)==33'sh0; 
  assign _T_79=_T_71&_T_78; 
  assign _T_82=_T_31&_T_79; 
  assign _T_84=_T_82|reset; 
  assign _T_88=4'h6==io_in_a_bits_size; 
  assign _T_89=~io_in_a_bits_source&_T_88; 
  assign _T_136=_T_68|_T_78; 
  assign _T_137=_T_26&_T_136; 
  assign _T_139=_T_89&_T_137; 
  assign _T_141=_T_139|reset; 
  assign _T_144=source_ok|reset; 
  assign _T_148=_mask_T|reset; 
  assign _T_151=is_aligned|reset; 
  assign _T_153=io_in_a_bits_param<=3'h2; 
  assign _T_155=_T_153|reset; 
  assign _T_158=~io_in_a_bits_mask==8'h0; 
  assign _T_160=_T_158|reset; 
  assign _T_166=io_in_a_bits_opcode==3'h7; 
  assign _T_299=io_in_a_bits_param!=3'h0; 
  assign _T_301=_T_299|reset; 
  assign _T_312=io_in_a_bits_opcode==3'h4; 
  assign _T_322=_T_31|reset; 
  assign _T_333=_T_26&_T_43; 
  assign _T_368=_T_38|_T_48; 
  assign _T_369=_T_368|_T_53; 
  assign _T_370=_T_369|_T_58; 
  assign _T_371=_T_370|_T_63; 
  assign _T_372=_T_371|_T_78; 
  assign _T_373=_T_71&_T_372; 
  assign _T_375=_T_333|_T_373; 
  assign _T_377=_T_375|reset; 
  assign _T_385=io_in_a_bits_param==3'h0; 
  assign _T_387=_T_385|reset; 
  assign _T_389=io_in_a_bits_mask==mask; 
  assign _T_391=_T_389|reset; 
  assign _T_397=io_in_a_bits_opcode==3'h0; 
  assign _T_440=_T_38|_T_53; 
  assign _T_441=_T_440|_T_58; 
  assign _T_442=_T_441|_T_78; 
  assign _T_443=_T_71&_T_442; 
  assign _T_452=io_in_a_bits_size<=4'h8; 
  assign _T_460=_T_452&_T_63; 
  assign _T_462=_T_333|_T_443; 
  assign _T_464=_T_462|_T_460; 
  assign _T_465=_T_31&_T_464; 
  assign _T_467=_T_465|reset; 
  assign _T_483=io_in_a_bits_opcode==3'h1; 
  assign _T_566=io_in_a_bits_mask&~mask; 
  assign _T_567=_T_566==8'h0; 
  assign _T_569=_T_567|reset; 
  assign _T_571=io_in_a_bits_opcode==3'h2; 
  assign _T_581=io_in_a_bits_size<=4'h3; 
  assign _T_605=_T_64|_T_53; 
  assign _T_606=_T_605|_T_58; 
  assign _T_607=_T_581&_T_606; 
  assign _T_629=_T_31&_T_607; 
  assign _T_631=_T_629|reset; 
  assign _T_639=io_in_a_bits_param<=3'h4; 
  assign _T_641=_T_639|reset; 
  assign _T_647=io_in_a_bits_opcode==3'h3; 
  assign _T_715=io_in_a_bits_param<=3'h3; 
  assign _T_717=_T_715|reset; 
  assign _T_723=io_in_a_bits_opcode==3'h5; 
  assign _T_781=_T_31&_T_333; 
  assign _T_783=_T_781|reset; 
  assign _T_791=io_in_a_bits_param<=3'h1; 
  assign _T_793=_T_791|reset; 
  assign _T_803=io_in_d_bits_opcode<=3'h6; 
  assign _T_805=_T_803|reset; 
  assign source_ok_1=~io_in_d_bits_source|io_in_d_bits_source; 
  assign _T_807=io_in_d_bits_opcode==3'h6; 
  assign _T_809=source_ok_1|reset; 
  assign _T_811=io_in_d_bits_size>=4'h3; 
  assign _T_813=_T_811|reset; 
  assign _T_815=io_in_d_bits_param==2'h0; 
  assign _T_817=_T_815|reset; 
  assign _T_821=~io_in_d_bits_corrupt|reset; 
  assign _T_825=~io_in_d_bits_denied|reset; 
  assign _T_827=io_in_d_bits_opcode==3'h4; 
  assign _T_838=io_in_d_bits_param<=2'h2; 
  assign _T_840=_T_838|reset; 
  assign _T_842=io_in_d_bits_param!=2'h2; 
  assign _T_844=_T_842|reset; 
  assign _T_855=io_in_d_bits_opcode==3'h5; 
  assign _T_875=~io_in_d_bits_denied|io_in_d_bits_corrupt; 
  assign _T_877=_T_875|reset; 
  assign _T_884=io_in_d_bits_opcode==3'h0; 
  assign _T_901=io_in_d_bits_opcode==3'h1; 
  assign _T_919=io_in_d_bits_opcode==3'h2; 
  assign _T_936=io_in_b_bits_opcode<=3'h6; 
  assign _T_938=_T_936|reset; 
  assign _T_943={1'b0,$signed(io_in_b_bits_address)}; 
  assign _address_ok_T=io_in_b_bits_address^32'h3000; 
  assign _address_ok_T_1={1'b0,$signed(_address_ok_T)}; 
  assign _address_ok_T_3=$signed(_address_ok_T_1)&-33'sh1000; 
  assign _address_ok_T_4=$signed(_address_ok_T_3)==33'sh0; 
  assign _address_ok_T_5=io_in_b_bits_address^32'hc000000; 
  assign _address_ok_T_6={1'b0,$signed(_address_ok_T_5)}; 
  assign _address_ok_T_8=$signed(_address_ok_T_6)&-33'sh4000000; 
  assign _address_ok_T_9=$signed(_address_ok_T_8)==33'sh0; 
  assign _address_ok_T_10=io_in_b_bits_address^32'h2000000; 
  assign _address_ok_T_11={1'b0,$signed(_address_ok_T_10)}; 
  assign _address_ok_T_13=$signed(_address_ok_T_11)&-33'sh10000; 
  assign _address_ok_T_14=$signed(_address_ok_T_13)==33'sh0; 
  assign _address_ok_T_18=$signed(_T_943)&-33'sh1000; 
  assign _address_ok_T_19=$signed(_address_ok_T_18)==33'sh0; 
  assign _address_ok_T_20=io_in_b_bits_address^32'h10000; 
  assign _address_ok_T_21={1'b0,$signed(_address_ok_T_20)}; 
  assign _address_ok_T_23=$signed(_address_ok_T_21)&-33'sh10000; 
  assign _address_ok_T_24=$signed(_address_ok_T_23)==33'sh0; 
  assign _address_ok_T_25=io_in_b_bits_address^32'h80000000; 
  assign _address_ok_T_26={1'b0,$signed(_address_ok_T_25)}; 
  assign _address_ok_T_28=$signed(_address_ok_T_26)&-33'sh10000000; 
  assign _address_ok_T_29=$signed(_address_ok_T_28)==33'sh0; 
  assign _address_ok_T_30=io_in_b_bits_address^32'h60000000; 
  assign _address_ok_T_31={1'b0,$signed(_address_ok_T_30)}; 
  assign _address_ok_T_33=$signed(_address_ok_T_31)&-33'sh20000000; 
  assign _address_ok_T_34=$signed(_address_ok_T_33)==33'sh0; 
  assign _address_ok_T_35=_address_ok_T_4|_address_ok_T_9; 
  assign _address_ok_T_36=_address_ok_T_35|_address_ok_T_14; 
  assign _address_ok_T_37=_address_ok_T_36|_address_ok_T_19; 
  assign _address_ok_T_38=_address_ok_T_37|_address_ok_T_24; 
  assign _address_ok_T_39=_address_ok_T_38|_address_ok_T_29; 
  assign address_ok=_address_ok_T_39|_address_ok_T_34; 
  assign _is_aligned_mask_T_4=27'hfff<<io_in_b_bits_size; 
  assign is_aligned_mask_1=~_is_aligned_mask_T_4[11:0]; 
  assign _GEN_87={20'b0,is_aligned_mask_1}; 
  assign _is_aligned_T_1=io_in_b_bits_address&_GEN_87; 
  assign is_aligned_1=_is_aligned_T_1==32'h0; 
  assign mask_sizeOH_shiftAmount_1=io_in_b_bits_size[1:0]; 
  assign _mask_sizeOH_T_4=4'h1<<mask_sizeOH_shiftAmount_1; 
  assign mask_sizeOH_1=_mask_sizeOH_T_4[2:0]|3'h1; 
  assign _mask_T_1=io_in_b_bits_size>=4'h3; 
  assign mask_size_3=mask_sizeOH_1[2]; 
  assign mask_bit_3=io_in_b_bits_address[2]; 
  assign mask_nbit_3=~mask_bit_3; 
  assign _mask_acc_T_14=mask_size_3&mask_nbit_3; 
  assign mask_acc_6=_mask_T_1|_mask_acc_T_14; 
  assign _mask_acc_T_15=mask_size_3&mask_bit_3; 
  assign mask_acc_7=_mask_T_1|_mask_acc_T_15; 
  assign mask_size_4=mask_sizeOH_1[1]; 
  assign mask_bit_4=io_in_b_bits_address[1]; 
  assign mask_nbit_4=~mask_bit_4; 
  assign mask_eq_16=mask_nbit_3&mask_nbit_4; 
  assign _mask_acc_T_16=mask_size_4&mask_eq_16; 
  assign mask_acc_8=mask_acc_6|_mask_acc_T_16; 
  assign mask_eq_17=mask_nbit_3&mask_bit_4; 
  assign _mask_acc_T_17=mask_size_4&mask_eq_17; 
  assign mask_acc_9=mask_acc_6|_mask_acc_T_17; 
  assign mask_eq_18=mask_bit_3&mask_nbit_4; 
  assign _mask_acc_T_18=mask_size_4&mask_eq_18; 
  assign mask_acc_10=mask_acc_7|_mask_acc_T_18; 
  assign mask_eq_19=mask_bit_3&mask_bit_4; 
  assign _mask_acc_T_19=mask_size_4&mask_eq_19; 
  assign mask_acc_11=mask_acc_7|_mask_acc_T_19; 
  assign mask_size_5=mask_sizeOH_1[0]; 
  assign mask_bit_5=io_in_b_bits_address[0]; 
  assign mask_nbit_5=~mask_bit_5; 
  assign mask_eq_20=mask_eq_16&mask_nbit_5; 
  assign _mask_acc_T_20=mask_size_5&mask_eq_20; 
  assign mask_lo_lo_lo_1=mask_acc_8|_mask_acc_T_20; 
  assign mask_eq_21=mask_eq_16&mask_bit_5; 
  assign _mask_acc_T_21=mask_size_5&mask_eq_21; 
  assign mask_lo_lo_hi_1=mask_acc_8|_mask_acc_T_21; 
  assign mask_eq_22=mask_eq_17&mask_nbit_5; 
  assign _mask_acc_T_22=mask_size_5&mask_eq_22; 
  assign mask_lo_hi_lo_1=mask_acc_9|_mask_acc_T_22; 
  assign mask_eq_23=mask_eq_17&mask_bit_5; 
  assign _mask_acc_T_23=mask_size_5&mask_eq_23; 
  assign mask_lo_hi_hi_1=mask_acc_9|_mask_acc_T_23; 
  assign mask_eq_24=mask_eq_18&mask_nbit_5; 
  assign _mask_acc_T_24=mask_size_5&mask_eq_24; 
  assign mask_hi_lo_lo_1=mask_acc_10|_mask_acc_T_24; 
  assign mask_eq_25=mask_eq_18&mask_bit_5; 
  assign _mask_acc_T_25=mask_size_5&mask_eq_25; 
  assign mask_hi_lo_hi_1=mask_acc_10|_mask_acc_T_25; 
  assign mask_eq_26=mask_eq_19&mask_nbit_5; 
  assign _mask_acc_T_26=mask_size_5&mask_eq_26; 
  assign mask_hi_hi_lo_1=mask_acc_11|_mask_acc_T_26; 
  assign mask_eq_27=mask_eq_19&mask_bit_5; 
  assign _mask_acc_T_27=mask_size_5&mask_eq_27; 
  assign mask_hi_hi_hi_1=mask_acc_11|_mask_acc_T_27; 
  assign mask_1={mask_hi_hi_hi_1,mask_hi_hi_lo_1,mask_hi_lo_hi_1,mask_hi_lo_lo_1,mask_lo_hi_hi_1,mask_lo_hi_lo_1,mask_lo_lo_hi_1,mask_lo_lo_lo_1}; 
  assign legal_source=io_in_b_bits_source==io_in_b_bits_source; 
  assign _T_960=io_in_b_bits_opcode==3'h6; 
  assign _T_963=4'h6==io_in_b_bits_size; 
  assign _T_964=~io_in_b_bits_source&_T_963; 
  assign _T_968=io_in_b_bits_size<=4'hc; 
  assign _T_1006=_address_ok_T_19|_address_ok_T_4; 
  assign _T_1007=_T_1006|_address_ok_T_24; 
  assign _T_1008=_T_1007|_address_ok_T_14; 
  assign _T_1009=_T_1008|_address_ok_T_9; 
  assign _T_1010=_T_1009|_address_ok_T_34; 
  assign _T_1011=_T_1010|_address_ok_T_29; 
  assign _T_1012=_T_968&_T_1011; 
  assign _T_1014=_T_964&_T_1012; 
  assign _T_1016=_T_1014|reset; 
  assign _T_1019=address_ok|reset; 
  assign _T_1022=legal_source|reset; 
  assign _T_1025=is_aligned_1|reset; 
  assign _T_1027=io_in_b_bits_param<=2'h2; 
  assign _T_1029=_T_1027|reset; 
  assign _T_1031=io_in_b_bits_mask==mask_1; 
  assign _T_1033=_T_1031|reset; 
  assign _T_1037=~io_in_b_bits_corrupt|reset; 
  assign _T_1039=io_in_b_bits_opcode==3'h4; 
  assign _T_1100=io_in_b_bits_param==2'h0; 
  assign _T_1102=_T_1100|reset; 
  assign _T_1112=io_in_b_bits_opcode==3'h0; 
  assign _T_1181=io_in_b_bits_opcode==3'h1; 
  assign _T_1247=io_in_b_bits_mask&~mask_1; 
  assign _T_1248=_T_1247==8'h0; 
  assign _T_1250=_T_1248|reset; 
  assign _T_1252=io_in_b_bits_opcode==3'h2; 
  assign _T_1321=io_in_b_bits_opcode==3'h3; 
  assign _T_1390=io_in_b_bits_opcode==3'h5; 
  assign source_ok_2=~io_in_c_bits_source|io_in_c_bits_source; 
  assign _is_aligned_mask_T_7=27'hfff<<io_in_c_bits_size; 
  assign is_aligned_mask_2=~_is_aligned_mask_T_7[11:0]; 
  assign _GEN_88={20'b0,is_aligned_mask_2}; 
  assign _is_aligned_T_2=io_in_c_bits_address&_GEN_88; 
  assign is_aligned_2=_is_aligned_T_2==32'h0; 
  assign _address_ok_T_40=io_in_c_bits_address^32'h3000; 
  assign _address_ok_T_41={1'b0,$signed(_address_ok_T_40)}; 
  assign _address_ok_T_43=$signed(_address_ok_T_41)&-33'sh1000; 
  assign _address_ok_T_44=$signed(_address_ok_T_43)==33'sh0; 
  assign _address_ok_T_45=io_in_c_bits_address^32'hc000000; 
  assign _address_ok_T_46={1'b0,$signed(_address_ok_T_45)}; 
  assign _address_ok_T_48=$signed(_address_ok_T_46)&-33'sh4000000; 
  assign _address_ok_T_49=$signed(_address_ok_T_48)==33'sh0; 
  assign _address_ok_T_50=io_in_c_bits_address^32'h2000000; 
  assign _address_ok_T_51={1'b0,$signed(_address_ok_T_50)}; 
  assign _address_ok_T_53=$signed(_address_ok_T_51)&-33'sh10000; 
  assign _address_ok_T_54=$signed(_address_ok_T_53)==33'sh0; 
  assign _address_ok_T_56={1'b0,$signed(io_in_c_bits_address)}; 
  assign _address_ok_T_58=$signed(_address_ok_T_56)&-33'sh1000; 
  assign _address_ok_T_59=$signed(_address_ok_T_58)==33'sh0; 
  assign _address_ok_T_60=io_in_c_bits_address^32'h10000; 
  assign _address_ok_T_61={1'b0,$signed(_address_ok_T_60)}; 
  assign _address_ok_T_63=$signed(_address_ok_T_61)&-33'sh10000; 
  assign _address_ok_T_64=$signed(_address_ok_T_63)==33'sh0; 
  assign _address_ok_T_65=io_in_c_bits_address^32'h80000000; 
  assign _address_ok_T_66={1'b0,$signed(_address_ok_T_65)}; 
  assign _address_ok_T_68=$signed(_address_ok_T_66)&-33'sh10000000; 
  assign _address_ok_T_69=$signed(_address_ok_T_68)==33'sh0; 
  assign _address_ok_T_70=io_in_c_bits_address^32'h60000000; 
  assign _address_ok_T_71={1'b0,$signed(_address_ok_T_70)}; 
  assign _address_ok_T_73=$signed(_address_ok_T_71)&-33'sh20000000; 
  assign _address_ok_T_74=$signed(_address_ok_T_73)==33'sh0; 
  assign _address_ok_T_75=_address_ok_T_44|_address_ok_T_49; 
  assign _address_ok_T_76=_address_ok_T_75|_address_ok_T_54; 
  assign _address_ok_T_77=_address_ok_T_76|_address_ok_T_59; 
  assign _address_ok_T_78=_address_ok_T_77|_address_ok_T_64; 
  assign _address_ok_T_79=_address_ok_T_78|_address_ok_T_69; 
  assign address_ok_1=_address_ok_T_79|_address_ok_T_74; 
  assign _T_1483=io_in_c_bits_opcode==3'h4; 
  assign _T_1485=address_ok_1|reset; 
  assign _T_1488=source_ok_2|reset; 
  assign _T_1490=io_in_c_bits_size>=4'h3; 
  assign _T_1492=_T_1490|reset; 
  assign _T_1495=is_aligned_2|reset; 
  assign _T_1497=io_in_c_bits_param<=3'h5; 
  assign _T_1499=_T_1497|reset; 
  assign _T_1505=io_in_c_bits_opcode==3'h5; 
  assign _T_1523=io_in_c_bits_opcode==3'h6; 
  assign _T_1525=io_in_c_bits_size<=4'hc; 
  assign _T_1530=_T_1525&source_ok_2; 
  assign _T_1563=_address_ok_T_59|_address_ok_T_44; 
  assign _T_1564=_T_1563|_address_ok_T_64; 
  assign _T_1565=_T_1564|_address_ok_T_54; 
  assign _T_1566=_T_1565|_address_ok_T_49; 
  assign _T_1567=_T_1566|_address_ok_T_74; 
  assign _T_1570=io_in_c_bits_size<=4'h6; 
  assign _T_1578=_T_1570&_address_ok_T_69; 
  assign _T_1581=_T_1530&_T_1578; 
  assign _T_1583=_T_1581|reset; 
  assign _T_1587=4'h6==io_in_c_bits_size; 
  assign _T_1588=~io_in_c_bits_source&_T_1587; 
  assign _T_1635=_T_1567|_address_ok_T_69; 
  assign _T_1636=_T_1525&_T_1635; 
  assign _T_1638=_T_1588&_T_1636; 
  assign _T_1640=_T_1638|reset; 
  assign _T_1660=io_in_c_bits_opcode==3'h7; 
  assign _T_1793=io_in_c_bits_opcode==3'h0; 
  assign _T_1803=io_in_c_bits_param==3'h0; 
  assign _T_1805=_T_1803|reset; 
  assign _T_1811=io_in_c_bits_opcode==3'h1; 
  assign _T_1825=io_in_c_bits_opcode==3'h2; 
  assign _a_first_T=io_in_a_ready&io_in_a_valid; 
  assign a_first_beats1_decode=is_aligned_mask[11:3]; 
  assign a_first_beats1_opdata=~io_in_a_bits_opcode[2]; 
  assign a_first_counter1=a_first_counter-9'h1; 
  assign a_first=a_first_counter==9'h0; 
  assign _T_1847=io_in_a_valid&~a_first; 
  assign _T_1848=io_in_a_bits_opcode==opcode; 
  assign _T_1850=_T_1848|reset; 
  assign _T_1852=io_in_a_bits_param==param; 
  assign _T_1854=_T_1852|reset; 
  assign _T_1856=io_in_a_bits_size==size; 
  assign _T_1858=_T_1856|reset; 
  assign _T_1860=io_in_a_bits_source==source; 
  assign _T_1862=_T_1860|reset; 
  assign _T_1864=io_in_a_bits_address==address; 
  assign _T_1866=_T_1864|reset; 
  assign _T_1869=_a_first_T&a_first; 
  assign _d_first_T=io_in_d_ready&io_in_d_valid; 
  assign _d_first_beats1_decode_T_1=27'hfff<<io_in_d_bits_size; 
  assign d_first_beats1_decode=~_d_first_beats1_decode_T_1[11:3]; 
  assign d_first_beats1_opdata=io_in_d_bits_opcode[0]; 
  assign d_first_counter1=d_first_counter-9'h1; 
  assign d_first=d_first_counter==9'h0; 
  assign _T_1871=io_in_d_valid&~d_first; 
  assign _T_1872=io_in_d_bits_opcode==opcode_1; 
  assign _T_1874=_T_1872|reset; 
  assign _T_1876=io_in_d_bits_param==param_1; 
  assign _T_1878=_T_1876|reset; 
  assign _T_1880=io_in_d_bits_size==size_1; 
  assign _T_1882=_T_1880|reset; 
  assign _T_1884=io_in_d_bits_source==source_1; 
  assign _T_1886=_T_1884|reset; 
  assign _T_1888=io_in_d_bits_sink==sink; 
  assign _T_1890=_T_1888|reset; 
  assign _T_1892=io_in_d_bits_denied==denied; 
  assign _T_1894=_T_1892|reset; 
  assign _T_1897=_d_first_T&d_first; 
  assign b_first_done=io_in_b_ready&io_in_b_valid; 
  assign b_first_counter1=b_first_counter-9'h1; 
  assign b_first=b_first_counter==9'h0; 
  assign _T_1899=io_in_b_valid&~b_first; 
  assign _T_1900=io_in_b_bits_opcode==opcode_2; 
  assign _T_1902=_T_1900|reset; 
  assign _T_1904=io_in_b_bits_param==param_2; 
  assign _T_1906=_T_1904|reset; 
  assign _T_1908=io_in_b_bits_size==size_2; 
  assign _T_1910=_T_1908|reset; 
  assign _T_1912=io_in_b_bits_source==source_2; 
  assign _T_1914=_T_1912|reset; 
  assign _T_1916=io_in_b_bits_address==address_1; 
  assign _T_1918=_T_1916|reset; 
  assign _T_1921=b_first_done&b_first; 
  assign _c_first_T=io_in_c_ready&io_in_c_valid; 
  assign c_first_beats1_decode=is_aligned_mask_2[11:3]; 
  assign c_first_beats1_opdata=io_in_c_bits_opcode[0]; 
  assign c_first_counter1=c_first_counter-9'h1; 
  assign c_first=c_first_counter==9'h0; 
  assign _T_1923=io_in_c_valid&~c_first; 
  assign _T_1924=io_in_c_bits_opcode==opcode_3; 
  assign _T_1926=_T_1924|reset; 
  assign _T_1928=io_in_c_bits_param==param_3; 
  assign _T_1930=_T_1928|reset; 
  assign _T_1932=io_in_c_bits_size==size_3; 
  assign _T_1934=_T_1932|reset; 
  assign _T_1936=io_in_c_bits_source==source_3; 
  assign _T_1938=_T_1936|reset; 
  assign _T_1940=io_in_c_bits_address==address_2; 
  assign _T_1942=_T_1940|reset; 
  assign _T_1945=_c_first_T&c_first; 
  assign a_first_counter1_1=a_first_counter_1-9'h1; 
  assign a_first_1=a_first_counter_1==9'h0; 
  assign d_first_counter1_1=d_first_counter_1-9'h1; 
  assign d_first_1=d_first_counter_1==9'h0; 
  assign _GEN_89={io_in_d_bits_source,2'h0}; 
  assign _a_opcode_lookup_T={1'b0,_GEN_89}; 
  assign _a_opcode_lookup_T_1=inflight_opcodes>>_a_opcode_lookup_T; 
  assign _a_opcode_lookup_T_5=16'h10-16'h1; 
  assign _GEN_90={8'b0,_a_opcode_lookup_T_1}; 
  assign _a_opcode_lookup_T_6=_GEN_90&_a_opcode_lookup_T_5; 
  assign _a_opcode_lookup_T_7={1'b0,_a_opcode_lookup_T_6[15:1]}; 
  assign _a_size_lookup_T={io_in_d_bits_source,3'h0}; 
  assign _a_size_lookup_T_1=inflight_sizes>>_a_size_lookup_T; 
  assign _a_size_lookup_T_5=16'h100-16'h1; 
  assign _a_size_lookup_T_6=_a_size_lookup_T_1&_a_size_lookup_T_5; 
  assign _a_size_lookup_T_7={1'b0,_a_size_lookup_T_6[15:1]}; 
  assign _T_1946=io_in_a_valid&a_first_1; 
  assign _a_set_wo_ready_T=2'h1<<io_in_a_bits_source; 
  assign a_set_wo_ready=_T_1946 ? _a_set_wo_ready_T:2'h0; 
  assign _T_1949=_a_first_T&a_first_1; 
  assign _a_opcodes_set_interm_T={io_in_a_bits_opcode,1'h0}; 
  assign _a_opcodes_set_interm_T_1=_a_opcodes_set_interm_T|4'h1; 
  assign _a_sizes_set_interm_T={io_in_a_bits_size,1'h0}; 
  assign _a_sizes_set_interm_T_1=_a_sizes_set_interm_T|5'h1; 
  assign _GEN_93={io_in_a_bits_source,2'h0}; 
  assign _a_opcodes_set_T={1'b0,_GEN_93}; 
  assign a_opcodes_set_interm=_T_1949 ? _a_opcodes_set_interm_T_1:4'h0; 
  assign _GEN_94={15'b0,a_opcodes_set_interm}; 
  assign _a_opcodes_set_T_1=_GEN_94<<_a_opcodes_set_T; 
  assign _a_sizes_set_T={io_in_a_bits_source,3'h0}; 
  assign a_sizes_set_interm=_T_1949 ? _a_sizes_set_interm_T_1:5'h0; 
  assign _GEN_95={15'b0,a_sizes_set_interm}; 
  assign _a_sizes_set_T_1=_GEN_95<<_a_sizes_set_T; 
  assign _T_1951=inflight>>io_in_a_bits_source; 
  assign _T_1955=~_T_1951[0]|reset; 
  assign a_set=_T_1949 ? _a_set_wo_ready_T:2'h0; 
  assign _GEN_31=_T_1949 ? _a_opcodes_set_T_1:19'h0; 
  assign _GEN_32=_T_1949 ? _a_sizes_set_T_1:20'h0; 
  assign _T_1957=io_in_d_valid&d_first_1; 
  assign _T_1960=_T_1957&~_T_807; 
  assign _d_clr_wo_ready_T=2'h1<<io_in_d_bits_source; 
  assign d_clr_wo_ready=_T_1960 ? _d_clr_wo_ready_T:2'h0; 
  assign _T_1962=_d_first_T&d_first_1; 
  assign _T_1965=_T_1962&~_T_807; 
  assign _GEN_97={15'b0,_a_opcode_lookup_T_5}; 
  assign _d_opcodes_clr_T_5=_GEN_97<<_a_opcode_lookup_T; 
  assign _GEN_98={15'b0,_a_size_lookup_T_5}; 
  assign _d_sizes_clr_T_5=_GEN_98<<_a_size_lookup_T; 
  assign d_clr=_T_1965 ? _d_clr_wo_ready_T:2'h0; 
  assign _GEN_35=_T_1965 ? _d_opcodes_clr_T_5:31'h0; 
  assign _GEN_36=_T_1965 ? _d_sizes_clr_T_5:31'h0; 
  assign _same_cycle_resp_T_2=io_in_a_bits_source==io_in_d_bits_source; 
  assign same_cycle_resp=_T_1946&_same_cycle_resp_T_2; 
  assign _T_1970=inflight>>io_in_d_bits_source; 
  assign _T_1972=_T_1970[0]|same_cycle_resp; 
  assign _T_1974=_T_1972|reset; 
  assign _GEN_39=3'h2==io_in_a_bits_opcode ? 3'h1:3'h0; 
  assign _GEN_40=3'h3==io_in_a_bits_opcode ? 3'h1:_GEN_39; 
  assign _GEN_41=3'h4==io_in_a_bits_opcode ? 3'h1:_GEN_40; 
  assign _GEN_42=3'h5==io_in_a_bits_opcode ? 3'h2:_GEN_41; 
  assign _GEN_43=3'h6==io_in_a_bits_opcode ? 3'h4:_GEN_42; 
  assign _GEN_44=3'h7==io_in_a_bits_opcode ? 3'h4:_GEN_43; 
  assign _T_1976=io_in_d_bits_opcode==_GEN_44; 
  assign _GEN_51=3'h6==io_in_a_bits_opcode ? 3'h5:_GEN_42; 
  assign _GEN_52=3'h7==io_in_a_bits_opcode ? 3'h4:_GEN_51; 
  assign _T_1977=io_in_d_bits_opcode==_GEN_52; 
  assign _T_1978=_T_1976|_T_1977; 
  assign _T_1980=_T_1978|reset; 
  assign _T_1982=io_in_a_bits_size==io_in_d_bits_size; 
  assign _T_1984=_T_1982|reset; 
  assign a_opcode_lookup=_a_opcode_lookup_T_7[3:0]; 
  assign _GEN_55=3'h2==a_opcode_lookup[2:0] ? 3'h1:3'h0; 
  assign _GEN_56=3'h3==a_opcode_lookup[2:0] ? 3'h1:_GEN_55; 
  assign _GEN_57=3'h4==a_opcode_lookup[2:0] ? 3'h1:_GEN_56; 
  assign _GEN_58=3'h5==a_opcode_lookup[2:0] ? 3'h2:_GEN_57; 
  assign _GEN_59=3'h6==a_opcode_lookup[2:0] ? 3'h4:_GEN_58; 
  assign _GEN_60=3'h7==a_opcode_lookup[2:0] ? 3'h4:_GEN_59; 
  assign _T_1987=io_in_d_bits_opcode==_GEN_60; 
  assign _GEN_67=3'h6==a_opcode_lookup[2:0] ? 3'h5:_GEN_58; 
  assign _GEN_68=3'h7==a_opcode_lookup[2:0] ? 3'h4:_GEN_67; 
  assign _T_1989=io_in_d_bits_opcode==_GEN_68; 
  assign _T_1990=_T_1987|_T_1989; 
  assign _T_1992=_T_1990|reset; 
  assign a_size_lookup=_a_size_lookup_T_7[7:0]; 
  assign _GEN_99={4'b0,io_in_d_bits_size}; 
  assign _T_1994=_GEN_99==a_size_lookup; 
  assign _T_1996=_T_1994|reset; 
  assign _T_1999=_T_1957&a_first_1; 
  assign _T_2000=_T_1999&io_in_a_valid; 
  assign _T_2002=_T_2000&_same_cycle_resp_T_2; 
  assign _T_2004=_T_2002&~_T_807; 
  assign _T_2006=~io_in_d_ready|io_in_a_ready; 
  assign _T_2008=_T_2006|reset; 
  assign _T_2010=a_set_wo_ready!=d_clr_wo_ready; 
  assign _T_2011=|a_set_wo_ready; 
  assign _T_2013=_T_2010|~_T_2011; 
  assign _T_2015=_T_2013|reset; 
  assign _inflight_T=inflight|a_set; 
  assign _inflight_T_2=_inflight_T&~d_clr; 
  assign a_opcodes_set=_GEN_31[7:0]; 
  assign _inflight_opcodes_T=inflight_opcodes|a_opcodes_set; 
  assign d_opcodes_clr=_GEN_35[7:0]; 
  assign _inflight_opcodes_T_2=_inflight_opcodes_T&~d_opcodes_clr; 
  assign a_sizes_set=_GEN_32[15:0]; 
  assign _inflight_sizes_T=inflight_sizes|a_sizes_set; 
  assign d_sizes_clr=_GEN_36[15:0]; 
  assign _inflight_sizes_T_2=_inflight_sizes_T&~d_sizes_clr; 
  assign _T_2017=|inflight; 
  assign _T_2019=plusarg_reader_out==32'h0; 
  assign _T_2020=~_T_2017|_T_2019; 
  assign _T_2021=watchdog<plusarg_reader_out; 
  assign _T_2022=_T_2020|_T_2021; 
  assign _T_2024=_T_2022|reset; 
  assign _watchdog_T_1=watchdog+32'h1; 
  assign _T_2028=_a_first_T|_d_first_T; 
  assign c_first_counter1_1=c_first_counter_1-9'h1; 
  assign c_first_1=c_first_counter_1==9'h0; 
  assign d_first_counter1_2=d_first_counter_2-9'h1; 
  assign d_first_2=d_first_counter_2==9'h0; 
  assign _c_size_lookup_T_1=inflight_sizes_1>>_a_size_lookup_T; 
  assign _c_size_lookup_T_6=_c_size_lookup_T_1&_a_size_lookup_T_5; 
  assign _c_size_lookup_T_7={1'b0,_c_size_lookup_T_6[15:1]}; 
  assign _T_2029=io_in_c_valid&c_first_1; 
  assign _T_2032=io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1]; 
  assign _T_2033=_T_2029&_T_2032; 
  assign _c_set_wo_ready_T=2'h1<<io_in_c_bits_source; 
  assign c_set_wo_ready=_T_2033 ? _c_set_wo_ready_T:2'h0; 
  assign _T_2035=_c_first_T&c_first_1; 
  assign _T_2039=_T_2035&_T_2032; 
  assign _c_sizes_set_interm_T={io_in_c_bits_size,1'h0}; 
  assign _c_sizes_set_interm_T_1=_c_sizes_set_interm_T|5'h1; 
  assign _c_sizes_set_T={io_in_c_bits_source,3'h0}; 
  assign c_sizes_set_interm=_T_2039 ? _c_sizes_set_interm_T_1:5'h0; 
  assign _GEN_106={15'b0,c_sizes_set_interm}; 
  assign _c_sizes_set_T_1=_GEN_106<<_c_sizes_set_T; 
  assign _T_2040=inflight_1>>io_in_c_bits_source; 
  assign _T_2044=~_T_2040[0]|reset; 
  assign c_set=_T_2039 ? _c_set_wo_ready_T:2'h0; 
  assign _GEN_77=_T_2039 ? _c_sizes_set_T_1:20'h0; 
  assign _T_2046=io_in_d_valid&d_first_2; 
  assign _T_2048=_T_2046&_T_807; 
  assign d_clr_wo_ready_1=_T_2048 ? _d_clr_wo_ready_T:2'h0; 
  assign _T_2050=_d_first_T&d_first_2; 
  assign _T_2052=_T_2050&_T_807; 
  assign d_clr_1=_T_2052 ? _d_clr_wo_ready_T:2'h0; 
  assign _GEN_81=_T_2052 ? _d_sizes_clr_T_5:31'h0; 
  assign _same_cycle_resp_T_8=io_in_c_bits_source==io_in_d_bits_source; 
  assign same_cycle_resp_1=_T_2033&_same_cycle_resp_T_8; 
  assign _T_2056=inflight_1>>io_in_d_bits_source; 
  assign _T_2058=_T_2056[0]|same_cycle_resp_1; 
  assign _T_2060=_T_2058|reset; 
  assign _T_2062=io_in_d_bits_size==io_in_c_bits_size; 
  assign _T_2064=_T_2062|reset; 
  assign c_size_lookup=_c_size_lookup_T_7[7:0]; 
  assign _T_2066=_GEN_99==c_size_lookup; 
  assign _T_2068=_T_2066|reset; 
  assign _T_2071=_T_2046&c_first_1; 
  assign _T_2072=_T_2071&io_in_c_valid; 
  assign _T_2074=_T_2072&_same_cycle_resp_T_8; 
  assign _T_2075=_T_2074&_T_807; 
  assign _T_2077=~io_in_d_ready|io_in_c_ready; 
  assign _T_2079=_T_2077|reset; 
  assign _T_2081=|c_set_wo_ready; 
  assign _T_2082=c_set_wo_ready!=d_clr_wo_ready_1; 
  assign _T_2084=_T_2082|reset; 
  assign _inflight_T_3=inflight_1|c_set; 
  assign _inflight_T_5=_inflight_T_3&~d_clr_1; 
  assign c_sizes_set=_GEN_77[15:0]; 
  assign _inflight_sizes_T_3=inflight_sizes_1|c_sizes_set; 
  assign d_sizes_clr_1=_GEN_81[15:0]; 
  assign _inflight_sizes_T_5=_inflight_sizes_T_3&~d_sizes_clr_1; 
  assign _T_2086=|inflight_1; 
  assign _T_2088=plusarg_reader_1_out==32'h0; 
  assign _T_2089=~_T_2086|_T_2088; 
  assign _T_2090=watchdog_1<plusarg_reader_1_out; 
  assign _T_2091=_T_2089|_T_2090; 
  assign _T_2093=_T_2091|reset; 
  assign _watchdog_T_3=watchdog_1+32'h1; 
  assign _T_2097=_c_first_T|_d_first_T; 
  assign d_first_counter1_3=d_first_counter_3-9'h1; 
  assign d_first_3=d_first_counter_3==9'h0; 
  assign _T_2099=_d_first_T&d_first_3; 
  assign _T_2103=io_in_d_bits_opcode[2]&~io_in_d_bits_opcode[1]; 
  assign _T_2104=_T_2099&_T_2103; 
  assign _d_set_T=4'h1<<io_in_d_bits_sink; 
  assign _T_2105=inflight_2>>io_in_d_bits_sink; 
  assign _T_2109=~_T_2105[0]|reset; 
  assign d_set=_T_2104 ? _d_set_T:4'h0; 
  assign _T_2111=io_in_e_ready&io_in_e_valid; 
  assign _e_clr_T=4'h1<<io_in_e_bits_sink; 
  assign _T_2114=d_set|inflight_2; 
  assign _T_2115=_T_2114>>io_in_e_bits_sink; 
  assign _T_2118=_T_2115[0]|reset; 
  assign e_clr=_T_2111 ? _e_clr_T:4'h0; 
  assign _inflight_T_6=inflight_2|d_set; 
  assign _inflight_T_8=_inflight_T_6&~e_clr; 
  assign _GEN_111=io_in_a_valid&_T_24; 
  assign _GEN_125=io_in_a_valid&_T_166; 
  assign _GEN_141=io_in_a_valid&_T_312; 
  assign _GEN_153=io_in_a_valid&_T_397; 
  assign _GEN_163=io_in_a_valid&_T_483; 
  assign _GEN_173=io_in_a_valid&_T_571; 
  assign _GEN_183=io_in_a_valid&_T_647; 
  assign _GEN_193=io_in_a_valid&_T_723; 
  assign _GEN_203=io_in_d_valid&_T_807; 
  assign _GEN_213=io_in_d_valid&_T_827; 
  assign _GEN_223=io_in_d_valid&_T_855; 
  assign _GEN_233=io_in_d_valid&_T_884; 
  assign _GEN_239=io_in_d_valid&_T_901; 
  assign _GEN_245=io_in_d_valid&_T_919; 
  assign _GEN_251=io_in_b_valid&_T_960; 
  assign _GEN_265=io_in_b_valid&_T_1039; 
  assign _GEN_279=io_in_b_valid&_T_1112; 
  assign _GEN_291=io_in_b_valid&_T_1181; 
  assign _GEN_303=io_in_b_valid&_T_1252; 
  assign _GEN_313=io_in_b_valid&_T_1321; 
  assign _GEN_323=io_in_b_valid&_T_1390; 
  assign _GEN_335=io_in_c_valid&_T_1483; 
  assign _GEN_345=io_in_c_valid&_T_1505; 
  assign _GEN_355=io_in_c_valid&_T_1523; 
  assign _GEN_367=io_in_c_valid&_T_1660; 
  assign _GEN_379=io_in_c_valid&_T_1793; 
  assign _GEN_387=io_in_c_valid&_T_1811; 
  assign _GEN_395=io_in_c_valid&_T_1825; 
  assign _GEN_403=_T_1960&same_cycle_resp; 
  assign _GEN_408=_T_1960&~same_cycle_resp; 
  assign _GEN_415=_T_2048&same_cycle_resp_1; 
  assign _GEN_418=_T_2048&~same_cycle_resp_1; 
  assign TLMonitor_23_covSum=30'h0; 
  assign io_covSum=TLMonitor_23_covSum; 
  assign stopEn0=_GEN_111&~_T_84; 
  assign stopEn1=_GEN_111&~_T_141; 
  assign stopEn2=_GEN_111&~_T_144; 
  assign stopEn3=_GEN_111&~_T_148; 
  assign stopEn4=_GEN_111&~_T_151; 
  assign stopEn5=_GEN_111&~_T_155; 
  assign stopEn6=_GEN_111&~_T_160; 
  assign stopEn7=_GEN_125&~_T_84; 
  assign stopEn8=_GEN_125&~_T_141; 
  assign stopEn9=_GEN_125&~_T_144; 
  assign stopEn10=_GEN_125&~_T_148; 
  assign stopEn11=_GEN_125&~_T_151; 
  assign stopEn12=_GEN_125&~_T_155; 
  assign stopEn13=_GEN_125&~_T_301; 
  assign stopEn14=_GEN_125&~_T_160; 
  assign stopEn15=_GEN_141&~_T_322; 
  assign stopEn16=_GEN_141&~_T_377; 
  assign stopEn17=_GEN_141&~_T_144; 
  assign stopEn18=_GEN_141&~_T_151; 
  assign stopEn19=_GEN_141&~_T_387; 
  assign stopEn20=_GEN_141&~_T_391; 
  assign stopEn21=_GEN_153&~_T_467; 
  assign stopEn22=_GEN_153&~_T_144; 
  assign stopEn23=_GEN_153&~_T_151; 
  assign stopEn24=_GEN_153&~_T_387; 
  assign stopEn25=_GEN_153&~_T_391; 
  assign stopEn26=_GEN_163&~_T_467; 
  assign stopEn27=_GEN_163&~_T_144; 
  assign stopEn28=_GEN_163&~_T_151; 
  assign stopEn29=_GEN_163&~_T_387; 
  assign stopEn30=_GEN_163&~_T_569; 
  assign stopEn31=_GEN_173&~_T_631; 
  assign stopEn32=_GEN_173&~_T_144; 
  assign stopEn33=_GEN_173&~_T_151; 
  assign stopEn34=_GEN_173&~_T_641; 
  assign stopEn35=_GEN_173&~_T_391; 
  assign stopEn36=_GEN_183&~_T_631; 
  assign stopEn37=_GEN_183&~_T_144; 
  assign stopEn38=_GEN_183&~_T_151; 
  assign stopEn39=_GEN_183&~_T_717; 
  assign stopEn40=_GEN_183&~_T_391; 
  assign stopEn41=_GEN_193&~_T_783; 
  assign stopEn42=_GEN_193&~_T_144; 
  assign stopEn43=_GEN_193&~_T_151; 
  assign stopEn44=_GEN_193&~_T_793; 
  assign stopEn45=_GEN_193&~_T_391; 
  assign stopEn46=io_in_d_valid&~_T_805; 
  assign stopEn47=_GEN_203&~_T_809; 
  assign stopEn48=_GEN_203&~_T_813; 
  assign stopEn49=_GEN_203&~_T_817; 
  assign stopEn50=_GEN_203&~_T_821; 
  assign stopEn51=_GEN_203&~_T_825; 
  assign stopEn52=_GEN_213&~_T_809; 
  assign stopEn53=_GEN_213&~_T_813; 
  assign stopEn54=_GEN_213&~_T_840; 
  assign stopEn55=_GEN_213&~_T_844; 
  assign stopEn56=_GEN_213&~_T_821; 
  assign stopEn57=_GEN_223&~_T_809; 
  assign stopEn58=_GEN_223&~_T_813; 
  assign stopEn59=_GEN_223&~_T_840; 
  assign stopEn60=_GEN_223&~_T_844; 
  assign stopEn61=_GEN_223&~_T_877; 
  assign stopEn62=_GEN_233&~_T_809; 
  assign stopEn63=_GEN_233&~_T_817; 
  assign stopEn64=_GEN_233&~_T_821; 
  assign stopEn65=_GEN_239&~_T_809; 
  assign stopEn66=_GEN_239&~_T_817; 
  assign stopEn67=_GEN_239&~_T_877; 
  assign stopEn68=_GEN_245&~_T_809; 
  assign stopEn69=_GEN_245&~_T_817; 
  assign stopEn70=_GEN_245&~_T_821; 
  assign stopEn71=io_in_b_valid&~_T_938; 
  assign stopEn72=_GEN_251&~_T_1016; 
  assign stopEn73=_GEN_251&~_T_1019; 
  assign stopEn74=_GEN_251&~_T_1022; 
  assign stopEn75=_GEN_251&~_T_1025; 
  assign stopEn76=_GEN_251&~_T_1029; 
  assign stopEn77=_GEN_251&~_T_1033; 
  assign stopEn78=_GEN_251&~_T_1037; 
  assign stopEn79=_GEN_265&~reset; 
  assign stopEn80=_GEN_265&~_T_1019; 
  assign stopEn81=_GEN_265&~_T_1022; 
  assign stopEn82=_GEN_265&~_T_1025; 
  assign stopEn83=_GEN_265&~_T_1102; 
  assign stopEn84=_GEN_265&~_T_1033; 
  assign stopEn85=_GEN_265&~_T_1037; 
  assign stopEn86=_GEN_279&~reset; 
  assign stopEn87=_GEN_279&~_T_1019; 
  assign stopEn88=_GEN_279&~_T_1022; 
  assign stopEn89=_GEN_279&~_T_1025; 
  assign stopEn90=_GEN_279&~_T_1102; 
  assign stopEn91=_GEN_279&~_T_1033; 
  assign stopEn92=_GEN_291&~reset; 
  assign stopEn93=_GEN_291&~_T_1019; 
  assign stopEn94=_GEN_291&~_T_1022; 
  assign stopEn95=_GEN_291&~_T_1025; 
  assign stopEn96=_GEN_291&~_T_1102; 
  assign stopEn97=_GEN_291&~_T_1250; 
  assign stopEn98=_GEN_303&~reset; 
  assign stopEn99=_GEN_303&~_T_1019; 
  assign stopEn100=_GEN_303&~_T_1022; 
  assign stopEn101=_GEN_303&~_T_1025; 
  assign stopEn102=_GEN_303&~_T_1033; 
  assign stopEn103=_GEN_313&~reset; 
  assign stopEn104=_GEN_313&~_T_1019; 
  assign stopEn105=_GEN_313&~_T_1022; 
  assign stopEn106=_GEN_313&~_T_1025; 
  assign stopEn107=_GEN_313&~_T_1033; 
  assign stopEn108=_GEN_323&~reset; 
  assign stopEn109=_GEN_323&~_T_1019; 
  assign stopEn110=_GEN_323&~_T_1022; 
  assign stopEn111=_GEN_323&~_T_1025; 
  assign stopEn112=_GEN_323&~_T_1033; 
  assign stopEn113=_GEN_323&~_T_1037; 
  assign stopEn114=_GEN_335&~_T_1485; 
  assign stopEn115=_GEN_335&~_T_1488; 
  assign stopEn116=_GEN_335&~_T_1492; 
  assign stopEn117=_GEN_335&~_T_1495; 
  assign stopEn118=_GEN_335&~_T_1499; 
  assign stopEn119=_GEN_345&~_T_1485; 
  assign stopEn120=_GEN_345&~_T_1488; 
  assign stopEn121=_GEN_345&~_T_1492; 
  assign stopEn122=_GEN_345&~_T_1495; 
  assign stopEn123=_GEN_345&~_T_1499; 
  assign stopEn124=_GEN_355&~_T_1583; 
  assign stopEn125=_GEN_355&~_T_1640; 
  assign stopEn126=_GEN_355&~_T_1488; 
  assign stopEn127=_GEN_355&~_T_1492; 
  assign stopEn128=_GEN_355&~_T_1495; 
  assign stopEn129=_GEN_355&~_T_1499; 
  assign stopEn130=_GEN_367&~_T_1583; 
  assign stopEn131=_GEN_367&~_T_1640; 
  assign stopEn132=_GEN_367&~_T_1488; 
  assign stopEn133=_GEN_367&~_T_1492; 
  assign stopEn134=_GEN_367&~_T_1495; 
  assign stopEn135=_GEN_367&~_T_1499; 
  assign stopEn136=_GEN_379&~_T_1485; 
  assign stopEn137=_GEN_379&~_T_1488; 
  assign stopEn138=_GEN_379&~_T_1495; 
  assign stopEn139=_GEN_379&~_T_1805; 
  assign stopEn140=_GEN_387&~_T_1485; 
  assign stopEn141=_GEN_387&~_T_1488; 
  assign stopEn142=_GEN_387&~_T_1495; 
  assign stopEn143=_GEN_387&~_T_1805; 
  assign stopEn144=_GEN_395&~_T_1485; 
  assign stopEn145=_GEN_395&~_T_1488; 
  assign stopEn146=_GEN_395&~_T_1495; 
  assign stopEn147=_GEN_395&~_T_1805; 
  assign stopEn148=_T_1847&~_T_1850; 
  assign stopEn149=_T_1847&~_T_1854; 
  assign stopEn150=_T_1847&~_T_1858; 
  assign stopEn151=_T_1847&~_T_1862; 
  assign stopEn152=_T_1847&~_T_1866; 
  assign stopEn153=_T_1871&~_T_1874; 
  assign stopEn154=_T_1871&~_T_1878; 
  assign stopEn155=_T_1871&~_T_1882; 
  assign stopEn156=_T_1871&~_T_1886; 
  assign stopEn157=_T_1871&~_T_1890; 
  assign stopEn158=_T_1871&~_T_1894; 
  assign stopEn159=_T_1899&~_T_1902; 
  assign stopEn160=_T_1899&~_T_1906; 
  assign stopEn161=_T_1899&~_T_1910; 
  assign stopEn162=_T_1899&~_T_1914; 
  assign stopEn163=_T_1899&~_T_1918; 
  assign stopEn164=_T_1923&~_T_1926; 
  assign stopEn165=_T_1923&~_T_1930; 
  assign stopEn166=_T_1923&~_T_1934; 
  assign stopEn167=_T_1923&~_T_1938; 
  assign stopEn168=_T_1923&~_T_1942; 
  assign stopEn169=_T_1949&~_T_1955; 
  assign stopEn170=_T_1960&~_T_1974; 
  assign stopEn171=_GEN_403&~_T_1980; 
  assign stopEn172=_GEN_403&~_T_1984; 
  assign stopEn173=_GEN_408&~_T_1992; 
  assign stopEn174=_GEN_408&~_T_1996; 
  assign stopEn175=_T_2004&~_T_2008; 
  assign stopEn176=~_T_2015; 
  assign stopEn177=~_T_2024; 
  assign stopEn178=_T_2039&~_T_2044; 
  assign stopEn179=_T_2048&~_T_2060; 
  assign stopEn180=_GEN_415&~_T_2064; 
  assign stopEn181=_GEN_418&~_T_2068; 
  assign stopEn182=_T_2075&~_T_2079; 
  assign stopEn183=_T_2081&~_T_2084; 
  assign stopEn184=~_T_2093; 
  assign stopEn185=_T_2104&~_T_2109; 
  assign stopEn186=_T_2111&~_T_2118; 
  assign TLMonitor_23_or63=stopEn0|stopEn1; 
  assign TLMonitor_23_or130=stopEn3|stopEn4; 
  assign TLMonitor_23_or64=stopEn2|TLMonitor_23_or130; 
  assign TLMonitor_23_or31=TLMonitor_23_or63|TLMonitor_23_or64; 
  assign TLMonitor_23_or132=stopEn6|stopEn7; 
  assign TLMonitor_23_or65=stopEn5|TLMonitor_23_or132; 
  assign TLMonitor_23_or134=stopEn9|stopEn10; 
  assign TLMonitor_23_or66=stopEn8|TLMonitor_23_or134; 
  assign TLMonitor_23_or32=TLMonitor_23_or65|TLMonitor_23_or66; 
  assign TLMonitor_23_or15=TLMonitor_23_or31|TLMonitor_23_or32; 
  assign TLMonitor_23_or136=stopEn12|stopEn13; 
  assign TLMonitor_23_or67=stopEn11|TLMonitor_23_or136; 
  assign TLMonitor_23_or138=stopEn15|stopEn16; 
  assign TLMonitor_23_or68=stopEn14|TLMonitor_23_or138; 
  assign TLMonitor_23_or33=TLMonitor_23_or67|TLMonitor_23_or68; 
  assign TLMonitor_23_or140=stopEn18|stopEn19; 
  assign TLMonitor_23_or69=stopEn17|TLMonitor_23_or140; 
  assign TLMonitor_23_or142=stopEn21|stopEn22; 
  assign TLMonitor_23_or70=stopEn20|TLMonitor_23_or142; 
  assign TLMonitor_23_or34=TLMonitor_23_or69|TLMonitor_23_or70; 
  assign TLMonitor_23_or16=TLMonitor_23_or33|TLMonitor_23_or34; 
  assign TLMonitor_23_or7=TLMonitor_23_or15|TLMonitor_23_or16; 
  assign TLMonitor_23_or144=stopEn24|stopEn25; 
  assign TLMonitor_23_or71=stopEn23|TLMonitor_23_or144; 
  assign TLMonitor_23_or146=stopEn27|stopEn28; 
  assign TLMonitor_23_or72=stopEn26|TLMonitor_23_or146; 
  assign TLMonitor_23_or35=TLMonitor_23_or71|TLMonitor_23_or72; 
  assign TLMonitor_23_or148=stopEn30|stopEn31; 
  assign TLMonitor_23_or73=stopEn29|TLMonitor_23_or148; 
  assign TLMonitor_23_or150=stopEn33|stopEn34; 
  assign TLMonitor_23_or74=stopEn32|TLMonitor_23_or150; 
  assign TLMonitor_23_or36=TLMonitor_23_or73|TLMonitor_23_or74; 
  assign TLMonitor_23_or17=TLMonitor_23_or35|TLMonitor_23_or36; 
  assign TLMonitor_23_or152=stopEn36|stopEn37; 
  assign TLMonitor_23_or75=stopEn35|TLMonitor_23_or152; 
  assign TLMonitor_23_or154=stopEn39|stopEn40; 
  assign TLMonitor_23_or76=stopEn38|TLMonitor_23_or154; 
  assign TLMonitor_23_or37=TLMonitor_23_or75|TLMonitor_23_or76; 
  assign TLMonitor_23_or156=stopEn42|stopEn43; 
  assign TLMonitor_23_or77=stopEn41|TLMonitor_23_or156; 
  assign TLMonitor_23_or158=stopEn45|stopEn46; 
  assign TLMonitor_23_or78=stopEn44|TLMonitor_23_or158; 
  assign TLMonitor_23_or38=TLMonitor_23_or77|TLMonitor_23_or78; 
  assign TLMonitor_23_or18=TLMonitor_23_or37|TLMonitor_23_or38; 
  assign TLMonitor_23_or8=TLMonitor_23_or17|TLMonitor_23_or18; 
  assign TLMonitor_23_or3=TLMonitor_23_or7|TLMonitor_23_or8; 
  assign TLMonitor_23_or79=stopEn47|stopEn48; 
  assign TLMonitor_23_or162=stopEn50|stopEn51; 
  assign TLMonitor_23_or80=stopEn49|TLMonitor_23_or162; 
  assign TLMonitor_23_or39=TLMonitor_23_or79|TLMonitor_23_or80; 
  assign TLMonitor_23_or164=stopEn53|stopEn54; 
  assign TLMonitor_23_or81=stopEn52|TLMonitor_23_or164; 
  assign TLMonitor_23_or166=stopEn56|stopEn57; 
  assign TLMonitor_23_or82=stopEn55|TLMonitor_23_or166; 
  assign TLMonitor_23_or40=TLMonitor_23_or81|TLMonitor_23_or82; 
  assign TLMonitor_23_or19=TLMonitor_23_or39|TLMonitor_23_or40; 
  assign TLMonitor_23_or168=stopEn59|stopEn60; 
  assign TLMonitor_23_or83=stopEn58|TLMonitor_23_or168; 
  assign TLMonitor_23_or170=stopEn62|stopEn63; 
  assign TLMonitor_23_or84=stopEn61|TLMonitor_23_or170; 
  assign TLMonitor_23_or41=TLMonitor_23_or83|TLMonitor_23_or84; 
  assign TLMonitor_23_or172=stopEn65|stopEn66; 
  assign TLMonitor_23_or85=stopEn64|TLMonitor_23_or172; 
  assign TLMonitor_23_or174=stopEn68|stopEn69; 
  assign TLMonitor_23_or86=stopEn67|TLMonitor_23_or174; 
  assign TLMonitor_23_or42=TLMonitor_23_or85|TLMonitor_23_or86; 
  assign TLMonitor_23_or20=TLMonitor_23_or41|TLMonitor_23_or42; 
  assign TLMonitor_23_or9=TLMonitor_23_or19|TLMonitor_23_or20; 
  assign TLMonitor_23_or176=stopEn71|stopEn72; 
  assign TLMonitor_23_or87=stopEn70|TLMonitor_23_or176; 
  assign TLMonitor_23_or178=stopEn74|stopEn75; 
  assign TLMonitor_23_or88=stopEn73|TLMonitor_23_or178; 
  assign TLMonitor_23_or43=TLMonitor_23_or87|TLMonitor_23_or88; 
  assign TLMonitor_23_or180=stopEn77|stopEn78; 
  assign TLMonitor_23_or89=stopEn76|TLMonitor_23_or180; 
  assign TLMonitor_23_or182=stopEn80|stopEn81; 
  assign TLMonitor_23_or90=stopEn79|TLMonitor_23_or182; 
  assign TLMonitor_23_or44=TLMonitor_23_or89|TLMonitor_23_or90; 
  assign TLMonitor_23_or21=TLMonitor_23_or43|TLMonitor_23_or44; 
  assign TLMonitor_23_or184=stopEn83|stopEn84; 
  assign TLMonitor_23_or91=stopEn82|TLMonitor_23_or184; 
  assign TLMonitor_23_or186=stopEn86|stopEn87; 
  assign TLMonitor_23_or92=stopEn85|TLMonitor_23_or186; 
  assign TLMonitor_23_or45=TLMonitor_23_or91|TLMonitor_23_or92; 
  assign TLMonitor_23_or188=stopEn89|stopEn90; 
  assign TLMonitor_23_or93=stopEn88|TLMonitor_23_or188; 
  assign TLMonitor_23_or190=stopEn92|stopEn93; 
  assign TLMonitor_23_or94=stopEn91|TLMonitor_23_or190; 
  assign TLMonitor_23_or46=TLMonitor_23_or93|TLMonitor_23_or94; 
  assign TLMonitor_23_or22=TLMonitor_23_or45|TLMonitor_23_or46; 
  assign TLMonitor_23_or10=TLMonitor_23_or21|TLMonitor_23_or22; 
  assign TLMonitor_23_or4=TLMonitor_23_or9|TLMonitor_23_or10; 
  assign TLMonitor_23_or1=TLMonitor_23_or3|TLMonitor_23_or4; 
  assign TLMonitor_23_or95=stopEn94|stopEn95; 
  assign TLMonitor_23_or194=stopEn97|stopEn98; 
  assign TLMonitor_23_or96=stopEn96|TLMonitor_23_or194; 
  assign TLMonitor_23_or47=TLMonitor_23_or95|TLMonitor_23_or96; 
  assign TLMonitor_23_or196=stopEn100|stopEn101; 
  assign TLMonitor_23_or97=stopEn99|TLMonitor_23_or196; 
  assign TLMonitor_23_or198=stopEn103|stopEn104; 
  assign TLMonitor_23_or98=stopEn102|TLMonitor_23_or198; 
  assign TLMonitor_23_or48=TLMonitor_23_or97|TLMonitor_23_or98; 
  assign TLMonitor_23_or23=TLMonitor_23_or47|TLMonitor_23_or48; 
  assign TLMonitor_23_or200=stopEn106|stopEn107; 
  assign TLMonitor_23_or99=stopEn105|TLMonitor_23_or200; 
  assign TLMonitor_23_or202=stopEn109|stopEn110; 
  assign TLMonitor_23_or100=stopEn108|TLMonitor_23_or202; 
  assign TLMonitor_23_or49=TLMonitor_23_or99|TLMonitor_23_or100; 
  assign TLMonitor_23_or204=stopEn112|stopEn113; 
  assign TLMonitor_23_or101=stopEn111|TLMonitor_23_or204; 
  assign TLMonitor_23_or206=stopEn115|stopEn116; 
  assign TLMonitor_23_or102=stopEn114|TLMonitor_23_or206; 
  assign TLMonitor_23_or50=TLMonitor_23_or101|TLMonitor_23_or102; 
  assign TLMonitor_23_or24=TLMonitor_23_or49|TLMonitor_23_or50; 
  assign TLMonitor_23_or11=TLMonitor_23_or23|TLMonitor_23_or24; 
  assign TLMonitor_23_or208=stopEn118|stopEn119; 
  assign TLMonitor_23_or103=stopEn117|TLMonitor_23_or208; 
  assign TLMonitor_23_or210=stopEn121|stopEn122; 
  assign TLMonitor_23_or104=stopEn120|TLMonitor_23_or210; 
  assign TLMonitor_23_or51=TLMonitor_23_or103|TLMonitor_23_or104; 
  assign TLMonitor_23_or212=stopEn124|stopEn125; 
  assign TLMonitor_23_or105=stopEn123|TLMonitor_23_or212; 
  assign TLMonitor_23_or214=stopEn127|stopEn128; 
  assign TLMonitor_23_or106=stopEn126|TLMonitor_23_or214; 
  assign TLMonitor_23_or52=TLMonitor_23_or105|TLMonitor_23_or106; 
  assign TLMonitor_23_or25=TLMonitor_23_or51|TLMonitor_23_or52; 
  assign TLMonitor_23_or216=stopEn130|stopEn131; 
  assign TLMonitor_23_or107=stopEn129|TLMonitor_23_or216; 
  assign TLMonitor_23_or218=stopEn133|stopEn134; 
  assign TLMonitor_23_or108=stopEn132|TLMonitor_23_or218; 
  assign TLMonitor_23_or53=TLMonitor_23_or107|TLMonitor_23_or108; 
  assign TLMonitor_23_or220=stopEn136|stopEn137; 
  assign TLMonitor_23_or109=stopEn135|TLMonitor_23_or220; 
  assign TLMonitor_23_or222=stopEn139|stopEn140; 
  assign TLMonitor_23_or110=stopEn138|TLMonitor_23_or222; 
  assign TLMonitor_23_or54=TLMonitor_23_or109|TLMonitor_23_or110; 
  assign TLMonitor_23_or26=TLMonitor_23_or53|TLMonitor_23_or54; 
  assign TLMonitor_23_or12=TLMonitor_23_or25|TLMonitor_23_or26; 
  assign TLMonitor_23_or5=TLMonitor_23_or11|TLMonitor_23_or12; 
  assign TLMonitor_23_or224=stopEn142|stopEn143; 
  assign TLMonitor_23_or111=stopEn141|TLMonitor_23_or224; 
  assign TLMonitor_23_or226=stopEn145|stopEn146; 
  assign TLMonitor_23_or112=stopEn144|TLMonitor_23_or226; 
  assign TLMonitor_23_or55=TLMonitor_23_or111|TLMonitor_23_or112; 
  assign TLMonitor_23_or228=stopEn148|stopEn149; 
  assign TLMonitor_23_or113=stopEn147|TLMonitor_23_or228; 
  assign TLMonitor_23_or230=stopEn151|stopEn152; 
  assign TLMonitor_23_or114=stopEn150|TLMonitor_23_or230; 
  assign TLMonitor_23_or56=TLMonitor_23_or113|TLMonitor_23_or114; 
  assign TLMonitor_23_or27=TLMonitor_23_or55|TLMonitor_23_or56; 
  assign TLMonitor_23_or232=stopEn154|stopEn155; 
  assign TLMonitor_23_or115=stopEn153|TLMonitor_23_or232; 
  assign TLMonitor_23_or234=stopEn157|stopEn158; 
  assign TLMonitor_23_or116=stopEn156|TLMonitor_23_or234; 
  assign TLMonitor_23_or57=TLMonitor_23_or115|TLMonitor_23_or116; 
  assign TLMonitor_23_or236=stopEn160|stopEn161; 
  assign TLMonitor_23_or117=stopEn159|TLMonitor_23_or236; 
  assign TLMonitor_23_or238=stopEn163|stopEn164; 
  assign TLMonitor_23_or118=stopEn162|TLMonitor_23_or238; 
  assign TLMonitor_23_or58=TLMonitor_23_or117|TLMonitor_23_or118; 
  assign TLMonitor_23_or28=TLMonitor_23_or57|TLMonitor_23_or58; 
  assign TLMonitor_23_or13=TLMonitor_23_or27|TLMonitor_23_or28; 
  assign TLMonitor_23_or240=stopEn166|stopEn167; 
  assign TLMonitor_23_or119=stopEn165|TLMonitor_23_or240; 
  assign TLMonitor_23_or242=stopEn169|stopEn170; 
  assign TLMonitor_23_or120=stopEn168|TLMonitor_23_or242; 
  assign TLMonitor_23_or59=TLMonitor_23_or119|TLMonitor_23_or120; 
  assign TLMonitor_23_or244=stopEn172|stopEn173; 
  assign TLMonitor_23_or121=stopEn171|TLMonitor_23_or244; 
  assign TLMonitor_23_or246=stopEn175|stopEn176; 
  assign TLMonitor_23_or122=stopEn174|TLMonitor_23_or246; 
  assign TLMonitor_23_or60=TLMonitor_23_or121|TLMonitor_23_or122; 
  assign TLMonitor_23_or29=TLMonitor_23_or59|TLMonitor_23_or60; 
  assign TLMonitor_23_or248=stopEn178|stopEn179; 
  assign TLMonitor_23_or123=stopEn177|TLMonitor_23_or248; 
  assign TLMonitor_23_or250=stopEn181|stopEn182; 
  assign TLMonitor_23_or124=stopEn180|TLMonitor_23_or250; 
  assign TLMonitor_23_or61=TLMonitor_23_or123|TLMonitor_23_or124; 
  assign TLMonitor_23_or252=stopEn184|stopEn185; 
  assign TLMonitor_23_or125=stopEn183|TLMonitor_23_or252; 
  assign TLMonitor_23_or254=plusarg_reader_metaAssert_wire|plusarg_reader_1_metaAssert_wire; 
  assign TLMonitor_23_or126=stopEn186|TLMonitor_23_or254; 
  assign TLMonitor_23_or62=TLMonitor_23_or125|TLMonitor_23_or126; 
  assign TLMonitor_23_or30=TLMonitor_23_or61|TLMonitor_23_or62; 
  assign TLMonitor_23_or14=TLMonitor_23_or29|TLMonitor_23_or30; 
  assign TLMonitor_23_or6=TLMonitor_23_or13|TLMonitor_23_or14; 
  assign TLMonitor_23_or2=TLMonitor_23_or5|TLMonitor_23_or6; 
  assign TLMonitor_23_or0=TLMonitor_23_or1|TLMonitor_23_or2; 
  assign metaAssert=TLMonitor_23_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              a_first_counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 a_first_counter <=9'h0;
               end 
             else 
               if (_a_first_T)
                  begin 
                    if (a_first)
                       begin 
                         if (a_first_beats1_opdata)
                            begin 
                              a_first_counter <=a_first_beats1_decode;
                            end 
                          else 
                            begin 
                              a_first_counter <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         a_first_counter <=a_first_counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              opcode <=3'h0;
            end 
          else 
            if (_T_1869)
               begin 
                 opcode <=io_in_a_bits_opcode;
               end 
         if (metaReset)
            begin 
              param <=3'h0;
            end 
          else 
            if (_T_1869)
               begin 
                 param <=io_in_a_bits_param;
               end 
         if (metaReset)
            begin 
              size <=4'h0;
            end 
          else 
            if (_T_1869)
               begin 
                 size <=io_in_a_bits_size;
               end 
         if (metaReset)
            begin 
              source <=1'h0;
            end 
          else 
            if (_T_1869)
               begin 
                 source <=io_in_a_bits_source;
               end 
         if (metaReset)
            begin 
              address <=32'h0;
            end 
          else 
            if (_T_1869)
               begin 
                 address <=io_in_a_bits_address;
               end 
         if (metaReset)
            begin 
              d_first_counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 d_first_counter <=9'h0;
               end 
             else 
               if (_d_first_T)
                  begin 
                    if (d_first)
                       begin 
                         if (d_first_beats1_opdata)
                            begin 
                              d_first_counter <=d_first_beats1_decode;
                            end 
                          else 
                            begin 
                              d_first_counter <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         d_first_counter <=d_first_counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              opcode_1 <=3'h0;
            end 
          else 
            if (_T_1897)
               begin 
                 opcode_1 <=io_in_d_bits_opcode;
               end 
         if (metaReset)
            begin 
              param_1 <=2'h0;
            end 
          else 
            if (_T_1897)
               begin 
                 param_1 <=io_in_d_bits_param;
               end 
         if (metaReset)
            begin 
              size_1 <=4'h0;
            end 
          else 
            if (_T_1897)
               begin 
                 size_1 <=io_in_d_bits_size;
               end 
         if (metaReset)
            begin 
              source_1 <=1'h0;
            end 
          else 
            if (_T_1897)
               begin 
                 source_1 <=io_in_d_bits_source;
               end 
         if (metaReset)
            begin 
              sink <=2'h0;
            end 
          else 
            if (_T_1897)
               begin 
                 sink <=io_in_d_bits_sink;
               end 
         if (metaReset)
            begin 
              denied <=1'h0;
            end 
          else 
            if (_T_1897)
               begin 
                 denied <=io_in_d_bits_denied;
               end 
         if (metaReset)
            begin 
              b_first_counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 b_first_counter <=9'h0;
               end 
             else 
               if (b_first_done)
                  begin 
                    if (b_first)
                       begin 
                         b_first_counter <=9'h0;
                       end 
                     else 
                       begin 
                         b_first_counter <=b_first_counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              opcode_2 <=3'h0;
            end 
          else 
            if (_T_1921)
               begin 
                 opcode_2 <=io_in_b_bits_opcode;
               end 
         if (metaReset)
            begin 
              param_2 <=2'h0;
            end 
          else 
            if (_T_1921)
               begin 
                 param_2 <=io_in_b_bits_param;
               end 
         if (metaReset)
            begin 
              size_2 <=4'h0;
            end 
          else 
            if (_T_1921)
               begin 
                 size_2 <=io_in_b_bits_size;
               end 
         if (metaReset)
            begin 
              source_2 <=1'h0;
            end 
          else 
            if (_T_1921)
               begin 
                 source_2 <=io_in_b_bits_source;
               end 
         if (metaReset)
            begin 
              address_1 <=32'h0;
            end 
          else 
            if (_T_1921)
               begin 
                 address_1 <=io_in_b_bits_address;
               end 
         if (metaReset)
            begin 
              c_first_counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 c_first_counter <=9'h0;
               end 
             else 
               if (_c_first_T)
                  begin 
                    if (c_first)
                       begin 
                         if (c_first_beats1_opdata)
                            begin 
                              c_first_counter <=c_first_beats1_decode;
                            end 
                          else 
                            begin 
                              c_first_counter <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         c_first_counter <=c_first_counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              opcode_3 <=3'h0;
            end 
          else 
            if (_T_1945)
               begin 
                 opcode_3 <=io_in_c_bits_opcode;
               end 
         if (metaReset)
            begin 
              param_3 <=3'h0;
            end 
          else 
            if (_T_1945)
               begin 
                 param_3 <=io_in_c_bits_param;
               end 
         if (metaReset)
            begin 
              size_3 <=4'h0;
            end 
          else 
            if (_T_1945)
               begin 
                 size_3 <=io_in_c_bits_size;
               end 
         if (metaReset)
            begin 
              source_3 <=1'h0;
            end 
          else 
            if (_T_1945)
               begin 
                 source_3 <=io_in_c_bits_source;
               end 
         if (metaReset)
            begin 
              address_2 <=32'h0;
            end 
          else 
            if (_T_1945)
               begin 
                 address_2 <=io_in_c_bits_address;
               end 
         if (metaReset)
            begin 
              inflight <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight <=2'h0;
               end 
             else 
               begin 
                 inflight <=_inflight_T_2;
               end 
         if (metaReset)
            begin 
              inflight_opcodes <=8'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_opcodes <=8'h0;
               end 
             else 
               begin 
                 inflight_opcodes <=_inflight_opcodes_T_2;
               end 
         if (metaReset)
            begin 
              inflight_sizes <=16'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_sizes <=16'h0;
               end 
             else 
               begin 
                 inflight_sizes <=_inflight_sizes_T_2;
               end 
         if (metaReset)
            begin 
              a_first_counter_1 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 a_first_counter_1 <=9'h0;
               end 
             else 
               if (_a_first_T)
                  begin 
                    if (a_first_1)
                       begin 
                         if (a_first_beats1_opdata)
                            begin 
                              a_first_counter_1 <=a_first_beats1_decode;
                            end 
                          else 
                            begin 
                              a_first_counter_1 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         a_first_counter_1 <=a_first_counter1_1;
                       end 
                  end 
         if (metaReset)
            begin 
              d_first_counter_1 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 d_first_counter_1 <=9'h0;
               end 
             else 
               if (_d_first_T)
                  begin 
                    if (d_first_1)
                       begin 
                         if (d_first_beats1_opdata)
                            begin 
                              d_first_counter_1 <=d_first_beats1_decode;
                            end 
                          else 
                            begin 
                              d_first_counter_1 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         d_first_counter_1 <=d_first_counter1_1;
                       end 
                  end 
         if (metaReset)
            begin 
              watchdog <=32'h0;
            end 
          else 
            if (reset)
               begin 
                 watchdog <=32'h0;
               end 
             else 
               if (_T_2028)
                  begin 
                    watchdog <=32'h0;
                  end 
                else 
                  begin 
                    watchdog <=_watchdog_T_1;
                  end 
         if (metaReset)
            begin 
              inflight_1 <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_1 <=2'h0;
               end 
             else 
               begin 
                 inflight_1 <=_inflight_T_5;
               end 
         if (metaReset)
            begin 
              inflight_sizes_1 <=16'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_sizes_1 <=16'h0;
               end 
             else 
               begin 
                 inflight_sizes_1 <=_inflight_sizes_T_5;
               end 
         if (metaReset)
            begin 
              c_first_counter_1 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 c_first_counter_1 <=9'h0;
               end 
             else 
               if (_c_first_T)
                  begin 
                    if (c_first_1)
                       begin 
                         if (c_first_beats1_opdata)
                            begin 
                              c_first_counter_1 <=c_first_beats1_decode;
                            end 
                          else 
                            begin 
                              c_first_counter_1 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         c_first_counter_1 <=c_first_counter1_1;
                       end 
                  end 
         if (metaReset)
            begin 
              d_first_counter_2 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 d_first_counter_2 <=9'h0;
               end 
             else 
               if (_d_first_T)
                  begin 
                    if (d_first_2)
                       begin 
                         if (d_first_beats1_opdata)
                            begin 
                              d_first_counter_2 <=d_first_beats1_decode;
                            end 
                          else 
                            begin 
                              d_first_counter_2 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         d_first_counter_2 <=d_first_counter1_2;
                       end 
                  end 
         if (metaReset)
            begin 
              watchdog_1 <=32'h0;
            end 
          else 
            if (reset)
               begin 
                 watchdog_1 <=32'h0;
               end 
             else 
               if (_T_2097)
                  begin 
                    watchdog_1 <=32'h0;
                  end 
                else 
                  begin 
                    watchdog_1 <=_watchdog_T_3;
                  end 
         if (metaReset)
            begin 
              inflight_2 <=4'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_2 <=4'h0;
               end 
             else 
               begin 
                 inflight_2 <=_inflight_T_8;
               end 
         if (metaReset)
            begin 
              d_first_counter_3 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 d_first_counter_3 <=9'h0;
               end 
             else 
               if (_d_first_T)
                  begin 
                    if (d_first_3)
                       begin 
                         if (d_first_beats1_opdata)
                            begin 
                              d_first_counter_3 <=d_first_beats1_decode;
                            end 
                          else 
                            begin 
                              d_first_counter_3 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         d_first_counter_3 <=d_first_counter1_3;
                       end 
                  end 
         if (_GEN_111&~_T_84)
            begin $display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_111&~_T_84)
            begin $display("fatal");
            end 
         if (_GEN_111&~_T_141)
            begin $display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_111&~_T_141)
            begin $display("fatal");
            end 
         if (_GEN_111&~_T_144)
            begin $display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_111&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_111&~_T_148)
            begin $display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_111&~_T_148)
            begin $display("fatal");
            end 
         if (_GEN_111&~_T_151)
            begin $display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_111&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_111&~_T_155)
            begin $display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_111&~_T_155)
            begin $display("fatal");
            end 
         if (_GEN_111&~_T_160)
            begin $display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_111&~_T_160)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_84)
            begin $display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_84)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_141)
            begin $display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_141)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_144)
            begin $display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_148)
            begin $display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_148)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_151)
            begin $display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_155)
            begin $display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_155)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_301)
            begin $display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_301)
            begin $display("fatal");
            end 
         if (_GEN_125&~_T_160)
            begin $display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_125&~_T_160)
            begin $display("fatal");
            end 
         if (_GEN_141&~_T_322)
            begin $display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_141&~_T_322)
            begin $display("fatal");
            end 
         if (_GEN_141&~_T_377)
            begin $display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_141&~_T_377)
            begin $display("fatal");
            end 
         if (_GEN_141&~_T_144)
            begin $display("Assertion failed: 'A' channel Get carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_141&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_141&~_T_151)
            begin $display("Assertion failed: 'A' channel Get address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_141&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_141&~_T_387)
            begin $display("Assertion failed: 'A' channel Get carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_141&~_T_387)
            begin $display("fatal");
            end 
         if (_GEN_141&~_T_391)
            begin $display("Assertion failed: 'A' channel Get contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_141&~_T_391)
            begin $display("fatal");
            end 
         if (_GEN_153&~_T_467)
            begin $display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_153&~_T_467)
            begin $display("fatal");
            end 
         if (_GEN_153&~_T_144)
            begin $display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_153&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_153&~_T_151)
            begin $display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_153&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_153&~_T_387)
            begin $display("Assertion failed: 'A' channel PutFull carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_153&~_T_387)
            begin $display("fatal");
            end 
         if (_GEN_153&~_T_391)
            begin $display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_153&~_T_391)
            begin $display("fatal");
            end 
         if (_GEN_163&~_T_467)
            begin $display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_163&~_T_467)
            begin $display("fatal");
            end 
         if (_GEN_163&~_T_144)
            begin $display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_163&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_163&~_T_151)
            begin $display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_163&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_163&~_T_387)
            begin $display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_163&~_T_387)
            begin $display("fatal");
            end 
         if (_GEN_163&~_T_569)
            begin $display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_163&~_T_569)
            begin $display("fatal");
            end 
         if (_GEN_173&~_T_631)
            begin $display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_173&~_T_631)
            begin $display("fatal");
            end 
         if (_GEN_173&~_T_144)
            begin $display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_173&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_173&~_T_151)
            begin $display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_173&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_173&~_T_641)
            begin $display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_173&~_T_641)
            begin $display("fatal");
            end 
         if (_GEN_173&~_T_391)
            begin $display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_173&~_T_391)
            begin $display("fatal");
            end 
         if (_GEN_183&~_T_631)
            begin $display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_183&~_T_631)
            begin $display("fatal");
            end 
         if (_GEN_183&~_T_144)
            begin $display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_183&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_183&~_T_151)
            begin $display("Assertion failed: 'A' channel Logical address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_183&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_183&~_T_717)
            begin $display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_183&~_T_717)
            begin $display("fatal");
            end 
         if (_GEN_183&~_T_391)
            begin $display("Assertion failed: 'A' channel Logical contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_183&~_T_391)
            begin $display("fatal");
            end 
         if (_GEN_193&~_T_783)
            begin $display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_193&~_T_783)
            begin $display("fatal");
            end 
         if (_GEN_193&~_T_144)
            begin $display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_193&~_T_144)
            begin $display("fatal");
            end 
         if (_GEN_193&~_T_151)
            begin $display("Assertion failed: 'A' channel Hint address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_193&~_T_151)
            begin $display("fatal");
            end 
         if (_GEN_193&~_T_793)
            begin $display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_193&~_T_793)
            begin $display("fatal");
            end 
         if (_GEN_193&~_T_391)
            begin $display("Assertion failed: 'A' channel Hint contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_193&~_T_391)
            begin $display("fatal");
            end 
         if (io_in_d_valid&~_T_805)
            begin $display("Assertion failed: 'D' channel has invalid opcode (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (io_in_d_valid&~_T_805)
            begin $display("fatal");
            end 
         if (_GEN_203&~_T_809)
            begin $display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_203&~_T_809)
            begin $display("fatal");
            end 
         if (_GEN_203&~_T_813)
            begin $display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_203&~_T_813)
            begin $display("fatal");
            end 
         if (_GEN_203&~_T_817)
            begin $display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_203&~_T_817)
            begin $display("fatal");
            end 
         if (_GEN_203&~_T_821)
            begin $display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_203&~_T_821)
            begin $display("fatal");
            end 
         if (_GEN_203&~_T_825)
            begin $display("Assertion failed: 'D' channel ReleaseAck is denied (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_203&~_T_825)
            begin $display("fatal");
            end 
         if (_GEN_213&~_T_809)
            begin $display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_213&~_T_809)
            begin $display("fatal");
            end 
         if (_GEN_213&~_T_813)
            begin $display("Assertion failed: 'D' channel Grant smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_213&~_T_813)
            begin $display("fatal");
            end 
         if (_GEN_213&~_T_840)
            begin $display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_213&~_T_840)
            begin $display("fatal");
            end 
         if (_GEN_213&~_T_844)
            begin $display("Assertion failed: 'D' channel Grant carries toN param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_213&~_T_844)
            begin $display("fatal");
            end 
         if (_GEN_213&~_T_821)
            begin $display("Assertion failed: 'D' channel Grant is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_213&~_T_821)
            begin $display("fatal");
            end 
         if (_GEN_223&~_T_809)
            begin $display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_223&~_T_809)
            begin $display("fatal");
            end 
         if (_GEN_223&~_T_813)
            begin $display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_223&~_T_813)
            begin $display("fatal");
            end 
         if (_GEN_223&~_T_840)
            begin $display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_223&~_T_840)
            begin $display("fatal");
            end 
         if (_GEN_223&~_T_844)
            begin $display("Assertion failed: 'D' channel GrantData carries toN param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_223&~_T_844)
            begin $display("fatal");
            end 
         if (_GEN_223&~_T_877)
            begin $display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_223&~_T_877)
            begin $display("fatal");
            end 
         if (_GEN_233&~_T_809)
            begin $display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_233&~_T_809)
            begin $display("fatal");
            end 
         if (_GEN_233&~_T_817)
            begin $display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_233&~_T_817)
            begin $display("fatal");
            end 
         if (_GEN_233&~_T_821)
            begin $display("Assertion failed: 'D' channel AccessAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_233&~_T_821)
            begin $display("fatal");
            end 
         if (_GEN_239&~_T_809)
            begin $display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_239&~_T_809)
            begin $display("fatal");
            end 
         if (_GEN_239&~_T_817)
            begin $display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_239&~_T_817)
            begin $display("fatal");
            end 
         if (_GEN_239&~_T_877)
            begin $display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_239&~_T_877)
            begin $display("fatal");
            end 
         if (_GEN_245&~_T_809)
            begin $display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_245&~_T_809)
            begin $display("fatal");
            end 
         if (_GEN_245&~_T_817)
            begin $display("Assertion failed: 'D' channel HintAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_245&~_T_817)
            begin $display("fatal");
            end 
         if (_GEN_245&~_T_821)
            begin $display("Assertion failed: 'D' channel HintAck is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_245&~_T_821)
            begin $display("fatal");
            end 
         if (io_in_b_valid&~_T_938)
            begin $display("Assertion failed: 'B' channel has invalid opcode (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (io_in_b_valid&~_T_938)
            begin $display("fatal");
            end 
         if (_GEN_251&~_T_1016)
            begin $display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_251&~_T_1016)
            begin $display("fatal");
            end 
         if (_GEN_251&~_T_1019)
            begin $display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_251&~_T_1019)
            begin $display("fatal");
            end 
         if (_GEN_251&~_T_1022)
            begin $display("Assertion failed: 'B' channel Probe carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_251&~_T_1022)
            begin $display("fatal");
            end 
         if (_GEN_251&~_T_1025)
            begin $display("Assertion failed: 'B' channel Probe address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_251&~_T_1025)
            begin $display("fatal");
            end 
         if (_GEN_251&~_T_1029)
            begin $display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_251&~_T_1029)
            begin $display("fatal");
            end 
         if (_GEN_251&~_T_1033)
            begin $display("Assertion failed: 'B' channel Probe contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_251&~_T_1033)
            begin $display("fatal");
            end 
         if (_GEN_251&~_T_1037)
            begin $display("Assertion failed: 'B' channel Probe is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_251&~_T_1037)
            begin $display("fatal");
            end 
         if (_GEN_265&~reset)
            begin $display("Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_265&~reset)
            begin $display("fatal");
            end 
         if (_GEN_265&~_T_1019)
            begin $display("Assertion failed: 'B' channel Get carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_265&~_T_1019)
            begin $display("fatal");
            end 
         if (_GEN_265&~_T_1022)
            begin $display("Assertion failed: 'B' channel Get carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_265&~_T_1022)
            begin $display("fatal");
            end 
         if (_GEN_265&~_T_1025)
            begin $display("Assertion failed: 'B' channel Get address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_265&~_T_1025)
            begin $display("fatal");
            end 
         if (_GEN_265&~_T_1102)
            begin $display("Assertion failed: 'B' channel Get carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_265&~_T_1102)
            begin $display("fatal");
            end 
         if (_GEN_265&~_T_1033)
            begin $display("Assertion failed: 'B' channel Get contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_265&~_T_1033)
            begin $display("fatal");
            end 
         if (_GEN_265&~_T_1037)
            begin $display("Assertion failed: 'B' channel Get is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_265&~_T_1037)
            begin $display("fatal");
            end 
         if (_GEN_279&~reset)
            begin $display("Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_279&~reset)
            begin $display("fatal");
            end 
         if (_GEN_279&~_T_1019)
            begin $display("Assertion failed: 'B' channel PutFull carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_279&~_T_1019)
            begin $display("fatal");
            end 
         if (_GEN_279&~_T_1022)
            begin $display("Assertion failed: 'B' channel PutFull carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_279&~_T_1022)
            begin $display("fatal");
            end 
         if (_GEN_279&~_T_1025)
            begin $display("Assertion failed: 'B' channel PutFull address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_279&~_T_1025)
            begin $display("fatal");
            end 
         if (_GEN_279&~_T_1102)
            begin $display("Assertion failed: 'B' channel PutFull carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_279&~_T_1102)
            begin $display("fatal");
            end 
         if (_GEN_279&~_T_1033)
            begin $display("Assertion failed: 'B' channel PutFull contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_279&~_T_1033)
            begin $display("fatal");
            end 
         if (_GEN_291&~reset)
            begin $display("Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_291&~reset)
            begin $display("fatal");
            end 
         if (_GEN_291&~_T_1019)
            begin $display("Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_291&~_T_1019)
            begin $display("fatal");
            end 
         if (_GEN_291&~_T_1022)
            begin $display("Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_291&~_T_1022)
            begin $display("fatal");
            end 
         if (_GEN_291&~_T_1025)
            begin $display("Assertion failed: 'B' channel PutPartial address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_291&~_T_1025)
            begin $display("fatal");
            end 
         if (_GEN_291&~_T_1102)
            begin $display("Assertion failed: 'B' channel PutPartial carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_291&~_T_1102)
            begin $display("fatal");
            end 
         if (_GEN_291&~_T_1250)
            begin $display("Assertion failed: 'B' channel PutPartial contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_291&~_T_1250)
            begin $display("fatal");
            end 
         if (_GEN_303&~reset)
            begin $display("Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_303&~reset)
            begin $display("fatal");
            end 
         if (_GEN_303&~_T_1019)
            begin $display("Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_303&~_T_1019)
            begin $display("fatal");
            end 
         if (_GEN_303&~_T_1022)
            begin $display("Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_303&~_T_1022)
            begin $display("fatal");
            end 
         if (_GEN_303&~_T_1025)
            begin $display("Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_303&~_T_1025)
            begin $display("fatal");
            end 
         if (_GEN_303&~_T_1033)
            begin $display("Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_303&~_T_1033)
            begin $display("fatal");
            end 
         if (_GEN_313&~reset)
            begin $display("Assertion failed: 'B' channel carries Logical type unsupported by client (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_313&~reset)
            begin $display("fatal");
            end 
         if (_GEN_313&~_T_1019)
            begin $display("Assertion failed: 'B' channel Logical carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_313&~_T_1019)
            begin $display("fatal");
            end 
         if (_GEN_313&~_T_1022)
            begin $display("Assertion failed: 'B' channel Logical carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_313&~_T_1022)
            begin $display("fatal");
            end 
         if (_GEN_313&~_T_1025)
            begin $display("Assertion failed: 'B' channel Logical address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_313&~_T_1025)
            begin $display("fatal");
            end 
         if (_GEN_313&~_T_1033)
            begin $display("Assertion failed: 'B' channel Logical contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_313&~_T_1033)
            begin $display("fatal");
            end 
         if (_GEN_323&~reset)
            begin $display("Assertion failed: 'B' channel carries Hint type unsupported by client (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_323&~reset)
            begin $display("fatal");
            end 
         if (_GEN_323&~_T_1019)
            begin $display("Assertion failed: 'B' channel Hint carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_323&~_T_1019)
            begin $display("fatal");
            end 
         if (_GEN_323&~_T_1022)
            begin $display("Assertion failed: 'B' channel Hint carries source that is not first source (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_323&~_T_1022)
            begin $display("fatal");
            end 
         if (_GEN_323&~_T_1025)
            begin $display("Assertion failed: 'B' channel Hint address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_323&~_T_1025)
            begin $display("fatal");
            end 
         if (_GEN_323&~_T_1033)
            begin $display("Assertion failed: 'B' channel Hint contains invalid mask (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_323&~_T_1033)
            begin $display("fatal");
            end 
         if (_GEN_323&~_T_1037)
            begin $display("Assertion failed: 'B' channel Hint is corrupt (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_323&~_T_1037)
            begin $display("fatal");
            end 
         if (_GEN_335&~_T_1485)
            begin $display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_335&~_T_1485)
            begin $display("fatal");
            end 
         if (_GEN_335&~_T_1488)
            begin $display("Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_335&~_T_1488)
            begin $display("fatal");
            end 
         if (_GEN_335&~_T_1492)
            begin $display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_335&~_T_1492)
            begin $display("fatal");
            end 
         if (_GEN_335&~_T_1495)
            begin $display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_335&~_T_1495)
            begin $display("fatal");
            end 
         if (_GEN_335&~_T_1499)
            begin $display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_335&~_T_1499)
            begin $display("fatal");
            end 
         if (_GEN_345&~_T_1485)
            begin $display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_345&~_T_1485)
            begin $display("fatal");
            end 
         if (_GEN_345&~_T_1488)
            begin $display("Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_345&~_T_1488)
            begin $display("fatal");
            end 
         if (_GEN_345&~_T_1492)
            begin $display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_345&~_T_1492)
            begin $display("fatal");
            end 
         if (_GEN_345&~_T_1495)
            begin $display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_345&~_T_1495)
            begin $display("fatal");
            end 
         if (_GEN_345&~_T_1499)
            begin $display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_345&~_T_1499)
            begin $display("fatal");
            end 
         if (_GEN_355&~_T_1583)
            begin $display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_355&~_T_1583)
            begin $display("fatal");
            end 
         if (_GEN_355&~_T_1640)
            begin $display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_355&~_T_1640)
            begin $display("fatal");
            end 
         if (_GEN_355&~_T_1488)
            begin $display("Assertion failed: 'C' channel Release carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_355&~_T_1488)
            begin $display("fatal");
            end 
         if (_GEN_355&~_T_1492)
            begin $display("Assertion failed: 'C' channel Release smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_355&~_T_1492)
            begin $display("fatal");
            end 
         if (_GEN_355&~_T_1495)
            begin $display("Assertion failed: 'C' channel Release address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_355&~_T_1495)
            begin $display("fatal");
            end 
         if (_GEN_355&~_T_1499)
            begin $display("Assertion failed: 'C' channel Release carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_355&~_T_1499)
            begin $display("fatal");
            end 
         if (_GEN_367&~_T_1583)
            begin $display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_367&~_T_1583)
            begin $display("fatal");
            end 
         if (_GEN_367&~_T_1640)
            begin $display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_367&~_T_1640)
            begin $display("fatal");
            end 
         if (_GEN_367&~_T_1488)
            begin $display("Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_367&~_T_1488)
            begin $display("fatal");
            end 
         if (_GEN_367&~_T_1492)
            begin $display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_367&~_T_1492)
            begin $display("fatal");
            end 
         if (_GEN_367&~_T_1495)
            begin $display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_367&~_T_1495)
            begin $display("fatal");
            end 
         if (_GEN_367&~_T_1499)
            begin $display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_367&~_T_1499)
            begin $display("fatal");
            end 
         if (_GEN_379&~_T_1485)
            begin $display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_379&~_T_1485)
            begin $display("fatal");
            end 
         if (_GEN_379&~_T_1488)
            begin $display("Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_379&~_T_1488)
            begin $display("fatal");
            end 
         if (_GEN_379&~_T_1495)
            begin $display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_379&~_T_1495)
            begin $display("fatal");
            end 
         if (_GEN_379&~_T_1805)
            begin $display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_379&~_T_1805)
            begin $display("fatal");
            end 
         if (_GEN_387&~_T_1485)
            begin $display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_387&~_T_1485)
            begin $display("fatal");
            end 
         if (_GEN_387&~_T_1488)
            begin $display("Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_387&~_T_1488)
            begin $display("fatal");
            end 
         if (_GEN_387&~_T_1495)
            begin $display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_387&~_T_1495)
            begin $display("fatal");
            end 
         if (_GEN_387&~_T_1805)
            begin $display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_387&~_T_1805)
            begin $display("fatal");
            end 
         if (_GEN_395&~_T_1485)
            begin $display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_395&~_T_1485)
            begin $display("fatal");
            end 
         if (_GEN_395&~_T_1488)
            begin $display("Assertion failed: 'C' channel HintAck carries invalid source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_395&~_T_1488)
            begin $display("fatal");
            end 
         if (_GEN_395&~_T_1495)
            begin $display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_395&~_T_1495)
            begin $display("fatal");
            end 
         if (_GEN_395&~_T_1805)
            begin $display("Assertion failed: 'C' channel HintAck carries invalid param (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_GEN_395&~_T_1805)
            begin $display("fatal");
            end 
         if (_T_1847&~_T_1850)
            begin $display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1847&~_T_1850)
            begin $display("fatal");
            end 
         if (_T_1847&~_T_1854)
            begin $display("Assertion failed: 'A' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1847&~_T_1854)
            begin $display("fatal");
            end 
         if (_T_1847&~_T_1858)
            begin $display("Assertion failed: 'A' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1847&~_T_1858)
            begin $display("fatal");
            end 
         if (_T_1847&~_T_1862)
            begin $display("Assertion failed: 'A' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1847&~_T_1862)
            begin $display("fatal");
            end 
         if (_T_1847&~_T_1866)
            begin $display("Assertion failed: 'A' channel address changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1847&~_T_1866)
            begin $display("fatal");
            end 
         if (_T_1871&~_T_1874)
            begin $display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1871&~_T_1874)
            begin $display("fatal");
            end 
         if (_T_1871&~_T_1878)
            begin $display("Assertion failed: 'D' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1871&~_T_1878)
            begin $display("fatal");
            end 
         if (_T_1871&~_T_1882)
            begin $display("Assertion failed: 'D' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1871&~_T_1882)
            begin $display("fatal");
            end 
         if (_T_1871&~_T_1886)
            begin $display("Assertion failed: 'D' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1871&~_T_1886)
            begin $display("fatal");
            end 
         if (_T_1871&~_T_1890)
            begin $display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1871&~_T_1890)
            begin $display("fatal");
            end 
         if (_T_1871&~_T_1894)
            begin $display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1871&~_T_1894)
            begin $display("fatal");
            end 
         if (_T_1899&~_T_1902)
            begin $display("Assertion failed: 'B' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1899&~_T_1902)
            begin $display("fatal");
            end 
         if (_T_1899&~_T_1906)
            begin $display("Assertion failed: 'B' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1899&~_T_1906)
            begin $display("fatal");
            end 
         if (_T_1899&~_T_1910)
            begin $display("Assertion failed: 'B' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1899&~_T_1910)
            begin $display("fatal");
            end 
         if (_T_1899&~_T_1914)
            begin $display("Assertion failed: 'B' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1899&~_T_1914)
            begin $display("fatal");
            end 
         if (_T_1899&~_T_1918)
            begin $display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1899&~_T_1918)
            begin $display("fatal");
            end 
         if (_T_1923&~_T_1926)
            begin $display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1923&~_T_1926)
            begin $display("fatal");
            end 
         if (_T_1923&~_T_1930)
            begin $display("Assertion failed: 'C' channel param changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1923&~_T_1930)
            begin $display("fatal");
            end 
         if (_T_1923&~_T_1934)
            begin $display("Assertion failed: 'C' channel size changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1923&~_T_1934)
            begin $display("fatal");
            end 
         if (_T_1923&~_T_1938)
            begin $display("Assertion failed: 'C' channel source changed within multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1923&~_T_1938)
            begin $display("fatal");
            end 
         if (_T_1923&~_T_1942)
            begin $display("Assertion failed: 'C' channel address changed with multibeat operation (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1923&~_T_1942)
            begin $display("fatal");
            end 
         if (_T_1949&~_T_1955)
            begin $display("Assertion failed: 'A' channel re-used a source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_1949&~_T_1955)
            begin $display("fatal");
            end 
         if (_T_1960&~_T_1974)
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1960&~_T_1974)
            begin $display("fatal");
            end 
         if (_GEN_403&~_T_1980)
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_403&~_T_1980)
            begin $display("fatal");
            end 
         if (_GEN_403&~_T_1984)
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_403&~_T_1984)
            begin $display("fatal");
            end 
         if (_GEN_408&~_T_1992)
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_408&~_T_1992)
            begin $display("fatal");
            end 
         if (_GEN_408&~_T_1996)
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_408&~_T_1996)
            begin $display("fatal");
            end 
         if (_T_2004&~_T_2008)
            begin $display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_2004&~_T_2008)
            begin $display("fatal");
            end 
         if (~_T_2015)
            begin $display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (~_T_2015)
            begin $display("fatal");
            end 
         if (~_T_2024)
            begin $display("Assertion failed: TileLink timeout expired (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~_T_2024)
            begin $display("fatal");
            end 
         if (_T_2039&~_T_2044)
            begin $display("Assertion failed: 'C' channel re-used a source ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_2039&~_T_2044)
            begin $display("fatal");
            end 
         if (_T_2048&~_T_2060)
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_2048&~_T_2060)
            begin $display("fatal");
            end 
         if (_GEN_415&~_T_2064)
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_415&~_T_2064)
            begin $display("fatal");
            end 
         if (_GEN_418&~_T_2068)
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_418&~_T_2068)
            begin $display("fatal");
            end 
         if (_T_2075&~_T_2079)
            begin $display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_2075&~_T_2079)
            begin $display("fatal");
            end 
         if (_T_2081&~_T_2084)
            begin $display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_2081&~_T_2084)
            begin $display("fatal");
            end 
         if (~_T_2093)
            begin $display("Assertion failed: TileLink timeout expired (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~_T_2093)
            begin $display("fatal");
            end 
         if (_T_2104&~_T_2109)
            begin $display("Assertion failed: 'D' channel re-used a sink ID (connected at HellaCache.scala:267:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_2104&~_T_2109)
            begin $display("fatal");
            end 
         if (_T_2111&~_T_2118)
            begin $display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at HellaCache.scala:267:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_2111&~_T_2118)
            begin $display("fatal");
            end 
         if (metaReset)
            begin 
              TLMonitor_23_metaAssert <=1'h0;
            end 
          else 
            begin 
              TLMonitor_23_metaAssert <=TLMonitor_23_metaAssert|TLMonitor_23_or0;
            end 
       end
  
endmodule
 
module TLMonitor_24 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [31:0] io_in_a_bits_address,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [31:0] plusarg_reader_out ;  
   wire [31:0] plusarg_reader_1_out ;  
   wire [31:0] _is_aligned_T ;  
   wire is_aligned ;  
   wire [32:0] _T_7 ;  
   wire [32:0] _T_26 ;  
   wire _T_27 ;  
   wire [31:0] _T_28 ;  
   wire [32:0] _T_29 ;  
   wire [32:0] _T_31 ;  
   wire _T_32 ;  
   wire [31:0] _T_33 ;  
   wire [32:0] _T_34 ;  
   wire [32:0] _T_36 ;  
   wire _T_37 ;  
   wire [31:0] _T_38 ;  
   wire [32:0] _T_39 ;  
   wire [32:0] _T_41 ;  
   wire _T_42 ;  
   wire [31:0] _T_43 ;  
   wire [32:0] _T_44 ;  
   wire [32:0] _T_46 ;  
   wire _T_47 ;  
   wire [31:0] _T_48 ;  
   wire [32:0] _T_49 ;  
   wire [32:0] _T_51 ;  
   wire _T_52 ;  
   wire [31:0] _T_63 ;  
   wire [32:0] _T_64 ;  
   wire [32:0] _T_66 ;  
   wire _T_67 ;  
   wire _T_134 ;  
   wire _T_341 ;  
   wire _T_342 ;  
   wire _T_343 ;  
   wire _T_344 ;  
   wire _T_345 ;  
   wire _T_348 ;  
   wire _T_350 ;  
   wire _T_766 ;  
   wire _T_768 ;  
   wire _T_770 ;  
   wire _T_774 ;  
   wire _T_776 ;  
   wire _T_778 ;  
   wire _T_780 ;  
   wire _T_784 ;  
   wire _T_788 ;  
   wire _T_790 ;  
   wire _T_801 ;  
   wire _T_803 ;  
   wire _T_805 ;  
   wire _T_807 ;  
   wire _T_818 ;  
   wire _T_838 ;  
   wire _T_840 ;  
   wire _T_847 ;  
   wire _T_864 ;  
   wire _T_882 ;  
   wire a_first_done ;  
   reg [8:0] a_first_counter ;  
   reg [31:0] _RAND_0 ;  
   wire [8:0] a_first_counter1 ;  
   wire a_first ;  
   reg [31:0] address ;  
   reg [31:0] _RAND_1 ;  
   wire _T_912 ;  
   wire _T_929 ;  
   wire _T_931 ;  
   wire _T_934 ;  
   wire [26:0] _d_first_beats1_decode_T_1 ;  
   wire [8:0] d_first_beats1_decode ;  
   wire d_first_beats1_opdata ;  
   reg [8:0] d_first_counter ;  
   reg [31:0] _RAND_2 ;  
   wire [8:0] d_first_counter1 ;  
   wire d_first ;  
   reg [2:0] opcode_1 ;  
   reg [31:0] _RAND_3 ;  
   reg [1:0] param_1 ;  
   reg [31:0] _RAND_4 ;  
   reg [3:0] size_1 ;  
   reg [31:0] _RAND_5 ;  
   reg [1:0] sink ;  
   reg [31:0] _RAND_6 ;  
   reg denied ;  
   reg [31:0] _RAND_7 ;  
   wire _T_936 ;  
   wire _T_937 ;  
   wire _T_939 ;  
   wire _T_941 ;  
   wire _T_943 ;  
   wire _T_945 ;  
   wire _T_947 ;  
   wire _T_953 ;  
   wire _T_955 ;  
   wire _T_957 ;  
   wire _T_959 ;  
   wire _T_962 ;  
   reg inflight ;  
   reg [31:0] _RAND_8 ;  
   reg [3:0] inflight_opcodes ;  
   reg [31:0] _RAND_9 ;  
   reg [7:0] inflight_sizes ;  
   reg [31:0] _RAND_10 ;  
   reg [8:0] a_first_counter_1 ;  
   reg [31:0] _RAND_11 ;  
   wire [8:0] a_first_counter1_1 ;  
   wire a_first_1 ;  
   reg [8:0] d_first_counter_1 ;  
   reg [31:0] _RAND_12 ;  
   wire [8:0] d_first_counter1_1 ;  
   wire d_first_1 ;  
   wire [15:0] _a_opcode_lookup_T_5 ;  
   wire [15:0] _GEN_71 ;  
   wire [15:0] _a_opcode_lookup_T_6 ;  
   wire [15:0] _a_opcode_lookup_T_7 ;  
   wire [15:0] _a_size_lookup_T_5 ;  
   wire [15:0] _GEN_73 ;  
   wire [15:0] _a_size_lookup_T_6 ;  
   wire [15:0] _a_size_lookup_T_7 ;  
   wire _T_963 ;  
   wire [1:0] _GEN_15 ;  
   wire _T_966 ;  
   wire [3:0] a_opcodes_set_interm ;  
   wire [18:0] _a_opcodes_set_T_1 ;  
   wire [4:0] a_sizes_set_interm ;  
   wire [19:0] _a_sizes_set_T_1 ;  
   wire _T_972 ;  
   wire [1:0] _GEN_16 ;  
   wire [18:0] _GEN_19 ;  
   wire [19:0] _GEN_20 ;  
   wire _T_974 ;  
   wire _T_977 ;  
   wire [1:0] _GEN_21 ;  
   wire [30:0] _d_opcodes_clr_T_5 ;  
   wire [30:0] _d_sizes_clr_T_5 ;  
   wire [30:0] _GEN_23 ;  
   wire [30:0] _GEN_24 ;  
   wire _T_989 ;  
   wire _T_991 ;  
   wire _T_995 ;  
   wire _T_997 ;  
   wire _T_999 ;  
   wire _T_1001 ;  
   wire [3:0] a_opcode_lookup ;  
   wire [2:0] _GEN_43 ;  
   wire [2:0] _GEN_44 ;  
   wire [2:0] _GEN_45 ;  
   wire [2:0] _GEN_46 ;  
   wire [2:0] _GEN_47 ;  
   wire [2:0] _GEN_48 ;  
   wire _T_1004 ;  
   wire [2:0] _GEN_55 ;  
   wire [2:0] _GEN_56 ;  
   wire _T_1006 ;  
   wire _T_1007 ;  
   wire _T_1009 ;  
   wire [7:0] a_size_lookup ;  
   wire [7:0] _GEN_75 ;  
   wire _T_1011 ;  
   wire _T_1013 ;  
   wire _T_1016 ;  
   wire _T_1017 ;  
   wire _T_1021 ;  
   wire _T_1025 ;  
   wire a_set_wo_ready ;  
   wire d_clr_wo_ready ;  
   wire _T_1027 ;  
   wire _T_1028 ;  
   wire _T_1030 ;  
   wire _T_1032 ;  
   wire a_set ;  
   wire _inflight_T ;  
   wire _inflight_T_2 ;  
   wire [3:0] a_opcodes_set ;  
   wire [3:0] _inflight_opcodes_T ;  
   wire [3:0] d_opcodes_clr ;  
   wire [3:0] _inflight_opcodes_T_2 ;  
   wire [7:0] a_sizes_set ;  
   wire [7:0] _inflight_sizes_T ;  
   wire [7:0] d_sizes_clr ;  
   wire [7:0] _inflight_sizes_T_2 ;  
   reg [31:0] watchdog ;  
   reg [31:0] _RAND_13 ;  
   wire _T_1034 ;  
   wire _T_1036 ;  
   wire _T_1037 ;  
   wire _T_1038 ;  
   wire _T_1039 ;  
   wire _T_1041 ;  
   wire [31:0] _watchdog_T_1 ;  
   wire _T_1045 ;  
   reg inflight_1 ;  
   reg [31:0] _RAND_14 ;  
   reg [7:0] inflight_sizes_1 ;  
   reg [31:0] _RAND_15 ;  
   reg [8:0] d_first_counter_2 ;  
   reg [31:0] _RAND_16 ;  
   wire [8:0] d_first_counter1_2 ;  
   wire d_first_2 ;  
   wire [15:0] _GEN_78 ;  
   wire [15:0] _c_size_lookup_T_6 ;  
   wire [15:0] _c_size_lookup_T_7 ;  
   wire _T_1063 ;  
   wire _T_1065 ;  
   wire [1:0] _GEN_66 ;  
   wire [30:0] _GEN_69 ;  
   wire _T_1077 ;  
   wire [7:0] c_size_lookup ;  
   wire _T_1083 ;  
   wire _T_1085 ;  
   wire _T_1098 ;  
   wire d_clr_wo_ready_1 ;  
   wire _T_1101 ;  
   wire _inflight_T_5 ;  
   wire [7:0] d_sizes_clr_1 ;  
   wire [7:0] _inflight_sizes_T_5 ;  
   reg [31:0] watchdog_1 ;  
   reg [31:0] _RAND_17 ;  
   wire _T_1103 ;  
   wire _T_1105 ;  
   wire _T_1106 ;  
   wire _T_1107 ;  
   wire _T_1108 ;  
   wire _T_1110 ;  
   wire [31:0] _watchdog_T_3 ;  
   wire _GEN_81 ;  
   wire _GEN_89 ;  
   wire _GEN_97 ;  
   wire _GEN_105 ;  
   wire _GEN_109 ;  
   wire _GEN_113 ;  
   wire _GEN_117 ;  
   wire _GEN_122 ;  
   wire [29:0] TLMonitor_24_covSum ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire stopEn2 ;  
   wire stopEn3 ;  
   wire stopEn4 ;  
   wire stopEn5 ;  
   wire stopEn6 ;  
   wire stopEn7 ;  
   wire stopEn8 ;  
   wire stopEn9 ;  
   wire stopEn10 ;  
   wire stopEn11 ;  
   wire stopEn12 ;  
   wire stopEn13 ;  
   wire stopEn14 ;  
   wire stopEn15 ;  
   wire stopEn16 ;  
   wire stopEn17 ;  
   wire stopEn18 ;  
   wire stopEn19 ;  
   wire stopEn20 ;  
   wire stopEn21 ;  
   wire stopEn22 ;  
   wire stopEn23 ;  
   wire stopEn24 ;  
   wire stopEn25 ;  
   wire stopEn26 ;  
   wire stopEn27 ;  
   wire stopEn28 ;  
   wire stopEn29 ;  
   wire stopEn30 ;  
   wire stopEn31 ;  
   wire stopEn32 ;  
   wire stopEn33 ;  
   wire stopEn34 ;  
   wire stopEn35 ;  
   wire stopEn36 ;  
   wire stopEn37 ;  
   wire stopEn38 ;  
   wire stopEn39 ;  
   wire plusarg_reader_metaAssert_wire ;  
   wire plusarg_reader_1_metaAssert_wire ;  
   wire TLMonitor_24_or15 ;  
   wire TLMonitor_24_or34 ;  
   wire TLMonitor_24_or16 ;  
   wire TLMonitor_24_or7 ;  
   wire TLMonitor_24_or17 ;  
   wire TLMonitor_24_or38 ;  
   wire TLMonitor_24_or18 ;  
   wire TLMonitor_24_or8 ;  
   wire TLMonitor_24_or3 ;  
   wire TLMonitor_24_or19 ;  
   wire TLMonitor_24_or42 ;  
   wire TLMonitor_24_or20 ;  
   wire TLMonitor_24_or9 ;  
   wire TLMonitor_24_or44 ;  
   wire TLMonitor_24_or21 ;  
   wire TLMonitor_24_or46 ;  
   wire TLMonitor_24_or22 ;  
   wire TLMonitor_24_or10 ;  
   wire TLMonitor_24_or4 ;  
   wire TLMonitor_24_or1 ;  
   wire TLMonitor_24_or23 ;  
   wire TLMonitor_24_or50 ;  
   wire TLMonitor_24_or24 ;  
   wire TLMonitor_24_or11 ;  
   wire TLMonitor_24_or25 ;  
   wire TLMonitor_24_or54 ;  
   wire TLMonitor_24_or26 ;  
   wire TLMonitor_24_or12 ;  
   wire TLMonitor_24_or5 ;  
   wire TLMonitor_24_or27 ;  
   wire TLMonitor_24_or58 ;  
   wire TLMonitor_24_or28 ;  
   wire TLMonitor_24_or13 ;  
   wire TLMonitor_24_or60 ;  
   wire TLMonitor_24_or29 ;  
   wire TLMonitor_24_or62 ;  
   wire TLMonitor_24_or30 ;  
   wire TLMonitor_24_or14 ;  
   wire TLMonitor_24_or6 ;  
   wire TLMonitor_24_or2 ;  
   wire TLMonitor_24_or0 ;  
   reg TLMonitor_24_metaAssert ;  
   reg [31:0] _RAND_18 ;  
  assign _is_aligned_T=io_in_a_bits_address&32'h3f; 
  assign is_aligned=_is_aligned_T==32'h0; 
  assign _T_7={1'b0,$signed(io_in_a_bits_address)}; 
  assign _T_26=$signed(_T_7)&-33'sh1000; 
  assign _T_27=$signed(_T_26)==33'sh0; 
  assign _T_28=io_in_a_bits_address^32'h3000; 
  assign _T_29={1'b0,$signed(_T_28)}; 
  assign _T_31=$signed(_T_29)&-33'sh1000; 
  assign _T_32=$signed(_T_31)==33'sh0; 
  assign _T_33=io_in_a_bits_address^32'h10000; 
  assign _T_34={1'b0,$signed(_T_33)}; 
  assign _T_36=$signed(_T_34)&-33'sh10000; 
  assign _T_37=$signed(_T_36)==33'sh0; 
  assign _T_38=io_in_a_bits_address^32'h2000000; 
  assign _T_39={1'b0,$signed(_T_38)}; 
  assign _T_41=$signed(_T_39)&-33'sh10000; 
  assign _T_42=$signed(_T_41)==33'sh0; 
  assign _T_43=io_in_a_bits_address^32'hc000000; 
  assign _T_44={1'b0,$signed(_T_43)}; 
  assign _T_46=$signed(_T_44)&-33'sh4000000; 
  assign _T_47=$signed(_T_46)==33'sh0; 
  assign _T_48=io_in_a_bits_address^32'h60000000; 
  assign _T_49={1'b0,$signed(_T_48)}; 
  assign _T_51=$signed(_T_49)&-33'sh20000000; 
  assign _T_52=$signed(_T_51)==33'sh0; 
  assign _T_63=io_in_a_bits_address^32'h80000000; 
  assign _T_64={1'b0,$signed(_T_63)}; 
  assign _T_66=$signed(_T_64)&-33'sh10000000; 
  assign _T_67=$signed(_T_66)==33'sh0; 
  assign _T_134=is_aligned|reset; 
  assign _T_341=_T_27|_T_37; 
  assign _T_342=_T_341|_T_42; 
  assign _T_343=_T_342|_T_47; 
  assign _T_344=_T_343|_T_52; 
  assign _T_345=_T_344|_T_67; 
  assign _T_348=_T_32|_T_345; 
  assign _T_350=_T_348|reset; 
  assign _T_766=io_in_d_bits_opcode<=3'h6; 
  assign _T_768=_T_766|reset; 
  assign _T_770=io_in_d_bits_opcode==3'h6; 
  assign _T_774=io_in_d_bits_size>=4'h3; 
  assign _T_776=_T_774|reset; 
  assign _T_778=io_in_d_bits_param==2'h0; 
  assign _T_780=_T_778|reset; 
  assign _T_784=~io_in_d_bits_corrupt|reset; 
  assign _T_788=~io_in_d_bits_denied|reset; 
  assign _T_790=io_in_d_bits_opcode==3'h4; 
  assign _T_801=io_in_d_bits_param<=2'h2; 
  assign _T_803=_T_801|reset; 
  assign _T_805=io_in_d_bits_param!=2'h2; 
  assign _T_807=_T_805|reset; 
  assign _T_818=io_in_d_bits_opcode==3'h5; 
  assign _T_838=~io_in_d_bits_denied|io_in_d_bits_corrupt; 
  assign _T_840=_T_838|reset; 
  assign _T_847=io_in_d_bits_opcode==3'h0; 
  assign _T_864=io_in_d_bits_opcode==3'h1; 
  assign _T_882=io_in_d_bits_opcode==3'h2; 
  assign a_first_done=io_in_a_ready&io_in_a_valid; 
  assign a_first_counter1=a_first_counter-9'h1; 
  assign a_first=a_first_counter==9'h0; 
  assign _T_912=io_in_a_valid&~a_first; 
  assign _T_929=io_in_a_bits_address==address; 
  assign _T_931=_T_929|reset; 
  assign _T_934=a_first_done&a_first; 
  assign _d_first_beats1_decode_T_1=27'hfff<<io_in_d_bits_size; 
  assign d_first_beats1_decode=~_d_first_beats1_decode_T_1[11:3]; 
  assign d_first_beats1_opdata=io_in_d_bits_opcode[0]; 
  assign d_first_counter1=d_first_counter-9'h1; 
  assign d_first=d_first_counter==9'h0; 
  assign _T_936=io_in_d_valid&~d_first; 
  assign _T_937=io_in_d_bits_opcode==opcode_1; 
  assign _T_939=_T_937|reset; 
  assign _T_941=io_in_d_bits_param==param_1; 
  assign _T_943=_T_941|reset; 
  assign _T_945=io_in_d_bits_size==size_1; 
  assign _T_947=_T_945|reset; 
  assign _T_953=io_in_d_bits_sink==sink; 
  assign _T_955=_T_953|reset; 
  assign _T_957=io_in_d_bits_denied==denied; 
  assign _T_959=_T_957|reset; 
  assign _T_962=io_in_d_valid&d_first; 
  assign a_first_counter1_1=a_first_counter_1-9'h1; 
  assign a_first_1=a_first_counter_1==9'h0; 
  assign d_first_counter1_1=d_first_counter_1-9'h1; 
  assign d_first_1=d_first_counter_1==9'h0; 
  assign _a_opcode_lookup_T_5=16'h10-16'h1; 
  assign _GEN_71={12'b0,inflight_opcodes}; 
  assign _a_opcode_lookup_T_6=_GEN_71&_a_opcode_lookup_T_5; 
  assign _a_opcode_lookup_T_7={1'b0,_a_opcode_lookup_T_6[15:1]}; 
  assign _a_size_lookup_T_5=16'h100-16'h1; 
  assign _GEN_73={8'b0,inflight_sizes}; 
  assign _a_size_lookup_T_6=_GEN_73&_a_size_lookup_T_5; 
  assign _a_size_lookup_T_7={1'b0,_a_size_lookup_T_6[15:1]}; 
  assign _T_963=io_in_a_valid&a_first_1; 
  assign _GEN_15=_T_963 ? 2'h1:2'h0; 
  assign _T_966=a_first_done&a_first_1; 
  assign a_opcodes_set_interm=_T_966 ? 4'h9:4'h0; 
  assign _a_opcodes_set_T_1={15'b0,a_opcodes_set_interm}; 
  assign a_sizes_set_interm=_T_966 ? 5'hd:5'h0; 
  assign _a_sizes_set_T_1={15'b0,a_sizes_set_interm}; 
  assign _T_972=~inflight|reset; 
  assign _GEN_16=_T_966 ? 2'h1:2'h0; 
  assign _GEN_19=_T_966 ? _a_opcodes_set_T_1:19'h0; 
  assign _GEN_20=_T_966 ? _a_sizes_set_T_1:20'h0; 
  assign _T_974=io_in_d_valid&d_first_1; 
  assign _T_977=_T_974&~_T_770; 
  assign _GEN_21=_T_977 ? 2'h1:2'h0; 
  assign _d_opcodes_clr_T_5={15'b0,_a_opcode_lookup_T_5}; 
  assign _d_sizes_clr_T_5={15'b0,_a_size_lookup_T_5}; 
  assign _GEN_23=_T_977 ? _d_opcodes_clr_T_5:31'h0; 
  assign _GEN_24=_T_977 ? _d_sizes_clr_T_5:31'h0; 
  assign _T_989=inflight|_T_963; 
  assign _T_991=_T_989|reset; 
  assign _T_995=_T_864|_T_864; 
  assign _T_997=_T_995|reset; 
  assign _T_999=4'h6==io_in_d_bits_size; 
  assign _T_1001=_T_999|reset; 
  assign a_opcode_lookup=_a_opcode_lookup_T_7[3:0]; 
  assign _GEN_43=3'h2==a_opcode_lookup[2:0] ? 3'h1:3'h0; 
  assign _GEN_44=3'h3==a_opcode_lookup[2:0] ? 3'h1:_GEN_43; 
  assign _GEN_45=3'h4==a_opcode_lookup[2:0] ? 3'h1:_GEN_44; 
  assign _GEN_46=3'h5==a_opcode_lookup[2:0] ? 3'h2:_GEN_45; 
  assign _GEN_47=3'h6==a_opcode_lookup[2:0] ? 3'h4:_GEN_46; 
  assign _GEN_48=3'h7==a_opcode_lookup[2:0] ? 3'h4:_GEN_47; 
  assign _T_1004=io_in_d_bits_opcode==_GEN_48; 
  assign _GEN_55=3'h6==a_opcode_lookup[2:0] ? 3'h5:_GEN_46; 
  assign _GEN_56=3'h7==a_opcode_lookup[2:0] ? 3'h4:_GEN_55; 
  assign _T_1006=io_in_d_bits_opcode==_GEN_56; 
  assign _T_1007=_T_1004|_T_1006; 
  assign _T_1009=_T_1007|reset; 
  assign a_size_lookup=_a_size_lookup_T_7[7:0]; 
  assign _GEN_75={4'b0,io_in_d_bits_size}; 
  assign _T_1011=_GEN_75==a_size_lookup; 
  assign _T_1013=_T_1011|reset; 
  assign _T_1016=_T_974&a_first_1; 
  assign _T_1017=_T_1016&io_in_a_valid; 
  assign _T_1021=_T_1017&~_T_770; 
  assign _T_1025=io_in_a_ready|reset; 
  assign a_set_wo_ready=_GEN_15[0]; 
  assign d_clr_wo_ready=_GEN_21[0]; 
  assign _T_1027=a_set_wo_ready!=d_clr_wo_ready; 
  assign _T_1028=|a_set_wo_ready; 
  assign _T_1030=_T_1027|~_T_1028; 
  assign _T_1032=_T_1030|reset; 
  assign a_set=_GEN_16[0]; 
  assign _inflight_T=inflight|a_set; 
  assign _inflight_T_2=_inflight_T&~d_clr_wo_ready; 
  assign a_opcodes_set=_GEN_19[3:0]; 
  assign _inflight_opcodes_T=inflight_opcodes|a_opcodes_set; 
  assign d_opcodes_clr=_GEN_23[3:0]; 
  assign _inflight_opcodes_T_2=_inflight_opcodes_T&~d_opcodes_clr; 
  assign a_sizes_set=_GEN_20[7:0]; 
  assign _inflight_sizes_T=inflight_sizes|a_sizes_set; 
  assign d_sizes_clr=_GEN_24[7:0]; 
  assign _inflight_sizes_T_2=_inflight_sizes_T&~d_sizes_clr; 
  assign _T_1034=|inflight; 
  assign _T_1036=plusarg_reader_out==32'h0; 
  assign _T_1037=~_T_1034|_T_1036; 
  assign _T_1038=watchdog<plusarg_reader_out; 
  assign _T_1039=_T_1037|_T_1038; 
  assign _T_1041=_T_1039|reset; 
  assign _watchdog_T_1=watchdog+32'h1; 
  assign _T_1045=a_first_done|io_in_d_valid; 
  assign d_first_counter1_2=d_first_counter_2-9'h1; 
  assign d_first_2=d_first_counter_2==9'h0; 
  assign _GEN_78={8'b0,inflight_sizes_1}; 
  assign _c_size_lookup_T_6=_GEN_78&_a_size_lookup_T_5; 
  assign _c_size_lookup_T_7={1'b0,_c_size_lookup_T_6[15:1]}; 
  assign _T_1063=io_in_d_valid&d_first_2; 
  assign _T_1065=_T_1063&_T_770; 
  assign _GEN_66=_T_1065 ? 2'h1:2'h0; 
  assign _GEN_69=_T_1065 ? _d_sizes_clr_T_5:31'h0; 
  assign _T_1077=inflight_1|reset; 
  assign c_size_lookup=_c_size_lookup_T_7[7:0]; 
  assign _T_1083=_GEN_75==c_size_lookup; 
  assign _T_1085=_T_1083|reset; 
  assign _T_1098=|1'h0; 
  assign d_clr_wo_ready_1=_GEN_66[0]; 
  assign _T_1101=d_clr_wo_ready_1|reset; 
  assign _inflight_T_5=inflight_1&~d_clr_wo_ready_1; 
  assign d_sizes_clr_1=_GEN_69[7:0]; 
  assign _inflight_sizes_T_5=inflight_sizes_1&~d_sizes_clr_1; 
  assign _T_1103=|inflight_1; 
  assign _T_1105=plusarg_reader_1_out==32'h0; 
  assign _T_1106=~_T_1103|_T_1105; 
  assign _T_1107=watchdog_1<plusarg_reader_1_out; 
  assign _T_1108=_T_1106|_T_1107; 
  assign _T_1110=_T_1108|reset; 
  assign _watchdog_T_3=watchdog_1+32'h1; 
  assign _GEN_81=io_in_d_valid&_T_770; 
  assign _GEN_89=io_in_d_valid&_T_790; 
  assign _GEN_97=io_in_d_valid&_T_818; 
  assign _GEN_105=io_in_d_valid&_T_847; 
  assign _GEN_109=io_in_d_valid&_T_864; 
  assign _GEN_113=io_in_d_valid&_T_882; 
  assign _GEN_117=_T_977&_T_963; 
  assign _GEN_122=_T_977&~_T_963; 
  assign TLMonitor_24_covSum=30'h0; 
  assign io_covSum=TLMonitor_24_covSum; 
  assign stopEn0=io_in_a_valid&~_T_350; 
  assign stopEn1=io_in_a_valid&~_T_134; 
  assign stopEn2=io_in_d_valid&~_T_768; 
  assign stopEn3=_GEN_81&~_T_776; 
  assign stopEn4=_GEN_81&~_T_780; 
  assign stopEn5=_GEN_81&~_T_784; 
  assign stopEn6=_GEN_81&~_T_788; 
  assign stopEn7=_GEN_89&~_T_776; 
  assign stopEn8=_GEN_89&~_T_803; 
  assign stopEn9=_GEN_89&~_T_807; 
  assign stopEn10=_GEN_89&~_T_784; 
  assign stopEn11=_GEN_97&~_T_776; 
  assign stopEn12=_GEN_97&~_T_803; 
  assign stopEn13=_GEN_97&~_T_807; 
  assign stopEn14=_GEN_97&~_T_840; 
  assign stopEn15=_GEN_105&~_T_780; 
  assign stopEn16=_GEN_105&~_T_784; 
  assign stopEn17=_GEN_109&~_T_780; 
  assign stopEn18=_GEN_109&~_T_840; 
  assign stopEn19=_GEN_113&~_T_780; 
  assign stopEn20=_GEN_113&~_T_784; 
  assign stopEn21=_T_912&~_T_931; 
  assign stopEn22=_T_936&~_T_939; 
  assign stopEn23=_T_936&~_T_943; 
  assign stopEn24=_T_936&~_T_947; 
  assign stopEn25=_T_936&~_T_955; 
  assign stopEn26=_T_936&~_T_959; 
  assign stopEn27=_T_966&~_T_972; 
  assign stopEn28=_T_977&~_T_991; 
  assign stopEn29=_GEN_117&~_T_997; 
  assign stopEn30=_GEN_117&~_T_1001; 
  assign stopEn31=_GEN_122&~_T_1009; 
  assign stopEn32=_GEN_122&~_T_1013; 
  assign stopEn33=_T_1021&~_T_1025; 
  assign stopEn34=~_T_1032; 
  assign stopEn35=~_T_1041; 
  assign stopEn36=_T_1065&~_T_1077; 
  assign stopEn37=_T_1065&~_T_1085; 
  assign stopEn38=_T_1098&~_T_1101; 
  assign stopEn39=~_T_1110; 
  assign TLMonitor_24_or15=stopEn0|stopEn1; 
  assign TLMonitor_24_or34=stopEn3|stopEn4; 
  assign TLMonitor_24_or16=stopEn2|TLMonitor_24_or34; 
  assign TLMonitor_24_or7=TLMonitor_24_or15|TLMonitor_24_or16; 
  assign TLMonitor_24_or17=stopEn5|stopEn6; 
  assign TLMonitor_24_or38=stopEn8|stopEn9; 
  assign TLMonitor_24_or18=stopEn7|TLMonitor_24_or38; 
  assign TLMonitor_24_or8=TLMonitor_24_or17|TLMonitor_24_or18; 
  assign TLMonitor_24_or3=TLMonitor_24_or7|TLMonitor_24_or8; 
  assign TLMonitor_24_or19=stopEn10|stopEn11; 
  assign TLMonitor_24_or42=stopEn13|stopEn14; 
  assign TLMonitor_24_or20=stopEn12|TLMonitor_24_or42; 
  assign TLMonitor_24_or9=TLMonitor_24_or19|TLMonitor_24_or20; 
  assign TLMonitor_24_or44=stopEn16|stopEn17; 
  assign TLMonitor_24_or21=stopEn15|TLMonitor_24_or44; 
  assign TLMonitor_24_or46=stopEn19|stopEn20; 
  assign TLMonitor_24_or22=stopEn18|TLMonitor_24_or46; 
  assign TLMonitor_24_or10=TLMonitor_24_or21|TLMonitor_24_or22; 
  assign TLMonitor_24_or4=TLMonitor_24_or9|TLMonitor_24_or10; 
  assign TLMonitor_24_or1=TLMonitor_24_or3|TLMonitor_24_or4; 
  assign TLMonitor_24_or23=stopEn21|stopEn22; 
  assign TLMonitor_24_or50=stopEn24|stopEn25; 
  assign TLMonitor_24_or24=stopEn23|TLMonitor_24_or50; 
  assign TLMonitor_24_or11=TLMonitor_24_or23|TLMonitor_24_or24; 
  assign TLMonitor_24_or25=stopEn26|stopEn27; 
  assign TLMonitor_24_or54=stopEn29|stopEn30; 
  assign TLMonitor_24_or26=stopEn28|TLMonitor_24_or54; 
  assign TLMonitor_24_or12=TLMonitor_24_or25|TLMonitor_24_or26; 
  assign TLMonitor_24_or5=TLMonitor_24_or11|TLMonitor_24_or12; 
  assign TLMonitor_24_or27=stopEn31|stopEn32; 
  assign TLMonitor_24_or58=stopEn34|stopEn35; 
  assign TLMonitor_24_or28=stopEn33|TLMonitor_24_or58; 
  assign TLMonitor_24_or13=TLMonitor_24_or27|TLMonitor_24_or28; 
  assign TLMonitor_24_or60=stopEn37|stopEn38; 
  assign TLMonitor_24_or29=stopEn36|TLMonitor_24_or60; 
  assign TLMonitor_24_or62=plusarg_reader_metaAssert_wire|plusarg_reader_1_metaAssert_wire; 
  assign TLMonitor_24_or30=stopEn39|TLMonitor_24_or62; 
  assign TLMonitor_24_or14=TLMonitor_24_or29|TLMonitor_24_or30; 
  assign TLMonitor_24_or6=TLMonitor_24_or13|TLMonitor_24_or14; 
  assign TLMonitor_24_or2=TLMonitor_24_or5|TLMonitor_24_or6; 
  assign TLMonitor_24_or0=TLMonitor_24_or1|TLMonitor_24_or2; 
  assign metaAssert=TLMonitor_24_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              a_first_counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 a_first_counter <=9'h0;
               end 
             else 
               if (a_first_done)
                  begin 
                    if (a_first)
                       begin 
                         a_first_counter <=9'h0;
                       end 
                     else 
                       begin 
                         a_first_counter <=a_first_counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              address <=32'h0;
            end 
          else 
            if (_T_934)
               begin 
                 address <=io_in_a_bits_address;
               end 
         if (metaReset)
            begin 
              d_first_counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 d_first_counter <=9'h0;
               end 
             else 
               if (io_in_d_valid)
                  begin 
                    if (d_first)
                       begin 
                         if (d_first_beats1_opdata)
                            begin 
                              d_first_counter <=d_first_beats1_decode;
                            end 
                          else 
                            begin 
                              d_first_counter <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         d_first_counter <=d_first_counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              opcode_1 <=3'h0;
            end 
          else 
            if (_T_962)
               begin 
                 opcode_1 <=io_in_d_bits_opcode;
               end 
         if (metaReset)
            begin 
              param_1 <=2'h0;
            end 
          else 
            if (_T_962)
               begin 
                 param_1 <=io_in_d_bits_param;
               end 
         if (metaReset)
            begin 
              size_1 <=4'h0;
            end 
          else 
            if (_T_962)
               begin 
                 size_1 <=io_in_d_bits_size;
               end 
         if (metaReset)
            begin 
              sink <=2'h0;
            end 
          else 
            if (_T_962)
               begin 
                 sink <=io_in_d_bits_sink;
               end 
         if (metaReset)
            begin 
              denied <=1'h0;
            end 
          else 
            if (_T_962)
               begin 
                 denied <=io_in_d_bits_denied;
               end 
         if (metaReset)
            begin 
              inflight <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight <=1'h0;
               end 
             else 
               begin 
                 inflight <=_inflight_T_2;
               end 
         if (metaReset)
            begin 
              inflight_opcodes <=4'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_opcodes <=4'h0;
               end 
             else 
               begin 
                 inflight_opcodes <=_inflight_opcodes_T_2;
               end 
         if (metaReset)
            begin 
              inflight_sizes <=8'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_sizes <=8'h0;
               end 
             else 
               begin 
                 inflight_sizes <=_inflight_sizes_T_2;
               end 
         if (metaReset)
            begin 
              a_first_counter_1 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 a_first_counter_1 <=9'h0;
               end 
             else 
               if (a_first_done)
                  begin 
                    if (a_first_1)
                       begin 
                         a_first_counter_1 <=9'h0;
                       end 
                     else 
                       begin 
                         a_first_counter_1 <=a_first_counter1_1;
                       end 
                  end 
         if (metaReset)
            begin 
              d_first_counter_1 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 d_first_counter_1 <=9'h0;
               end 
             else 
               if (io_in_d_valid)
                  begin 
                    if (d_first_1)
                       begin 
                         if (d_first_beats1_opdata)
                            begin 
                              d_first_counter_1 <=d_first_beats1_decode;
                            end 
                          else 
                            begin 
                              d_first_counter_1 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         d_first_counter_1 <=d_first_counter1_1;
                       end 
                  end 
         if (metaReset)
            begin 
              watchdog <=32'h0;
            end 
          else 
            if (reset)
               begin 
                 watchdog <=32'h0;
               end 
             else 
               if (_T_1045)
                  begin 
                    watchdog <=32'h0;
                  end 
                else 
                  begin 
                    watchdog <=_watchdog_T_1;
                  end 
         if (metaReset)
            begin 
              inflight_1 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_1 <=1'h0;
               end 
             else 
               begin 
                 inflight_1 <=_inflight_T_5;
               end 
         if (metaReset)
            begin 
              inflight_sizes_1 <=8'h0;
            end 
          else 
            if (reset)
               begin 
                 inflight_sizes_1 <=8'h0;
               end 
             else 
               begin 
                 inflight_sizes_1 <=_inflight_sizes_T_5;
               end 
         if (metaReset)
            begin 
              d_first_counter_2 <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 d_first_counter_2 <=9'h0;
               end 
             else 
               if (io_in_d_valid)
                  begin 
                    if (d_first_2)
                       begin 
                         if (d_first_beats1_opdata)
                            begin 
                              d_first_counter_2 <=d_first_beats1_decode;
                            end 
                          else 
                            begin 
                              d_first_counter_2 <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         d_first_counter_2 <=d_first_counter1_2;
                       end 
                  end 
         if (metaReset)
            begin 
              watchdog_1 <=32'h0;
            end 
          else 
            if (reset)
               begin 
                 watchdog_1 <=32'h0;
               end 
             else 
               if (io_in_d_valid)
                  begin 
                    watchdog_1 <=32'h0;
                  end 
                else 
                  begin 
                    watchdog_1 <=_watchdog_T_3;
                  end 
         if (io_in_a_valid&~_T_350)
            begin $display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (io_in_a_valid&~_T_350)
            begin $display("fatal");
            end 
         if (io_in_a_valid&~_T_134)
            begin $display("Assertion failed: 'A' channel Get address not aligned to size (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (io_in_a_valid&~_T_134)
            begin $display("fatal");
            end 
         if (io_in_d_valid&~_T_768)
            begin $display("Assertion failed: 'D' channel has invalid opcode (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (io_in_d_valid&~_T_768)
            begin $display("fatal");
            end 
         if (_GEN_81&~_T_776)
            begin $display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_81&~_T_776)
            begin $display("fatal");
            end 
         if (_GEN_81&~_T_780)
            begin $display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_81&~_T_780)
            begin $display("fatal");
            end 
         if (_GEN_81&~_T_784)
            begin $display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_81&~_T_784)
            begin $display("fatal");
            end 
         if (_GEN_81&~_T_788)
            begin $display("Assertion failed: 'D' channel ReleaseAck is denied (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_81&~_T_788)
            begin $display("fatal");
            end 
         if (_GEN_89&~_T_776)
            begin $display("Assertion failed: 'D' channel Grant smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_89&~_T_776)
            begin $display("fatal");
            end 
         if (_GEN_89&~_T_803)
            begin $display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_89&~_T_803)
            begin $display("fatal");
            end 
         if (_GEN_89&~_T_807)
            begin $display("Assertion failed: 'D' channel Grant carries toN param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_89&~_T_807)
            begin $display("fatal");
            end 
         if (_GEN_89&~_T_784)
            begin $display("Assertion failed: 'D' channel Grant is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_89&~_T_784)
            begin $display("fatal");
            end 
         if (_GEN_97&~_T_776)
            begin $display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_97&~_T_776)
            begin $display("fatal");
            end 
         if (_GEN_97&~_T_803)
            begin $display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_97&~_T_803)
            begin $display("fatal");
            end 
         if (_GEN_97&~_T_807)
            begin $display("Assertion failed: 'D' channel GrantData carries toN param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_97&~_T_807)
            begin $display("fatal");
            end 
         if (_GEN_97&~_T_840)
            begin $display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_97&~_T_840)
            begin $display("fatal");
            end 
         if (_GEN_105&~_T_780)
            begin $display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_105&~_T_780)
            begin $display("fatal");
            end 
         if (_GEN_105&~_T_784)
            begin $display("Assertion failed: 'D' channel AccessAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_105&~_T_784)
            begin $display("fatal");
            end 
         if (_GEN_109&~_T_780)
            begin $display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_109&~_T_780)
            begin $display("fatal");
            end 
         if (_GEN_109&~_T_840)
            begin $display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_109&~_T_840)
            begin $display("fatal");
            end 
         if (_GEN_113&~_T_780)
            begin $display("Assertion failed: 'D' channel HintAck carries invalid param (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_113&~_T_780)
            begin $display("fatal");
            end 
         if (_GEN_113&~_T_784)
            begin $display("Assertion failed: 'D' channel HintAck is corrupt (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_113&~_T_784)
            begin $display("fatal");
            end 
         if (_T_912&~_T_931)
            begin $display("Assertion failed: 'A' channel address changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_912&~_T_931)
            begin $display("fatal");
            end 
         if (_T_936&~_T_939)
            begin $display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_936&~_T_939)
            begin $display("fatal");
            end 
         if (_T_936&~_T_943)
            begin $display("Assertion failed: 'D' channel param changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_936&~_T_943)
            begin $display("fatal");
            end 
         if (_T_936&~_T_947)
            begin $display("Assertion failed: 'D' channel size changed within multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_936&~_T_947)
            begin $display("fatal");
            end 
         if (_T_936&~_T_955)
            begin $display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_936&~_T_955)
            begin $display("fatal");
            end 
         if (_T_936&~_T_959)
            begin $display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_936&~_T_959)
            begin $display("fatal");
            end 
         if (_T_966&~_T_972)
            begin $display("Assertion failed: 'A' channel re-used a source ID (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (_T_966&~_T_972)
            begin $display("fatal");
            end 
         if (_T_977&~_T_991)
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_977&~_T_991)
            begin $display("fatal");
            end 
         if (_GEN_117&~_T_997)
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_117&~_T_997)
            begin $display("fatal");
            end 
         if (_GEN_117&~_T_1001)
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_117&~_T_1001)
            begin $display("fatal");
            end 
         if (_GEN_122&~_T_1009)
            begin $display("Assertion failed: 'D' channel contains improper opcode response (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_122&~_T_1009)
            begin $display("fatal");
            end 
         if (_GEN_122&~_T_1013)
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_GEN_122&~_T_1013)
            begin $display("fatal");
            end 
         if (_T_1021&~_T_1025)
            begin $display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1021&~_T_1025)
            begin $display("fatal");
            end 
         if (~_T_1032)
            begin $display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (~_T_1032)
            begin $display("fatal");
            end 
         if (~_T_1041)
            begin $display("Assertion failed: TileLink timeout expired (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~_T_1041)
            begin $display("fatal");
            end 
         if (_T_1065&~_T_1077)
            begin $display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1065&~_T_1077)
            begin $display("fatal");
            end 
         if (_T_1065&~_T_1085)
            begin $display("Assertion failed: 'D' channel contains improper response size (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1065&~_T_1085)
            begin $display("fatal");
            end 
         if (_T_1098&~_T_1101)
            begin $display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at Frontend.scala:351:21)\n    at Monitor.scala:49 assert(cond, message)\n");
            end 
         if (_T_1098&~_T_1101)
            begin $display("fatal");
            end 
         if (~_T_1110)
            begin $display("Assertion failed: TileLink timeout expired (connected at Frontend.scala:351:21)\n    at Monitor.scala:42 assert(cond, message)\n");
            end 
         if (~_T_1110)
            begin $display("fatal");
            end 
         if (metaReset)
            begin 
              TLMonitor_24_metaAssert <=1'h0;
            end 
          else 
            begin 
              TLMonitor_24_metaAssert <=TLMonitor_24_metaAssert|TLMonitor_24_or0;
            end 
       end
  
endmodule
 
module TLB (
  input clock,
  input reset,
  output io_req_ready,
  input io_req_valid,
  input [39:0] io_req_bits_vaddr,
  input io_req_bits_passthrough,
  input [1:0] io_req_bits_size,
  input [4:0] io_req_bits_cmd,
  output io_resp_miss,
  output [31:0] io_resp_paddr,
  output io_resp_pf_ld,
  output io_resp_pf_st,
  output io_resp_ae_ld,
  output io_resp_ae_st,
  output io_resp_ma_ld,
  output io_resp_ma_st,
  output io_resp_cacheable,
  input io_sfence_valid,
  input io_sfence_bits_rs1,
  input io_sfence_bits_rs2,
  input [38:0] io_sfence_bits_addr,
  input io_ptw_req_ready,
  output io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input io_ptw_resp_valid,
  input io_ptw_resp_bits_ae,
  input [53:0] io_ptw_resp_bits_pte_ppn,
  input io_ptw_resp_bits_pte_d,
  input io_ptw_resp_bits_pte_a,
  input io_ptw_resp_bits_pte_g,
  input io_ptw_resp_bits_pte_u,
  input io_ptw_resp_bits_pte_x,
  input io_ptw_resp_bits_pte_w,
  input io_ptw_resp_bits_pte_r,
  input io_ptw_resp_bits_pte_v,
  input [1:0] io_ptw_resp_bits_level,
  input io_ptw_resp_bits_homogeneous,
  input [3:0] io_ptw_ptbr_mode,
  input io_ptw_status_debug,
  input [1:0] io_ptw_status_dprv,
  input io_ptw_status_mxr,
  input io_ptw_status_sum,
  input io_ptw_pmp_0_cfg_l,
  input [1:0] io_ptw_pmp_0_cfg_a,
  input io_ptw_pmp_0_cfg_x,
  input io_ptw_pmp_0_cfg_w,
  input io_ptw_pmp_0_cfg_r,
  input [29:0] io_ptw_pmp_0_addr,
  input [31:0] io_ptw_pmp_0_mask,
  input io_ptw_pmp_1_cfg_l,
  input [1:0] io_ptw_pmp_1_cfg_a,
  input io_ptw_pmp_1_cfg_x,
  input io_ptw_pmp_1_cfg_w,
  input io_ptw_pmp_1_cfg_r,
  input [29:0] io_ptw_pmp_1_addr,
  input [31:0] io_ptw_pmp_1_mask,
  input io_ptw_pmp_2_cfg_l,
  input [1:0] io_ptw_pmp_2_cfg_a,
  input io_ptw_pmp_2_cfg_x,
  input io_ptw_pmp_2_cfg_w,
  input io_ptw_pmp_2_cfg_r,
  input [29:0] io_ptw_pmp_2_addr,
  input [31:0] io_ptw_pmp_2_mask,
  input io_ptw_pmp_3_cfg_l,
  input [1:0] io_ptw_pmp_3_cfg_a,
  input io_ptw_pmp_3_cfg_x,
  input io_ptw_pmp_3_cfg_w,
  input io_ptw_pmp_3_cfg_r,
  input [29:0] io_ptw_pmp_3_addr,
  input [31:0] io_ptw_pmp_3_mask,
  input io_ptw_pmp_4_cfg_l,
  input [1:0] io_ptw_pmp_4_cfg_a,
  input io_ptw_pmp_4_cfg_x,
  input io_ptw_pmp_4_cfg_w,
  input io_ptw_pmp_4_cfg_r,
  input [29:0] io_ptw_pmp_4_addr,
  input [31:0] io_ptw_pmp_4_mask,
  input io_ptw_pmp_5_cfg_l,
  input [1:0] io_ptw_pmp_5_cfg_a,
  input io_ptw_pmp_5_cfg_x,
  input io_ptw_pmp_5_cfg_w,
  input io_ptw_pmp_5_cfg_r,
  input [29:0] io_ptw_pmp_5_addr,
  input [31:0] io_ptw_pmp_5_mask,
  input io_ptw_pmp_6_cfg_l,
  input [1:0] io_ptw_pmp_6_cfg_a,
  input io_ptw_pmp_6_cfg_x,
  input io_ptw_pmp_6_cfg_w,
  input io_ptw_pmp_6_cfg_r,
  input [29:0] io_ptw_pmp_6_addr,
  input [31:0] io_ptw_pmp_6_mask,
  input io_ptw_pmp_7_cfg_l,
  input [1:0] io_ptw_pmp_7_cfg_a,
  input io_ptw_pmp_7_cfg_x,
  input io_ptw_pmp_7_cfg_w,
  input io_ptw_pmp_7_cfg_r,
  input [29:0] io_ptw_pmp_7_addr,
  input [31:0] io_ptw_pmp_7_mask,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [19:0] mpu_ppn_barrier_io_x_ppn ;  
   wire mpu_ppn_barrier_io_x_u ;  
   wire mpu_ppn_barrier_io_x_ae ;  
   wire mpu_ppn_barrier_io_x_sw ;  
   wire mpu_ppn_barrier_io_x_sx ;  
   wire mpu_ppn_barrier_io_x_sr ;  
   wire mpu_ppn_barrier_io_x_pw ;  
   wire mpu_ppn_barrier_io_x_px ;  
   wire mpu_ppn_barrier_io_x_pr ;  
   wire mpu_ppn_barrier_io_x_ppp ;  
   wire mpu_ppn_barrier_io_x_pal ;  
   wire mpu_ppn_barrier_io_x_paa ;  
   wire mpu_ppn_barrier_io_x_eff ;  
   wire mpu_ppn_barrier_io_x_c ;  
   wire [19:0] mpu_ppn_barrier_io_y_ppn ;  
   wire mpu_ppn_barrier_io_y_u ;  
   wire mpu_ppn_barrier_io_y_ae ;  
   wire mpu_ppn_barrier_io_y_sw ;  
   wire mpu_ppn_barrier_io_y_sx ;  
   wire mpu_ppn_barrier_io_y_sr ;  
   wire mpu_ppn_barrier_io_y_pw ;  
   wire mpu_ppn_barrier_io_y_px ;  
   wire mpu_ppn_barrier_io_y_pr ;  
   wire mpu_ppn_barrier_io_y_ppp ;  
   wire mpu_ppn_barrier_io_y_pal ;  
   wire mpu_ppn_barrier_io_y_paa ;  
   wire mpu_ppn_barrier_io_y_eff ;  
   wire mpu_ppn_barrier_io_y_c ;  
   wire [29:0] mpu_ppn_barrier_io_covSum ;  
   wire mpu_ppn_barrier_metaAssert ;  
   wire [1:0] pmp_io_prv ;  
   wire pmp_io_pmp_0_cfg_l ;  
   wire [1:0] pmp_io_pmp_0_cfg_a ;  
   wire pmp_io_pmp_0_cfg_x ;  
   wire pmp_io_pmp_0_cfg_w ;  
   wire pmp_io_pmp_0_cfg_r ;  
   wire [29:0] pmp_io_pmp_0_addr ;  
   wire [31:0] pmp_io_pmp_0_mask ;  
   wire pmp_io_pmp_1_cfg_l ;  
   wire [1:0] pmp_io_pmp_1_cfg_a ;  
   wire pmp_io_pmp_1_cfg_x ;  
   wire pmp_io_pmp_1_cfg_w ;  
   wire pmp_io_pmp_1_cfg_r ;  
   wire [29:0] pmp_io_pmp_1_addr ;  
   wire [31:0] pmp_io_pmp_1_mask ;  
   wire pmp_io_pmp_2_cfg_l ;  
   wire [1:0] pmp_io_pmp_2_cfg_a ;  
   wire pmp_io_pmp_2_cfg_x ;  
   wire pmp_io_pmp_2_cfg_w ;  
   wire pmp_io_pmp_2_cfg_r ;  
   wire [29:0] pmp_io_pmp_2_addr ;  
   wire [31:0] pmp_io_pmp_2_mask ;  
   wire pmp_io_pmp_3_cfg_l ;  
   wire [1:0] pmp_io_pmp_3_cfg_a ;  
   wire pmp_io_pmp_3_cfg_x ;  
   wire pmp_io_pmp_3_cfg_w ;  
   wire pmp_io_pmp_3_cfg_r ;  
   wire [29:0] pmp_io_pmp_3_addr ;  
   wire [31:0] pmp_io_pmp_3_mask ;  
   wire pmp_io_pmp_4_cfg_l ;  
   wire [1:0] pmp_io_pmp_4_cfg_a ;  
   wire pmp_io_pmp_4_cfg_x ;  
   wire pmp_io_pmp_4_cfg_w ;  
   wire pmp_io_pmp_4_cfg_r ;  
   wire [29:0] pmp_io_pmp_4_addr ;  
   wire [31:0] pmp_io_pmp_4_mask ;  
   wire pmp_io_pmp_5_cfg_l ;  
   wire [1:0] pmp_io_pmp_5_cfg_a ;  
   wire pmp_io_pmp_5_cfg_x ;  
   wire pmp_io_pmp_5_cfg_w ;  
   wire pmp_io_pmp_5_cfg_r ;  
   wire [29:0] pmp_io_pmp_5_addr ;  
   wire [31:0] pmp_io_pmp_5_mask ;  
   wire pmp_io_pmp_6_cfg_l ;  
   wire [1:0] pmp_io_pmp_6_cfg_a ;  
   wire pmp_io_pmp_6_cfg_x ;  
   wire pmp_io_pmp_6_cfg_w ;  
   wire pmp_io_pmp_6_cfg_r ;  
   wire [29:0] pmp_io_pmp_6_addr ;  
   wire [31:0] pmp_io_pmp_6_mask ;  
   wire pmp_io_pmp_7_cfg_l ;  
   wire [1:0] pmp_io_pmp_7_cfg_a ;  
   wire pmp_io_pmp_7_cfg_x ;  
   wire pmp_io_pmp_7_cfg_w ;  
   wire pmp_io_pmp_7_cfg_r ;  
   wire [29:0] pmp_io_pmp_7_addr ;  
   wire [31:0] pmp_io_pmp_7_mask ;  
   wire [31:0] pmp_io_addr ;  
   wire [1:0] pmp_io_size ;  
   wire pmp_io_r ;  
   wire pmp_io_w ;  
   wire pmp_io_x ;  
   wire [29:0] pmp_io_covSum ;  
   wire pmp_metaAssert ;  
   wire [19:0] entries_barrier_io_x_ppn ;  
   wire entries_barrier_io_x_u ;  
   wire entries_barrier_io_x_ae ;  
   wire entries_barrier_io_x_sw ;  
   wire entries_barrier_io_x_sx ;  
   wire entries_barrier_io_x_sr ;  
   wire entries_barrier_io_x_pw ;  
   wire entries_barrier_io_x_px ;  
   wire entries_barrier_io_x_pr ;  
   wire entries_barrier_io_x_ppp ;  
   wire entries_barrier_io_x_pal ;  
   wire entries_barrier_io_x_paa ;  
   wire entries_barrier_io_x_eff ;  
   wire entries_barrier_io_x_c ;  
   wire [19:0] entries_barrier_io_y_ppn ;  
   wire entries_barrier_io_y_u ;  
   wire entries_barrier_io_y_ae ;  
   wire entries_barrier_io_y_sw ;  
   wire entries_barrier_io_y_sx ;  
   wire entries_barrier_io_y_sr ;  
   wire entries_barrier_io_y_pw ;  
   wire entries_barrier_io_y_px ;  
   wire entries_barrier_io_y_pr ;  
   wire entries_barrier_io_y_ppp ;  
   wire entries_barrier_io_y_pal ;  
   wire entries_barrier_io_y_paa ;  
   wire entries_barrier_io_y_eff ;  
   wire entries_barrier_io_y_c ;  
   wire [29:0] entries_barrier_io_covSum ;  
   wire entries_barrier_metaAssert ;  
   wire [19:0] entries_barrier_1_io_x_ppn ;  
   wire entries_barrier_1_io_x_u ;  
   wire entries_barrier_1_io_x_ae ;  
   wire entries_barrier_1_io_x_sw ;  
   wire entries_barrier_1_io_x_sx ;  
   wire entries_barrier_1_io_x_sr ;  
   wire entries_barrier_1_io_x_pw ;  
   wire entries_barrier_1_io_x_px ;  
   wire entries_barrier_1_io_x_pr ;  
   wire entries_barrier_1_io_x_ppp ;  
   wire entries_barrier_1_io_x_pal ;  
   wire entries_barrier_1_io_x_paa ;  
   wire entries_barrier_1_io_x_eff ;  
   wire entries_barrier_1_io_x_c ;  
   wire [19:0] entries_barrier_1_io_y_ppn ;  
   wire entries_barrier_1_io_y_u ;  
   wire entries_barrier_1_io_y_ae ;  
   wire entries_barrier_1_io_y_sw ;  
   wire entries_barrier_1_io_y_sx ;  
   wire entries_barrier_1_io_y_sr ;  
   wire entries_barrier_1_io_y_pw ;  
   wire entries_barrier_1_io_y_px ;  
   wire entries_barrier_1_io_y_pr ;  
   wire entries_barrier_1_io_y_ppp ;  
   wire entries_barrier_1_io_y_pal ;  
   wire entries_barrier_1_io_y_paa ;  
   wire entries_barrier_1_io_y_eff ;  
   wire entries_barrier_1_io_y_c ;  
   wire [29:0] entries_barrier_1_io_covSum ;  
   wire entries_barrier_1_metaAssert ;  
   wire [19:0] entries_barrier_2_io_x_ppn ;  
   wire entries_barrier_2_io_x_u ;  
   wire entries_barrier_2_io_x_ae ;  
   wire entries_barrier_2_io_x_sw ;  
   wire entries_barrier_2_io_x_sx ;  
   wire entries_barrier_2_io_x_sr ;  
   wire entries_barrier_2_io_x_pw ;  
   wire entries_barrier_2_io_x_px ;  
   wire entries_barrier_2_io_x_pr ;  
   wire entries_barrier_2_io_x_ppp ;  
   wire entries_barrier_2_io_x_pal ;  
   wire entries_barrier_2_io_x_paa ;  
   wire entries_barrier_2_io_x_eff ;  
   wire entries_barrier_2_io_x_c ;  
   wire [19:0] entries_barrier_2_io_y_ppn ;  
   wire entries_barrier_2_io_y_u ;  
   wire entries_barrier_2_io_y_ae ;  
   wire entries_barrier_2_io_y_sw ;  
   wire entries_barrier_2_io_y_sx ;  
   wire entries_barrier_2_io_y_sr ;  
   wire entries_barrier_2_io_y_pw ;  
   wire entries_barrier_2_io_y_px ;  
   wire entries_barrier_2_io_y_pr ;  
   wire entries_barrier_2_io_y_ppp ;  
   wire entries_barrier_2_io_y_pal ;  
   wire entries_barrier_2_io_y_paa ;  
   wire entries_barrier_2_io_y_eff ;  
   wire entries_barrier_2_io_y_c ;  
   wire [29:0] entries_barrier_2_io_covSum ;  
   wire entries_barrier_2_metaAssert ;  
   wire [19:0] entries_barrier_3_io_x_ppn ;  
   wire entries_barrier_3_io_x_u ;  
   wire entries_barrier_3_io_x_ae ;  
   wire entries_barrier_3_io_x_sw ;  
   wire entries_barrier_3_io_x_sx ;  
   wire entries_barrier_3_io_x_sr ;  
   wire entries_barrier_3_io_x_pw ;  
   wire entries_barrier_3_io_x_px ;  
   wire entries_barrier_3_io_x_pr ;  
   wire entries_barrier_3_io_x_ppp ;  
   wire entries_barrier_3_io_x_pal ;  
   wire entries_barrier_3_io_x_paa ;  
   wire entries_barrier_3_io_x_eff ;  
   wire entries_barrier_3_io_x_c ;  
   wire [19:0] entries_barrier_3_io_y_ppn ;  
   wire entries_barrier_3_io_y_u ;  
   wire entries_barrier_3_io_y_ae ;  
   wire entries_barrier_3_io_y_sw ;  
   wire entries_barrier_3_io_y_sx ;  
   wire entries_barrier_3_io_y_sr ;  
   wire entries_barrier_3_io_y_pw ;  
   wire entries_barrier_3_io_y_px ;  
   wire entries_barrier_3_io_y_pr ;  
   wire entries_barrier_3_io_y_ppp ;  
   wire entries_barrier_3_io_y_pal ;  
   wire entries_barrier_3_io_y_paa ;  
   wire entries_barrier_3_io_y_eff ;  
   wire entries_barrier_3_io_y_c ;  
   wire [29:0] entries_barrier_3_io_covSum ;  
   wire entries_barrier_3_metaAssert ;  
   wire [19:0] entries_barrier_4_io_x_ppn ;  
   wire entries_barrier_4_io_x_u ;  
   wire entries_barrier_4_io_x_ae ;  
   wire entries_barrier_4_io_x_sw ;  
   wire entries_barrier_4_io_x_sx ;  
   wire entries_barrier_4_io_x_sr ;  
   wire entries_barrier_4_io_x_pw ;  
   wire entries_barrier_4_io_x_px ;  
   wire entries_barrier_4_io_x_pr ;  
   wire entries_barrier_4_io_x_ppp ;  
   wire entries_barrier_4_io_x_pal ;  
   wire entries_barrier_4_io_x_paa ;  
   wire entries_barrier_4_io_x_eff ;  
   wire entries_barrier_4_io_x_c ;  
   wire [19:0] entries_barrier_4_io_y_ppn ;  
   wire entries_barrier_4_io_y_u ;  
   wire entries_barrier_4_io_y_ae ;  
   wire entries_barrier_4_io_y_sw ;  
   wire entries_barrier_4_io_y_sx ;  
   wire entries_barrier_4_io_y_sr ;  
   wire entries_barrier_4_io_y_pw ;  
   wire entries_barrier_4_io_y_px ;  
   wire entries_barrier_4_io_y_pr ;  
   wire entries_barrier_4_io_y_ppp ;  
   wire entries_barrier_4_io_y_pal ;  
   wire entries_barrier_4_io_y_paa ;  
   wire entries_barrier_4_io_y_eff ;  
   wire entries_barrier_4_io_y_c ;  
   wire [29:0] entries_barrier_4_io_covSum ;  
   wire entries_barrier_4_metaAssert ;  
   wire [19:0] entries_barrier_5_io_x_ppn ;  
   wire entries_barrier_5_io_x_u ;  
   wire entries_barrier_5_io_x_ae ;  
   wire entries_barrier_5_io_x_sw ;  
   wire entries_barrier_5_io_x_sx ;  
   wire entries_barrier_5_io_x_sr ;  
   wire entries_barrier_5_io_x_pw ;  
   wire entries_barrier_5_io_x_px ;  
   wire entries_barrier_5_io_x_pr ;  
   wire entries_barrier_5_io_x_ppp ;  
   wire entries_barrier_5_io_x_pal ;  
   wire entries_barrier_5_io_x_paa ;  
   wire entries_barrier_5_io_x_eff ;  
   wire entries_barrier_5_io_x_c ;  
   wire [19:0] entries_barrier_5_io_y_ppn ;  
   wire entries_barrier_5_io_y_u ;  
   wire entries_barrier_5_io_y_ae ;  
   wire entries_barrier_5_io_y_sw ;  
   wire entries_barrier_5_io_y_sx ;  
   wire entries_barrier_5_io_y_sr ;  
   wire entries_barrier_5_io_y_pw ;  
   wire entries_barrier_5_io_y_px ;  
   wire entries_barrier_5_io_y_pr ;  
   wire entries_barrier_5_io_y_ppp ;  
   wire entries_barrier_5_io_y_pal ;  
   wire entries_barrier_5_io_y_paa ;  
   wire entries_barrier_5_io_y_eff ;  
   wire entries_barrier_5_io_y_c ;  
   wire [29:0] entries_barrier_5_io_covSum ;  
   wire entries_barrier_5_metaAssert ;  
   wire [19:0] entries_barrier_6_io_x_ppn ;  
   wire entries_barrier_6_io_x_u ;  
   wire entries_barrier_6_io_x_ae ;  
   wire entries_barrier_6_io_x_sw ;  
   wire entries_barrier_6_io_x_sx ;  
   wire entries_barrier_6_io_x_sr ;  
   wire entries_barrier_6_io_x_pw ;  
   wire entries_barrier_6_io_x_px ;  
   wire entries_barrier_6_io_x_pr ;  
   wire entries_barrier_6_io_x_ppp ;  
   wire entries_barrier_6_io_x_pal ;  
   wire entries_barrier_6_io_x_paa ;  
   wire entries_barrier_6_io_x_eff ;  
   wire entries_barrier_6_io_x_c ;  
   wire [19:0] entries_barrier_6_io_y_ppn ;  
   wire entries_barrier_6_io_y_u ;  
   wire entries_barrier_6_io_y_ae ;  
   wire entries_barrier_6_io_y_sw ;  
   wire entries_barrier_6_io_y_sx ;  
   wire entries_barrier_6_io_y_sr ;  
   wire entries_barrier_6_io_y_pw ;  
   wire entries_barrier_6_io_y_px ;  
   wire entries_barrier_6_io_y_pr ;  
   wire entries_barrier_6_io_y_ppp ;  
   wire entries_barrier_6_io_y_pal ;  
   wire entries_barrier_6_io_y_paa ;  
   wire entries_barrier_6_io_y_eff ;  
   wire entries_barrier_6_io_y_c ;  
   wire [29:0] entries_barrier_6_io_covSum ;  
   wire entries_barrier_6_metaAssert ;  
   wire [19:0] entries_barrier_7_io_x_ppn ;  
   wire entries_barrier_7_io_x_u ;  
   wire entries_barrier_7_io_x_ae ;  
   wire entries_barrier_7_io_x_sw ;  
   wire entries_barrier_7_io_x_sx ;  
   wire entries_barrier_7_io_x_sr ;  
   wire entries_barrier_7_io_x_pw ;  
   wire entries_barrier_7_io_x_px ;  
   wire entries_barrier_7_io_x_pr ;  
   wire entries_barrier_7_io_x_ppp ;  
   wire entries_barrier_7_io_x_pal ;  
   wire entries_barrier_7_io_x_paa ;  
   wire entries_barrier_7_io_x_eff ;  
   wire entries_barrier_7_io_x_c ;  
   wire [19:0] entries_barrier_7_io_y_ppn ;  
   wire entries_barrier_7_io_y_u ;  
   wire entries_barrier_7_io_y_ae ;  
   wire entries_barrier_7_io_y_sw ;  
   wire entries_barrier_7_io_y_sx ;  
   wire entries_barrier_7_io_y_sr ;  
   wire entries_barrier_7_io_y_pw ;  
   wire entries_barrier_7_io_y_px ;  
   wire entries_barrier_7_io_y_pr ;  
   wire entries_barrier_7_io_y_ppp ;  
   wire entries_barrier_7_io_y_pal ;  
   wire entries_barrier_7_io_y_paa ;  
   wire entries_barrier_7_io_y_eff ;  
   wire entries_barrier_7_io_y_c ;  
   wire [29:0] entries_barrier_7_io_covSum ;  
   wire entries_barrier_7_metaAssert ;  
   wire [19:0] entries_barrier_8_io_x_ppn ;  
   wire entries_barrier_8_io_x_u ;  
   wire entries_barrier_8_io_x_ae ;  
   wire entries_barrier_8_io_x_sw ;  
   wire entries_barrier_8_io_x_sx ;  
   wire entries_barrier_8_io_x_sr ;  
   wire entries_barrier_8_io_x_pw ;  
   wire entries_barrier_8_io_x_px ;  
   wire entries_barrier_8_io_x_pr ;  
   wire entries_barrier_8_io_x_ppp ;  
   wire entries_barrier_8_io_x_pal ;  
   wire entries_barrier_8_io_x_paa ;  
   wire entries_barrier_8_io_x_eff ;  
   wire entries_barrier_8_io_x_c ;  
   wire [19:0] entries_barrier_8_io_y_ppn ;  
   wire entries_barrier_8_io_y_u ;  
   wire entries_barrier_8_io_y_ae ;  
   wire entries_barrier_8_io_y_sw ;  
   wire entries_barrier_8_io_y_sx ;  
   wire entries_barrier_8_io_y_sr ;  
   wire entries_barrier_8_io_y_pw ;  
   wire entries_barrier_8_io_y_px ;  
   wire entries_barrier_8_io_y_pr ;  
   wire entries_barrier_8_io_y_ppp ;  
   wire entries_barrier_8_io_y_pal ;  
   wire entries_barrier_8_io_y_paa ;  
   wire entries_barrier_8_io_y_eff ;  
   wire entries_barrier_8_io_y_c ;  
   wire [29:0] entries_barrier_8_io_covSum ;  
   wire entries_barrier_8_metaAssert ;  
   wire [19:0] entries_barrier_9_io_x_ppn ;  
   wire entries_barrier_9_io_x_u ;  
   wire entries_barrier_9_io_x_ae ;  
   wire entries_barrier_9_io_x_sw ;  
   wire entries_barrier_9_io_x_sx ;  
   wire entries_barrier_9_io_x_sr ;  
   wire entries_barrier_9_io_x_pw ;  
   wire entries_barrier_9_io_x_px ;  
   wire entries_barrier_9_io_x_pr ;  
   wire entries_barrier_9_io_x_ppp ;  
   wire entries_barrier_9_io_x_pal ;  
   wire entries_barrier_9_io_x_paa ;  
   wire entries_barrier_9_io_x_eff ;  
   wire entries_barrier_9_io_x_c ;  
   wire [19:0] entries_barrier_9_io_y_ppn ;  
   wire entries_barrier_9_io_y_u ;  
   wire entries_barrier_9_io_y_ae ;  
   wire entries_barrier_9_io_y_sw ;  
   wire entries_barrier_9_io_y_sx ;  
   wire entries_barrier_9_io_y_sr ;  
   wire entries_barrier_9_io_y_pw ;  
   wire entries_barrier_9_io_y_px ;  
   wire entries_barrier_9_io_y_pr ;  
   wire entries_barrier_9_io_y_ppp ;  
   wire entries_barrier_9_io_y_pal ;  
   wire entries_barrier_9_io_y_paa ;  
   wire entries_barrier_9_io_y_eff ;  
   wire entries_barrier_9_io_y_c ;  
   wire [29:0] entries_barrier_9_io_covSum ;  
   wire entries_barrier_9_metaAssert ;  
   wire [19:0] entries_barrier_10_io_x_ppn ;  
   wire entries_barrier_10_io_x_u ;  
   wire entries_barrier_10_io_x_ae ;  
   wire entries_barrier_10_io_x_sw ;  
   wire entries_barrier_10_io_x_sx ;  
   wire entries_barrier_10_io_x_sr ;  
   wire entries_barrier_10_io_x_pw ;  
   wire entries_barrier_10_io_x_px ;  
   wire entries_barrier_10_io_x_pr ;  
   wire entries_barrier_10_io_x_ppp ;  
   wire entries_barrier_10_io_x_pal ;  
   wire entries_barrier_10_io_x_paa ;  
   wire entries_barrier_10_io_x_eff ;  
   wire entries_barrier_10_io_x_c ;  
   wire [19:0] entries_barrier_10_io_y_ppn ;  
   wire entries_barrier_10_io_y_u ;  
   wire entries_barrier_10_io_y_ae ;  
   wire entries_barrier_10_io_y_sw ;  
   wire entries_barrier_10_io_y_sx ;  
   wire entries_barrier_10_io_y_sr ;  
   wire entries_barrier_10_io_y_pw ;  
   wire entries_barrier_10_io_y_px ;  
   wire entries_barrier_10_io_y_pr ;  
   wire entries_barrier_10_io_y_ppp ;  
   wire entries_barrier_10_io_y_pal ;  
   wire entries_barrier_10_io_y_paa ;  
   wire entries_barrier_10_io_y_eff ;  
   wire entries_barrier_10_io_y_c ;  
   wire [29:0] entries_barrier_10_io_covSum ;  
   wire entries_barrier_10_metaAssert ;  
   wire [19:0] entries_barrier_11_io_x_ppn ;  
   wire entries_barrier_11_io_x_u ;  
   wire entries_barrier_11_io_x_ae ;  
   wire entries_barrier_11_io_x_sw ;  
   wire entries_barrier_11_io_x_sx ;  
   wire entries_barrier_11_io_x_sr ;  
   wire entries_barrier_11_io_x_pw ;  
   wire entries_barrier_11_io_x_px ;  
   wire entries_barrier_11_io_x_pr ;  
   wire entries_barrier_11_io_x_ppp ;  
   wire entries_barrier_11_io_x_pal ;  
   wire entries_barrier_11_io_x_paa ;  
   wire entries_barrier_11_io_x_eff ;  
   wire entries_barrier_11_io_x_c ;  
   wire [19:0] entries_barrier_11_io_y_ppn ;  
   wire entries_barrier_11_io_y_u ;  
   wire entries_barrier_11_io_y_ae ;  
   wire entries_barrier_11_io_y_sw ;  
   wire entries_barrier_11_io_y_sx ;  
   wire entries_barrier_11_io_y_sr ;  
   wire entries_barrier_11_io_y_pw ;  
   wire entries_barrier_11_io_y_px ;  
   wire entries_barrier_11_io_y_pr ;  
   wire entries_barrier_11_io_y_ppp ;  
   wire entries_barrier_11_io_y_pal ;  
   wire entries_barrier_11_io_y_paa ;  
   wire entries_barrier_11_io_y_eff ;  
   wire entries_barrier_11_io_y_c ;  
   wire [29:0] entries_barrier_11_io_covSum ;  
   wire entries_barrier_11_metaAssert ;  
   wire [19:0] entries_barrier_12_io_x_ppn ;  
   wire entries_barrier_12_io_x_u ;  
   wire entries_barrier_12_io_x_ae ;  
   wire entries_barrier_12_io_x_sw ;  
   wire entries_barrier_12_io_x_sx ;  
   wire entries_barrier_12_io_x_sr ;  
   wire entries_barrier_12_io_x_pw ;  
   wire entries_barrier_12_io_x_px ;  
   wire entries_barrier_12_io_x_pr ;  
   wire entries_barrier_12_io_x_ppp ;  
   wire entries_barrier_12_io_x_pal ;  
   wire entries_barrier_12_io_x_paa ;  
   wire entries_barrier_12_io_x_eff ;  
   wire entries_barrier_12_io_x_c ;  
   wire [19:0] entries_barrier_12_io_y_ppn ;  
   wire entries_barrier_12_io_y_u ;  
   wire entries_barrier_12_io_y_ae ;  
   wire entries_barrier_12_io_y_sw ;  
   wire entries_barrier_12_io_y_sx ;  
   wire entries_barrier_12_io_y_sr ;  
   wire entries_barrier_12_io_y_pw ;  
   wire entries_barrier_12_io_y_px ;  
   wire entries_barrier_12_io_y_pr ;  
   wire entries_barrier_12_io_y_ppp ;  
   wire entries_barrier_12_io_y_pal ;  
   wire entries_barrier_12_io_y_paa ;  
   wire entries_barrier_12_io_y_eff ;  
   wire entries_barrier_12_io_y_c ;  
   wire [29:0] entries_barrier_12_io_covSum ;  
   wire entries_barrier_12_metaAssert ;  
   wire [26:0] vpn ;  
   reg [26:0] sectored_entries_0_0_tag ;  
   reg [31:0] _RAND_0 ;  
   reg [34:0] sectored_entries_0_0_data_0 ;  
   reg [63:0] _RAND_1 ;  
   reg [34:0] sectored_entries_0_0_data_1 ;  
   reg [63:0] _RAND_2 ;  
   reg [34:0] sectored_entries_0_0_data_2 ;  
   reg [63:0] _RAND_3 ;  
   reg [34:0] sectored_entries_0_0_data_3 ;  
   reg [63:0] _RAND_4 ;  
   reg sectored_entries_0_0_valid_0 ;  
   reg [31:0] _RAND_5 ;  
   reg sectored_entries_0_0_valid_1 ;  
   reg [31:0] _RAND_6 ;  
   reg sectored_entries_0_0_valid_2 ;  
   reg [31:0] _RAND_7 ;  
   reg sectored_entries_0_0_valid_3 ;  
   reg [31:0] _RAND_8 ;  
   reg [26:0] sectored_entries_0_1_tag ;  
   reg [31:0] _RAND_9 ;  
   reg [34:0] sectored_entries_0_1_data_0 ;  
   reg [63:0] _RAND_10 ;  
   reg [34:0] sectored_entries_0_1_data_1 ;  
   reg [63:0] _RAND_11 ;  
   reg [34:0] sectored_entries_0_1_data_2 ;  
   reg [63:0] _RAND_12 ;  
   reg [34:0] sectored_entries_0_1_data_3 ;  
   reg [63:0] _RAND_13 ;  
   reg sectored_entries_0_1_valid_0 ;  
   reg [31:0] _RAND_14 ;  
   reg sectored_entries_0_1_valid_1 ;  
   reg [31:0] _RAND_15 ;  
   reg sectored_entries_0_1_valid_2 ;  
   reg [31:0] _RAND_16 ;  
   reg sectored_entries_0_1_valid_3 ;  
   reg [31:0] _RAND_17 ;  
   reg [26:0] sectored_entries_0_2_tag ;  
   reg [31:0] _RAND_18 ;  
   reg [34:0] sectored_entries_0_2_data_0 ;  
   reg [63:0] _RAND_19 ;  
   reg [34:0] sectored_entries_0_2_data_1 ;  
   reg [63:0] _RAND_20 ;  
   reg [34:0] sectored_entries_0_2_data_2 ;  
   reg [63:0] _RAND_21 ;  
   reg [34:0] sectored_entries_0_2_data_3 ;  
   reg [63:0] _RAND_22 ;  
   reg sectored_entries_0_2_valid_0 ;  
   reg [31:0] _RAND_23 ;  
   reg sectored_entries_0_2_valid_1 ;  
   reg [31:0] _RAND_24 ;  
   reg sectored_entries_0_2_valid_2 ;  
   reg [31:0] _RAND_25 ;  
   reg sectored_entries_0_2_valid_3 ;  
   reg [31:0] _RAND_26 ;  
   reg [26:0] sectored_entries_0_3_tag ;  
   reg [31:0] _RAND_27 ;  
   reg [34:0] sectored_entries_0_3_data_0 ;  
   reg [63:0] _RAND_28 ;  
   reg [34:0] sectored_entries_0_3_data_1 ;  
   reg [63:0] _RAND_29 ;  
   reg [34:0] sectored_entries_0_3_data_2 ;  
   reg [63:0] _RAND_30 ;  
   reg [34:0] sectored_entries_0_3_data_3 ;  
   reg [63:0] _RAND_31 ;  
   reg sectored_entries_0_3_valid_0 ;  
   reg [31:0] _RAND_32 ;  
   reg sectored_entries_0_3_valid_1 ;  
   reg [31:0] _RAND_33 ;  
   reg sectored_entries_0_3_valid_2 ;  
   reg [31:0] _RAND_34 ;  
   reg sectored_entries_0_3_valid_3 ;  
   reg [31:0] _RAND_35 ;  
   reg [26:0] sectored_entries_0_4_tag ;  
   reg [31:0] _RAND_36 ;  
   reg [34:0] sectored_entries_0_4_data_0 ;  
   reg [63:0] _RAND_37 ;  
   reg [34:0] sectored_entries_0_4_data_1 ;  
   reg [63:0] _RAND_38 ;  
   reg [34:0] sectored_entries_0_4_data_2 ;  
   reg [63:0] _RAND_39 ;  
   reg [34:0] sectored_entries_0_4_data_3 ;  
   reg [63:0] _RAND_40 ;  
   reg sectored_entries_0_4_valid_0 ;  
   reg [31:0] _RAND_41 ;  
   reg sectored_entries_0_4_valid_1 ;  
   reg [31:0] _RAND_42 ;  
   reg sectored_entries_0_4_valid_2 ;  
   reg [31:0] _RAND_43 ;  
   reg sectored_entries_0_4_valid_3 ;  
   reg [31:0] _RAND_44 ;  
   reg [26:0] sectored_entries_0_5_tag ;  
   reg [31:0] _RAND_45 ;  
   reg [34:0] sectored_entries_0_5_data_0 ;  
   reg [63:0] _RAND_46 ;  
   reg [34:0] sectored_entries_0_5_data_1 ;  
   reg [63:0] _RAND_47 ;  
   reg [34:0] sectored_entries_0_5_data_2 ;  
   reg [63:0] _RAND_48 ;  
   reg [34:0] sectored_entries_0_5_data_3 ;  
   reg [63:0] _RAND_49 ;  
   reg sectored_entries_0_5_valid_0 ;  
   reg [31:0] _RAND_50 ;  
   reg sectored_entries_0_5_valid_1 ;  
   reg [31:0] _RAND_51 ;  
   reg sectored_entries_0_5_valid_2 ;  
   reg [31:0] _RAND_52 ;  
   reg sectored_entries_0_5_valid_3 ;  
   reg [31:0] _RAND_53 ;  
   reg [26:0] sectored_entries_0_6_tag ;  
   reg [31:0] _RAND_54 ;  
   reg [34:0] sectored_entries_0_6_data_0 ;  
   reg [63:0] _RAND_55 ;  
   reg [34:0] sectored_entries_0_6_data_1 ;  
   reg [63:0] _RAND_56 ;  
   reg [34:0] sectored_entries_0_6_data_2 ;  
   reg [63:0] _RAND_57 ;  
   reg [34:0] sectored_entries_0_6_data_3 ;  
   reg [63:0] _RAND_58 ;  
   reg sectored_entries_0_6_valid_0 ;  
   reg [31:0] _RAND_59 ;  
   reg sectored_entries_0_6_valid_1 ;  
   reg [31:0] _RAND_60 ;  
   reg sectored_entries_0_6_valid_2 ;  
   reg [31:0] _RAND_61 ;  
   reg sectored_entries_0_6_valid_3 ;  
   reg [31:0] _RAND_62 ;  
   reg [26:0] sectored_entries_0_7_tag ;  
   reg [31:0] _RAND_63 ;  
   reg [34:0] sectored_entries_0_7_data_0 ;  
   reg [63:0] _RAND_64 ;  
   reg [34:0] sectored_entries_0_7_data_1 ;  
   reg [63:0] _RAND_65 ;  
   reg [34:0] sectored_entries_0_7_data_2 ;  
   reg [63:0] _RAND_66 ;  
   reg [34:0] sectored_entries_0_7_data_3 ;  
   reg [63:0] _RAND_67 ;  
   reg sectored_entries_0_7_valid_0 ;  
   reg [31:0] _RAND_68 ;  
   reg sectored_entries_0_7_valid_1 ;  
   reg [31:0] _RAND_69 ;  
   reg sectored_entries_0_7_valid_2 ;  
   reg [31:0] _RAND_70 ;  
   reg sectored_entries_0_7_valid_3 ;  
   reg [31:0] _RAND_71 ;  
   reg [1:0] superpage_entries_0_level ;  
   reg [31:0] _RAND_72 ;  
   reg [26:0] superpage_entries_0_tag ;  
   reg [31:0] _RAND_73 ;  
   reg [34:0] superpage_entries_0_data_0 ;  
   reg [63:0] _RAND_74 ;  
   reg superpage_entries_0_valid_0 ;  
   reg [31:0] _RAND_75 ;  
   reg [1:0] superpage_entries_1_level ;  
   reg [31:0] _RAND_76 ;  
   reg [26:0] superpage_entries_1_tag ;  
   reg [31:0] _RAND_77 ;  
   reg [34:0] superpage_entries_1_data_0 ;  
   reg [63:0] _RAND_78 ;  
   reg superpage_entries_1_valid_0 ;  
   reg [31:0] _RAND_79 ;  
   reg [1:0] superpage_entries_2_level ;  
   reg [31:0] _RAND_80 ;  
   reg [26:0] superpage_entries_2_tag ;  
   reg [31:0] _RAND_81 ;  
   reg [34:0] superpage_entries_2_data_0 ;  
   reg [63:0] _RAND_82 ;  
   reg superpage_entries_2_valid_0 ;  
   reg [31:0] _RAND_83 ;  
   reg [1:0] superpage_entries_3_level ;  
   reg [31:0] _RAND_84 ;  
   reg [26:0] superpage_entries_3_tag ;  
   reg [31:0] _RAND_85 ;  
   reg [34:0] superpage_entries_3_data_0 ;  
   reg [63:0] _RAND_86 ;  
   reg superpage_entries_3_valid_0 ;  
   reg [31:0] _RAND_87 ;  
   reg [1:0] special_entry_level ;  
   reg [31:0] _RAND_88 ;  
   reg [26:0] special_entry_tag ;  
   reg [31:0] _RAND_89 ;  
   reg [34:0] special_entry_data_0 ;  
   reg [63:0] _RAND_90 ;  
   reg special_entry_valid_0 ;  
   reg [31:0] _RAND_91 ;  
   reg [1:0] state ;  
   reg [31:0] _RAND_92 ;  
   reg [26:0] r_refill_tag ;  
   reg [31:0] _RAND_93 ;  
   reg [1:0] r_superpage_repl_addr ;  
   reg [31:0] _RAND_94 ;  
   reg [2:0] r_sectored_repl_addr ;  
   reg [31:0] _RAND_95 ;  
   reg [2:0] r_sectored_hit_addr ;  
   reg [31:0] _RAND_96 ;  
   reg r_sectored_hit ;  
   reg [31:0] _RAND_97 ;  
   wire priv_s ;  
   wire priv_uses_vm ;  
   wire _vm_enabled_T_2 ;  
   wire vm_enabled ;  
   wire [19:0] refill_ppn ;  
   wire _invalidate_refill_T ;  
   wire _invalidate_refill_T_1 ;  
   wire _invalidate_refill_T_2 ;  
   wire invalidate_refill ;  
   wire [1:0] mpu_ppn_hi ;  
   wire mpu_ppn_ignore ;  
   wire [26:0] _mpu_ppn_T_17 ;  
   wire [26:0] _GEN_919 ;  
   wire [26:0] _mpu_ppn_T_18 ;  
   wire [8:0] mpu_ppn_lo ;  
   wire mpu_ppn_ignore_1 ;  
   wire [26:0] _mpu_ppn_T_19 ;  
   wire [26:0] _mpu_ppn_T_20 ;  
   wire [8:0] mpu_ppn_lo_1 ;  
   wire [19:0] _mpu_ppn_T_21 ;  
   wire [27:0] _mpu_ppn_T_23 ;  
   wire [27:0] mpu_ppn ;  
   wire [11:0] mpu_physaddr_lo ;  
   wire [39:0] mpu_physaddr ;  
   wire _mpu_priv_T ;  
   wire [2:0] _mpu_priv_T_2 ;  
   wire [2:0] mpu_priv ;  
   wire [39:0] _legal_address_T ;  
   wire [40:0] _legal_address_T_1 ;  
   wire [40:0] _legal_address_T_3 ;  
   wire _legal_address_T_4 ;  
   wire [39:0] _legal_address_T_5 ;  
   wire [40:0] _legal_address_T_6 ;  
   wire [40:0] _legal_address_T_8 ;  
   wire _legal_address_T_9 ;  
   wire [39:0] _legal_address_T_10 ;  
   wire [40:0] _legal_address_T_11 ;  
   wire [40:0] _legal_address_T_13 ;  
   wire _legal_address_T_14 ;  
   wire [40:0] _legal_address_T_16 ;  
   wire [40:0] _legal_address_T_18 ;  
   wire _legal_address_T_19 ;  
   wire [39:0] _legal_address_T_20 ;  
   wire [40:0] _legal_address_T_21 ;  
   wire [40:0] _legal_address_T_23 ;  
   wire _legal_address_T_24 ;  
   wire [39:0] _legal_address_T_25 ;  
   wire [40:0] _legal_address_T_26 ;  
   wire [40:0] _legal_address_T_28 ;  
   wire _legal_address_T_29 ;  
   wire [39:0] _legal_address_T_30 ;  
   wire [40:0] _legal_address_T_31 ;  
   wire [40:0] _legal_address_T_33 ;  
   wire _legal_address_T_34 ;  
   wire _legal_address_T_35 ;  
   wire _legal_address_T_36 ;  
   wire _legal_address_T_37 ;  
   wire _legal_address_T_38 ;  
   wire _legal_address_T_39 ;  
   wire legal_address ;  
   wire [40:0] _cacheable_T_8 ;  
   wire _cacheable_T_9 ;  
   wire cacheable ;  
   wire [39:0] _homogeneous_T_54 ;  
   wire [40:0] _homogeneous_T_55 ;  
   wire [40:0] _homogeneous_T_57 ;  
   wire _homogeneous_T_58 ;  
   wire [40:0] _homogeneous_T_71 ;  
   wire _homogeneous_T_72 ;  
   wire _homogeneous_T_79 ;  
   wire _deny_access_to_debug_T ;  
   wire deny_access_to_debug ;  
   wire _prot_r_T_7 ;  
   wire prot_r ;  
   wire [39:0] _prot_w_T_10 ;  
   wire [40:0] _prot_w_T_11 ;  
   wire [40:0] _prot_w_T_13 ;  
   wire _prot_w_T_14 ;  
   wire [40:0] _prot_w_T_18 ;  
   wire _prot_w_T_19 ;  
   wire _prot_w_T_21 ;  
   wire _prot_w_T_22 ;  
   wire _prot_w_T_31 ;  
   wire _prot_w_T_33 ;  
   wire prot_w ;  
   wire prot_al ;  
   wire [40:0] _prot_x_T_3 ;  
   wire _prot_x_T_4 ;  
   wire _prot_x_T_15 ;  
   wire _prot_x_T_16 ;  
   wire _prot_x_T_31 ;  
   wire _prot_x_T_33 ;  
   wire prot_x ;  
   wire [40:0] _prot_eff_T_20 ;  
   wire _prot_eff_T_21 ;  
   wire [40:0] _prot_eff_T_25 ;  
   wire _prot_eff_T_26 ;  
   wire _prot_eff_T_37 ;  
   wire _prot_eff_T_38 ;  
   wire _prot_eff_T_39 ;  
   wire prot_eff ;  
   wire _sector_hits_T ;  
   wire _sector_hits_T_1 ;  
   wire _sector_hits_T_2 ;  
   wire [26:0] _sector_hits_T_3 ;  
   wire _sector_hits_T_5 ;  
   wire sector_hits_0 ;  
   wire _sector_hits_T_6 ;  
   wire _sector_hits_T_7 ;  
   wire _sector_hits_T_8 ;  
   wire [26:0] _sector_hits_T_9 ;  
   wire _sector_hits_T_11 ;  
   wire sector_hits_1 ;  
   wire _sector_hits_T_12 ;  
   wire _sector_hits_T_13 ;  
   wire _sector_hits_T_14 ;  
   wire [26:0] _sector_hits_T_15 ;  
   wire _sector_hits_T_17 ;  
   wire sector_hits_2 ;  
   wire _sector_hits_T_18 ;  
   wire _sector_hits_T_19 ;  
   wire _sector_hits_T_20 ;  
   wire [26:0] _sector_hits_T_21 ;  
   wire _sector_hits_T_23 ;  
   wire sector_hits_3 ;  
   wire _sector_hits_T_24 ;  
   wire _sector_hits_T_25 ;  
   wire _sector_hits_T_26 ;  
   wire [26:0] _sector_hits_T_27 ;  
   wire _sector_hits_T_29 ;  
   wire sector_hits_4 ;  
   wire _sector_hits_T_30 ;  
   wire _sector_hits_T_31 ;  
   wire _sector_hits_T_32 ;  
   wire [26:0] _sector_hits_T_33 ;  
   wire _sector_hits_T_35 ;  
   wire sector_hits_5 ;  
   wire _sector_hits_T_36 ;  
   wire _sector_hits_T_37 ;  
   wire _sector_hits_T_38 ;  
   wire [26:0] _sector_hits_T_39 ;  
   wire _sector_hits_T_41 ;  
   wire sector_hits_6 ;  
   wire _sector_hits_T_42 ;  
   wire _sector_hits_T_43 ;  
   wire _sector_hits_T_44 ;  
   wire [26:0] _sector_hits_T_45 ;  
   wire _sector_hits_T_47 ;  
   wire sector_hits_7 ;  
   wire _superpage_hits_T_2 ;  
   wire _superpage_hits_T_4 ;  
   wire superpage_hits_ignore_1 ;  
   wire _superpage_hits_T_7 ;  
   wire _superpage_hits_T_8 ;  
   wire superpage_hits_0 ;  
   wire _superpage_hits_T_16 ;  
   wire _superpage_hits_T_18 ;  
   wire superpage_hits_ignore_4 ;  
   wire _superpage_hits_T_21 ;  
   wire _superpage_hits_T_22 ;  
   wire superpage_hits_1 ;  
   wire _superpage_hits_T_30 ;  
   wire _superpage_hits_T_32 ;  
   wire superpage_hits_ignore_7 ;  
   wire _superpage_hits_T_35 ;  
   wire _superpage_hits_T_36 ;  
   wire superpage_hits_2 ;  
   wire _superpage_hits_T_44 ;  
   wire _superpage_hits_T_46 ;  
   wire superpage_hits_ignore_10 ;  
   wire _superpage_hits_T_49 ;  
   wire _superpage_hits_T_50 ;  
   wire superpage_hits_3 ;  
   wire [1:0] hitsVec_idx ;  
   wire _GEN_1 ;  
   wire _GEN_2 ;  
   wire _GEN_3 ;  
   wire _hitsVec_T_3 ;  
   wire hitsVec_0 ;  
   wire _GEN_5 ;  
   wire _GEN_6 ;  
   wire _GEN_7 ;  
   wire _hitsVec_T_7 ;  
   wire hitsVec_1 ;  
   wire _GEN_9 ;  
   wire _GEN_10 ;  
   wire _GEN_11 ;  
   wire _hitsVec_T_11 ;  
   wire hitsVec_2 ;  
   wire _GEN_13 ;  
   wire _GEN_14 ;  
   wire _GEN_15 ;  
   wire _hitsVec_T_15 ;  
   wire hitsVec_3 ;  
   wire _GEN_17 ;  
   wire _GEN_18 ;  
   wire _GEN_19 ;  
   wire _hitsVec_T_19 ;  
   wire hitsVec_4 ;  
   wire _GEN_21 ;  
   wire _GEN_22 ;  
   wire _GEN_23 ;  
   wire _hitsVec_T_23 ;  
   wire hitsVec_5 ;  
   wire _GEN_25 ;  
   wire _GEN_26 ;  
   wire _GEN_27 ;  
   wire _hitsVec_T_27 ;  
   wire hitsVec_6 ;  
   wire _GEN_29 ;  
   wire _GEN_30 ;  
   wire _GEN_31 ;  
   wire _hitsVec_T_31 ;  
   wire hitsVec_7 ;  
   wire hitsVec_8 ;  
   wire hitsVec_9 ;  
   wire hitsVec_10 ;  
   wire hitsVec_11 ;  
   wire _hitsVec_T_94 ;  
   wire _hitsVec_T_96 ;  
   wire _hitsVec_T_99 ;  
   wire _hitsVec_T_100 ;  
   wire _hitsVec_T_101 ;  
   wire _hitsVec_T_104 ;  
   wire _hitsVec_T_105 ;  
   wire _hitsVec_T_106 ;  
   wire hitsVec_12 ;  
   wire [5:0] real_hits_lo ;  
   wire [12:0] real_hits ;  
   wire hits_hi ;  
   wire [13:0] hits ;  
   wire newEntry_g ;  
   wire _newEntry_sr_T_1 ;  
   wire _newEntry_sr_T_2 ;  
   wire _newEntry_sr_T_3 ;  
   wire _newEntry_sr_T_4 ;  
   wire newEntry_sr ;  
   wire _newEntry_sw_T_5 ;  
   wire newEntry_sw ;  
   wire newEntry_sx ;  
   wire [7:0] special_entry_data_0_lo ;  
   wire [34:0] _special_entry_data_0_T ;  
   wire _GEN_32 ;  
   wire _T_2 ;  
   wire _T_3 ;  
   wire _GEN_35 ;  
   wire _T_4 ;  
   wire _GEN_39 ;  
   wire _T_5 ;  
   wire _GEN_43 ;  
   wire _T_6 ;  
   wire _GEN_47 ;  
   wire [2:0] waddr ;  
   wire _T_7 ;  
   wire _GEN_49 ;  
   wire _GEN_50 ;  
   wire _GEN_51 ;  
   wire _GEN_52 ;  
   wire [1:0] idx ;  
   wire _GEN_921 ;  
   wire _GEN_53 ;  
   wire _GEN_922 ;  
   wire _GEN_54 ;  
   wire _GEN_923 ;  
   wire _GEN_55 ;  
   wire _GEN_924 ;  
   wire _GEN_56 ;  
   wire _GEN_61 ;  
   wire _GEN_62 ;  
   wire _GEN_63 ;  
   wire _GEN_64 ;  
   wire _GEN_65 ;  
   wire _GEN_66 ;  
   wire _GEN_67 ;  
   wire _GEN_68 ;  
   wire _T_9 ;  
   wire _GEN_75 ;  
   wire _GEN_76 ;  
   wire _GEN_77 ;  
   wire _GEN_78 ;  
   wire _GEN_79 ;  
   wire _GEN_80 ;  
   wire _GEN_81 ;  
   wire _GEN_82 ;  
   wire _GEN_87 ;  
   wire _GEN_88 ;  
   wire _GEN_89 ;  
   wire _GEN_90 ;  
   wire _GEN_91 ;  
   wire _GEN_92 ;  
   wire _GEN_93 ;  
   wire _GEN_94 ;  
   wire _T_11 ;  
   wire _GEN_101 ;  
   wire _GEN_102 ;  
   wire _GEN_103 ;  
   wire _GEN_104 ;  
   wire _GEN_105 ;  
   wire _GEN_106 ;  
   wire _GEN_107 ;  
   wire _GEN_108 ;  
   wire _GEN_113 ;  
   wire _GEN_114 ;  
   wire _GEN_115 ;  
   wire _GEN_116 ;  
   wire _GEN_117 ;  
   wire _GEN_118 ;  
   wire _GEN_119 ;  
   wire _GEN_120 ;  
   wire _T_13 ;  
   wire _GEN_127 ;  
   wire _GEN_128 ;  
   wire _GEN_129 ;  
   wire _GEN_130 ;  
   wire _GEN_131 ;  
   wire _GEN_132 ;  
   wire _GEN_133 ;  
   wire _GEN_134 ;  
   wire _GEN_139 ;  
   wire _GEN_140 ;  
   wire _GEN_141 ;  
   wire _GEN_142 ;  
   wire _GEN_143 ;  
   wire _GEN_144 ;  
   wire _GEN_145 ;  
   wire _GEN_146 ;  
   wire _T_15 ;  
   wire _GEN_153 ;  
   wire _GEN_154 ;  
   wire _GEN_155 ;  
   wire _GEN_156 ;  
   wire _GEN_157 ;  
   wire _GEN_158 ;  
   wire _GEN_159 ;  
   wire _GEN_160 ;  
   wire _GEN_165 ;  
   wire _GEN_166 ;  
   wire _GEN_167 ;  
   wire _GEN_168 ;  
   wire _GEN_169 ;  
   wire _GEN_170 ;  
   wire _GEN_171 ;  
   wire _GEN_172 ;  
   wire _T_17 ;  
   wire _GEN_179 ;  
   wire _GEN_180 ;  
   wire _GEN_181 ;  
   wire _GEN_182 ;  
   wire _GEN_183 ;  
   wire _GEN_184 ;  
   wire _GEN_185 ;  
   wire _GEN_186 ;  
   wire _GEN_191 ;  
   wire _GEN_192 ;  
   wire _GEN_193 ;  
   wire _GEN_194 ;  
   wire _GEN_195 ;  
   wire _GEN_196 ;  
   wire _GEN_197 ;  
   wire _GEN_198 ;  
   wire _T_19 ;  
   wire _GEN_205 ;  
   wire _GEN_206 ;  
   wire _GEN_207 ;  
   wire _GEN_208 ;  
   wire _GEN_209 ;  
   wire _GEN_210 ;  
   wire _GEN_211 ;  
   wire _GEN_212 ;  
   wire _GEN_217 ;  
   wire _GEN_218 ;  
   wire _GEN_219 ;  
   wire _GEN_220 ;  
   wire _GEN_221 ;  
   wire _GEN_222 ;  
   wire _GEN_223 ;  
   wire _GEN_224 ;  
   wire _T_21 ;  
   wire _GEN_231 ;  
   wire _GEN_232 ;  
   wire _GEN_233 ;  
   wire _GEN_234 ;  
   wire _GEN_235 ;  
   wire _GEN_236 ;  
   wire _GEN_237 ;  
   wire _GEN_238 ;  
   wire _GEN_243 ;  
   wire _GEN_244 ;  
   wire _GEN_245 ;  
   wire _GEN_246 ;  
   wire _GEN_247 ;  
   wire _GEN_248 ;  
   wire _GEN_249 ;  
   wire _GEN_250 ;  
   wire _GEN_259 ;  
   wire _GEN_263 ;  
   wire _GEN_267 ;  
   wire _GEN_271 ;  
   wire _GEN_273 ;  
   wire _GEN_274 ;  
   wire _GEN_275 ;  
   wire _GEN_276 ;  
   wire _GEN_283 ;  
   wire _GEN_284 ;  
   wire _GEN_285 ;  
   wire _GEN_286 ;  
   wire _GEN_293 ;  
   wire _GEN_294 ;  
   wire _GEN_295 ;  
   wire _GEN_296 ;  
   wire _GEN_303 ;  
   wire _GEN_304 ;  
   wire _GEN_305 ;  
   wire _GEN_306 ;  
   wire _GEN_313 ;  
   wire _GEN_314 ;  
   wire _GEN_315 ;  
   wire _GEN_316 ;  
   wire _GEN_323 ;  
   wire _GEN_324 ;  
   wire _GEN_325 ;  
   wire _GEN_326 ;  
   wire _GEN_333 ;  
   wire _GEN_334 ;  
   wire _GEN_335 ;  
   wire _GEN_336 ;  
   wire _GEN_343 ;  
   wire _GEN_344 ;  
   wire _GEN_345 ;  
   wire _GEN_346 ;  
   wire _GEN_355 ;  
   wire _GEN_359 ;  
   wire _GEN_363 ;  
   wire _GEN_367 ;  
   wire _GEN_371 ;  
   wire _GEN_373 ;  
   wire _GEN_374 ;  
   wire _GEN_375 ;  
   wire _GEN_376 ;  
   wire _GEN_383 ;  
   wire _GEN_384 ;  
   wire _GEN_385 ;  
   wire _GEN_386 ;  
   wire _GEN_393 ;  
   wire _GEN_394 ;  
   wire _GEN_395 ;  
   wire _GEN_396 ;  
   wire _GEN_403 ;  
   wire _GEN_404 ;  
   wire _GEN_405 ;  
   wire _GEN_406 ;  
   wire _GEN_413 ;  
   wire _GEN_414 ;  
   wire _GEN_415 ;  
   wire _GEN_416 ;  
   wire _GEN_423 ;  
   wire _GEN_424 ;  
   wire _GEN_425 ;  
   wire _GEN_426 ;  
   wire _GEN_433 ;  
   wire _GEN_434 ;  
   wire _GEN_435 ;  
   wire _GEN_436 ;  
   wire _GEN_443 ;  
   wire _GEN_444 ;  
   wire _GEN_445 ;  
   wire _GEN_446 ;  
   wire _GEN_455 ;  
   wire _GEN_459 ;  
   wire _GEN_463 ;  
   wire _GEN_467 ;  
   wire _GEN_471 ;  
   wire _GEN_473 ;  
   wire _GEN_474 ;  
   wire _GEN_475 ;  
   wire _GEN_476 ;  
   wire _GEN_483 ;  
   wire _GEN_484 ;  
   wire _GEN_485 ;  
   wire _GEN_486 ;  
   wire _GEN_493 ;  
   wire _GEN_494 ;  
   wire _GEN_495 ;  
   wire _GEN_496 ;  
   wire _GEN_503 ;  
   wire _GEN_504 ;  
   wire _GEN_505 ;  
   wire _GEN_506 ;  
   wire _GEN_513 ;  
   wire _GEN_514 ;  
   wire _GEN_515 ;  
   wire _GEN_516 ;  
   wire _GEN_523 ;  
   wire _GEN_524 ;  
   wire _GEN_525 ;  
   wire _GEN_526 ;  
   wire _GEN_533 ;  
   wire _GEN_534 ;  
   wire _GEN_535 ;  
   wire _GEN_536 ;  
   wire _GEN_543 ;  
   wire _GEN_544 ;  
   wire _GEN_545 ;  
   wire _GEN_546 ;  
   wire [34:0] _GEN_554 ;  
   wire [34:0] _GEN_555 ;  
   wire [34:0] _GEN_556 ;  
   wire [34:0] _GEN_558 ;  
   wire [34:0] _GEN_559 ;  
   wire [34:0] _GEN_560 ;  
   wire [34:0] _GEN_562 ;  
   wire [34:0] _GEN_563 ;  
   wire [34:0] _GEN_564 ;  
   wire [34:0] _GEN_566 ;  
   wire [34:0] _GEN_567 ;  
   wire [34:0] _GEN_568 ;  
   wire [34:0] _GEN_570 ;  
   wire [34:0] _GEN_571 ;  
   wire [34:0] _GEN_572 ;  
   wire [34:0] _GEN_574 ;  
   wire [34:0] _GEN_575 ;  
   wire [34:0] _GEN_576 ;  
   wire [34:0] _GEN_578 ;  
   wire [34:0] _GEN_579 ;  
   wire [34:0] _GEN_580 ;  
   wire [34:0] _GEN_582 ;  
   wire [34:0] _GEN_583 ;  
   wire [34:0] _GEN_584 ;  
   wire [1:0] ppn_hi ;  
   wire [26:0] _ppn_T_1 ;  
   wire [26:0] _GEN_953 ;  
   wire [26:0] _ppn_T_2 ;  
   wire [8:0] ppn_lo ;  
   wire [26:0] _ppn_T_4 ;  
   wire [8:0] ppn_lo_1 ;  
   wire [19:0] _ppn_T_5 ;  
   wire [1:0] ppn_hi_2 ;  
   wire [26:0] _ppn_T_6 ;  
   wire [26:0] _GEN_955 ;  
   wire [26:0] _ppn_T_7 ;  
   wire [8:0] ppn_lo_2 ;  
   wire [26:0] _ppn_T_9 ;  
   wire [8:0] ppn_lo_3 ;  
   wire [19:0] _ppn_T_10 ;  
   wire [1:0] ppn_hi_4 ;  
   wire [26:0] _ppn_T_11 ;  
   wire [26:0] _GEN_957 ;  
   wire [26:0] _ppn_T_12 ;  
   wire [8:0] ppn_lo_4 ;  
   wire [26:0] _ppn_T_14 ;  
   wire [8:0] ppn_lo_5 ;  
   wire [19:0] _ppn_T_15 ;  
   wire [1:0] ppn_hi_6 ;  
   wire [26:0] _ppn_T_16 ;  
   wire [26:0] _GEN_959 ;  
   wire [26:0] _ppn_T_17 ;  
   wire [8:0] ppn_lo_6 ;  
   wire [26:0] _ppn_T_19 ;  
   wire [8:0] ppn_lo_7 ;  
   wire [19:0] _ppn_T_20 ;  
   wire [1:0] ppn_hi_8 ;  
   wire [26:0] _GEN_961 ;  
   wire [26:0] _ppn_T_22 ;  
   wire [8:0] ppn_lo_8 ;  
   wire [26:0] _ppn_T_24 ;  
   wire [8:0] ppn_lo_9 ;  
   wire [19:0] _ppn_T_25 ;  
   wire [19:0] _ppn_T_27 ;  
   wire [19:0] _ppn_T_28 ;  
   wire [19:0] _ppn_T_29 ;  
   wire [19:0] _ppn_T_30 ;  
   wire [19:0] _ppn_T_31 ;  
   wire [19:0] _ppn_T_32 ;  
   wire [19:0] _ppn_T_33 ;  
   wire [19:0] _ppn_T_34 ;  
   wire [19:0] _ppn_T_35 ;  
   wire [19:0] _ppn_T_36 ;  
   wire [19:0] _ppn_T_37 ;  
   wire [19:0] _ppn_T_38 ;  
   wire [19:0] _ppn_T_39 ;  
   wire [19:0] _ppn_T_40 ;  
   wire [19:0] _ppn_T_41 ;  
   wire [19:0] _ppn_T_42 ;  
   wire [19:0] _ppn_T_43 ;  
   wire [19:0] _ppn_T_44 ;  
   wire [19:0] _ppn_T_45 ;  
   wire [19:0] _ppn_T_46 ;  
   wire [19:0] _ppn_T_47 ;  
   wire [19:0] _ppn_T_48 ;  
   wire [19:0] _ppn_T_49 ;  
   wire [19:0] _ppn_T_50 ;  
   wire [19:0] _ppn_T_51 ;  
   wire [19:0] _ppn_T_52 ;  
   wire [19:0] ppn ;  
   wire [5:0] ptw_ae_array_lo ;  
   wire [13:0] ptw_ae_array ;  
   wire _priv_rw_ok_T_1 ;  
   wire [5:0] priv_rw_ok_lo ;  
   wire [12:0] _priv_rw_ok_T_2 ;  
   wire [12:0] _priv_rw_ok_T_3 ;  
   wire [12:0] _priv_rw_ok_T_6 ;  
   wire [12:0] priv_rw_ok ;  
   wire [5:0] r_array_lo ;  
   wire [12:0] _r_array_T ;  
   wire [5:0] r_array_lo_1 ;  
   wire [12:0] _r_array_T_1 ;  
   wire [12:0] _r_array_T_2 ;  
   wire [12:0] _r_array_T_3 ;  
   wire [12:0] r_array_lo_2 ;  
   wire [13:0] r_array ;  
   wire [5:0] w_array_lo ;  
   wire [12:0] _w_array_T ;  
   wire [12:0] w_array_lo_1 ;  
   wire [13:0] w_array ;  
   wire [1:0] pr_array_hi ;  
   wire [5:0] pr_array_lo ;  
   wire [13:0] _pr_array_T_1 ;  
   wire [13:0] pr_array ;  
   wire [1:0] pw_array_hi ;  
   wire [5:0] pw_array_lo ;  
   wire [13:0] _pw_array_T_1 ;  
   wire [13:0] pw_array ;  
   wire [1:0] eff_array_hi ;  
   wire [5:0] eff_array_lo ;  
   wire [13:0] eff_array ;  
   wire [1:0] c_array_hi ;  
   wire [5:0] c_array_lo ;  
   wire [13:0] c_array ;  
   wire [1:0] ppp_array_hi ;  
   wire [5:0] ppp_array_lo ;  
   wire [13:0] ppp_array ;  
   wire [1:0] paa_array_hi ;  
   wire [5:0] paa_array_lo ;  
   wire [13:0] paa_array ;  
   wire [5:0] pal_array_lo ;  
   wire [13:0] pal_array ;  
   wire [13:0] ppp_array_if_cached ;  
   wire [13:0] paa_array_if_cached ;  
   wire [13:0] pal_array_if_cached ;  
   wire [3:0] _misaligned_T ;  
   wire [3:0] _misaligned_T_2 ;  
   wire [39:0] _GEN_963 ;  
   wire [39:0] _misaligned_T_3 ;  
   wire misaligned ;  
   wire [39:0] bad_va_maskedVAddr ;  
   wire _bad_va_T_1 ;  
   wire _bad_va_T_2 ;  
   wire _bad_va_T_3 ;  
   wire bad_va ;  
   wire _cmd_lrsc_T ;  
   wire _cmd_lrsc_T_1 ;  
   wire cmd_lrsc ;  
   wire _cmd_amo_logical_T ;  
   wire _cmd_amo_logical_T_1 ;  
   wire _cmd_amo_logical_T_2 ;  
   wire _cmd_amo_logical_T_3 ;  
   wire _cmd_amo_logical_T_4 ;  
   wire _cmd_amo_logical_T_5 ;  
   wire cmd_amo_logical ;  
   wire _cmd_amo_arithmetic_T ;  
   wire _cmd_amo_arithmetic_T_1 ;  
   wire _cmd_amo_arithmetic_T_2 ;  
   wire _cmd_amo_arithmetic_T_3 ;  
   wire _cmd_amo_arithmetic_T_4 ;  
   wire _cmd_amo_arithmetic_T_5 ;  
   wire _cmd_amo_arithmetic_T_6 ;  
   wire _cmd_amo_arithmetic_T_7 ;  
   wire cmd_amo_arithmetic ;  
   wire cmd_put_partial ;  
   wire _cmd_read_T ;  
   wire _cmd_read_T_2 ;  
   wire _cmd_read_T_4 ;  
   wire _cmd_read_T_21 ;  
   wire cmd_read ;  
   wire _cmd_write_T ;  
   wire _cmd_write_T_2 ;  
   wire _cmd_write_T_4 ;  
   wire cmd_write ;  
   wire _cmd_write_perms_T ;  
   wire _cmd_write_perms_T_1 ;  
   wire _cmd_write_perms_T_2 ;  
   wire cmd_write_perms ;  
   wire [13:0] _ae_array_T ;  
   wire [13:0] _ae_array_T_2 ;  
   wire [13:0] ae_array ;  
   wire [13:0] _ae_ld_array_T_1 ;  
   wire [13:0] ae_ld_array ;  
   wire [13:0] _ae_st_array_T_1 ;  
   wire [13:0] _ae_st_array_T_2 ;  
   wire [13:0] _ae_st_array_T_4 ;  
   wire [13:0] _ae_st_array_T_5 ;  
   wire [13:0] _ae_st_array_T_7 ;  
   wire [13:0] _ae_st_array_T_8 ;  
   wire [13:0] _ae_st_array_T_10 ;  
   wire [13:0] ae_st_array ;  
   wire _ma_ld_array_T ;  
   wire [13:0] ma_ld_array ;  
   wire _ma_st_array_T ;  
   wire [13:0] ma_st_array ;  
   wire [13:0] _pf_ld_array_T ;  
   wire [13:0] pf_ld_array ;  
   wire [13:0] _pf_st_array_T ;  
   wire [13:0] pf_st_array ;  
   wire tlb_hit ;  
   wire _tlb_miss_T_1 ;  
   wire tlb_miss ;  
   reg [6:0] state_vec_0 ;  
   reg [31:0] _RAND_98 ;  
   reg [2:0] state_reg_1 ;  
   reg [31:0] _RAND_99 ;  
   wire _T_23 ;  
   wire _T_24 ;  
   wire _T_25 ;  
   wire _T_26 ;  
   wire _T_27 ;  
   wire _T_28 ;  
   wire _T_29 ;  
   wire _T_30 ;  
   wire [7:0] _T_31 ;  
   wire [3:0] hi_1 ;  
   wire [3:0] lo_1 ;  
   wire hi_2 ;  
   wire [3:0] _T_32 ;  
   wire [1:0] hi_3 ;  
   wire [1:0] lo_2 ;  
   wire hi_4 ;  
   wire [1:0] _T_33 ;  
   wire lo_3 ;  
   wire [2:0] state_vec_0_touch_way_sized ;  
   wire state_vec_0_hi_hi ;  
   wire [2:0] state_vec_0_left_subtree_state ;  
   wire [2:0] state_vec_0_right_subtree_state ;  
   wire state_vec_0_hi_hi_1 ;  
   wire state_vec_0_left_subtree_state_1 ;  
   wire state_vec_0_right_subtree_state_1 ;  
   wire state_vec_0_hi_lo ;  
   wire state_vec_0_lo ;  
   wire [2:0] _state_vec_0_T_7 ;  
   wire [2:0] state_vec_0_hi_lo_1 ;  
   wire state_vec_0_left_subtree_state_2 ;  
   wire state_vec_0_right_subtree_state_2 ;  
   wire state_vec_0_hi_lo_2 ;  
   wire state_vec_0_lo_1 ;  
   wire [2:0] _state_vec_0_T_15 ;  
   wire [2:0] state_vec_0_lo_2 ;  
   wire [6:0] _state_vec_0_T_16 ;  
   wire _T_35 ;  
   wire _T_36 ;  
   wire _T_37 ;  
   wire [3:0] _T_38 ;  
   wire [1:0] hi_6 ;  
   wire [1:0] lo_6 ;  
   wire hi_7 ;  
   wire [1:0] _T_39 ;  
   wire lo_7 ;  
   wire [1:0] state_reg_touch_way_sized ;  
   wire state_reg_hi_hi ;  
   wire state_reg_left_subtree_state ;  
   wire state_reg_right_subtree_state ;  
   wire state_reg_hi_lo ;  
   wire state_reg_lo ;  
   wire [2:0] _state_reg_T_6 ;  
   wire multipleHits_leftOne ;  
   wire multipleHits_leftOne_1 ;  
   wire multipleHits_rightOne ;  
   wire multipleHits_rightOne_1 ;  
   wire multipleHits_rightTwo ;  
   wire multipleHits_leftOne_2 ;  
   wire _multipleHits_T_9 ;  
   wire multipleHits_leftTwo ;  
   wire multipleHits_leftOne_3 ;  
   wire multipleHits_leftOne_4 ;  
   wire multipleHits_rightOne_2 ;  
   wire multipleHits_rightOne_3 ;  
   wire multipleHits_rightTwo_1 ;  
   wire multipleHits_rightOne_4 ;  
   wire _multipleHits_T_18 ;  
   wire multipleHits_rightTwo_2 ;  
   wire multipleHits_leftOne_5 ;  
   wire _multipleHits_T_19 ;  
   wire _multipleHits_T_20 ;  
   wire multipleHits_leftTwo_1 ;  
   wire multipleHits_leftOne_6 ;  
   wire multipleHits_leftOne_7 ;  
   wire multipleHits_rightOne_5 ;  
   wire multipleHits_rightOne_6 ;  
   wire multipleHits_rightTwo_3 ;  
   wire multipleHits_leftOne_8 ;  
   wire _multipleHits_T_30 ;  
   wire multipleHits_leftTwo_2 ;  
   wire multipleHits_leftOne_9 ;  
   wire multipleHits_rightOne_7 ;  
   wire multipleHits_leftOne_10 ;  
   wire multipleHits_leftTwo_3 ;  
   wire multipleHits_leftOne_11 ;  
   wire multipleHits_rightOne_8 ;  
   wire multipleHits_rightOne_9 ;  
   wire multipleHits_rightTwo_4 ;  
   wire multipleHits_rightOne_10 ;  
   wire _multipleHits_T_42 ;  
   wire _multipleHits_T_43 ;  
   wire multipleHits_rightTwo_5 ;  
   wire multipleHits_rightOne_11 ;  
   wire _multipleHits_T_44 ;  
   wire _multipleHits_T_45 ;  
   wire multipleHits_rightTwo_6 ;  
   wire _multipleHits_T_47 ;  
   wire _multipleHits_T_48 ;  
   wire multipleHits ;  
   wire _io_resp_pf_ld_T ;  
   wire [13:0] _io_resp_pf_ld_T_1 ;  
   wire _io_resp_pf_ld_T_2 ;  
   wire _io_resp_pf_st_T ;  
   wire [13:0] _io_resp_pf_st_T_1 ;  
   wire _io_resp_pf_st_T_2 ;  
   wire [13:0] _io_resp_ae_ld_T ;  
   wire [13:0] _io_resp_ae_st_T ;  
   wire [13:0] _io_resp_ma_ld_T ;  
   wire [13:0] _io_resp_ma_st_T ;  
   wire [13:0] _io_resp_cacheable_T ;  
   wire _io_resp_miss_T ;  
   wire _T_41 ;  
   wire _T_42 ;  
   wire r_superpage_repl_addr_hi ;  
   wire r_superpage_repl_addr_lo ;  
   wire [1:0] _r_superpage_repl_addr_T_2 ;  
   wire [3:0] r_superpage_repl_addr_valids ;  
   wire _r_superpage_repl_addr_T_3 ;  
   wire _r_superpage_repl_addr_T_5 ;  
   wire _r_superpage_repl_addr_T_6 ;  
   wire _r_superpage_repl_addr_T_7 ;  
   wire r_sectored_repl_addr_hi ;  
   wire r_sectored_repl_addr_hi_1 ;  
   wire r_sectored_repl_addr_lo ;  
   wire [1:0] _r_sectored_repl_addr_T_2 ;  
   wire r_sectored_repl_addr_hi_2 ;  
   wire r_sectored_repl_addr_lo_1 ;  
   wire [1:0] _r_sectored_repl_addr_T_5 ;  
   wire [1:0] r_sectored_repl_addr_lo_2 ;  
   wire [2:0] _r_sectored_repl_addr_T_6 ;  
   wire [7:0] r_sectored_repl_addr_valids ;  
   wire _r_sectored_repl_addr_T_7 ;  
   wire _r_sectored_repl_addr_T_9 ;  
   wire _r_sectored_repl_addr_T_10 ;  
   wire _r_sectored_repl_addr_T_11 ;  
   wire _r_sectored_repl_addr_T_12 ;  
   wire _r_sectored_repl_addr_T_13 ;  
   wire _r_sectored_repl_addr_T_14 ;  
   wire _r_sectored_repl_addr_T_15 ;  
   wire _T_44 ;  
   wire _T_45 ;  
   wire _T_48 ;  
   wire _T_49 ;  
   wire _T_51 ;  
   wire _T_59 ;  
   wire _GEN_617 ;  
   wire _GEN_618 ;  
   wire _GEN_619 ;  
   wire _GEN_620 ;  
   wire _GEN_621 ;  
   wire _GEN_622 ;  
   wire _GEN_623 ;  
   wire _GEN_624 ;  
   wire _T_198 ;  
   wire _GEN_645 ;  
   wire _GEN_646 ;  
   wire _GEN_647 ;  
   wire _GEN_648 ;  
   wire _GEN_649 ;  
   wire _GEN_650 ;  
   wire _GEN_651 ;  
   wire _GEN_652 ;  
   wire _T_337 ;  
   wire _GEN_673 ;  
   wire _GEN_674 ;  
   wire _GEN_675 ;  
   wire _GEN_676 ;  
   wire _GEN_677 ;  
   wire _GEN_678 ;  
   wire _GEN_679 ;  
   wire _GEN_680 ;  
   wire _T_476 ;  
   wire _GEN_701 ;  
   wire _GEN_702 ;  
   wire _GEN_703 ;  
   wire _GEN_704 ;  
   wire _GEN_705 ;  
   wire _GEN_706 ;  
   wire _GEN_707 ;  
   wire _GEN_708 ;  
   wire _T_615 ;  
   wire _GEN_729 ;  
   wire _GEN_730 ;  
   wire _GEN_731 ;  
   wire _GEN_732 ;  
   wire _GEN_733 ;  
   wire _GEN_734 ;  
   wire _GEN_735 ;  
   wire _GEN_736 ;  
   wire _T_754 ;  
   wire _GEN_757 ;  
   wire _GEN_758 ;  
   wire _GEN_759 ;  
   wire _GEN_760 ;  
   wire _GEN_761 ;  
   wire _GEN_762 ;  
   wire _GEN_763 ;  
   wire _GEN_764 ;  
   wire _T_893 ;  
   wire _GEN_785 ;  
   wire _GEN_786 ;  
   wire _GEN_787 ;  
   wire _GEN_788 ;  
   wire _GEN_789 ;  
   wire _GEN_790 ;  
   wire _GEN_791 ;  
   wire _GEN_792 ;  
   wire _T_1032 ;  
   wire _GEN_813 ;  
   wire _GEN_814 ;  
   wire _GEN_815 ;  
   wire _GEN_816 ;  
   wire _GEN_817 ;  
   wire _GEN_818 ;  
   wire _GEN_819 ;  
   wire _GEN_820 ;  
   wire _GEN_826 ;  
   wire _GEN_827 ;  
   wire _GEN_830 ;  
   wire _GEN_831 ;  
   wire _GEN_834 ;  
   wire _GEN_835 ;  
   wire _GEN_838 ;  
   wire _GEN_839 ;  
   wire _GEN_842 ;  
   wire _GEN_843 ;  
   wire _T_1326 ;  
   reg [19:0] TLB_state ;  
   reg [31:0] _RAND_100 ;  
   reg TLB_cov[0:1048575] ;  
   reg [31:0] _RAND_101 ;  
   wire TLB_cov_read_data ;  
   wire [19:0] TLB_cov_read_addr ;  
   wire TLB_cov_write_data ;  
   wire [19:0] TLB_cov_write_addr ;  
   wire TLB_cov_write_mask ;  
   wire TLB_cov_write_en ;  
   reg [29:0] TLB_covSum ;  
   reg [31:0] _RAND_102 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire mux_cond_4 ;  
   wire mux_cond_5 ;  
   wire mux_cond_6 ;  
   wire mux_cond_7 ;  
   wire mux_cond_8 ;  
   wire mux_cond_9 ;  
   wire mux_cond_10 ;  
   wire mux_cond_11 ;  
   wire mux_cond_12 ;  
   wire mux_cond_13 ;  
   wire mux_cond_14 ;  
   wire mux_cond_15 ;  
   wire mux_cond_16 ;  
   wire mux_cond_17 ;  
   wire mux_cond_18 ;  
   wire mux_cond_19 ;  
   wire mux_cond_20 ;  
   wire mux_cond_21 ;  
   wire mux_cond_22 ;  
   wire mux_cond_23 ;  
   wire mux_cond_24 ;  
   wire mux_cond_25 ;  
   wire mux_cond_26 ;  
   wire mux_cond_27 ;  
   wire mux_cond_28 ;  
   wire mux_cond_29 ;  
   wire mux_cond_30 ;  
   wire mux_cond_31 ;  
   wire mux_cond_32 ;  
   wire mux_cond_33 ;  
   wire mux_cond_34 ;  
   wire mux_cond_35 ;  
   wire mux_cond_36 ;  
   wire mux_cond_37 ;  
   wire mux_cond_38 ;  
   wire mux_cond_39 ;  
   wire mux_cond_40 ;  
   wire mux_cond_41 ;  
   wire mux_cond_42 ;  
   wire mux_cond_43 ;  
   wire mux_cond_44 ;  
   wire mux_cond_45 ;  
   wire mux_cond_46 ;  
   wire mux_cond_47 ;  
   wire mux_cond_48 ;  
   wire mux_cond_49 ;  
   wire mux_cond_50 ;  
   wire mux_cond_51 ;  
   wire mux_cond_52 ;  
   wire mux_cond_53 ;  
   wire mux_cond_54 ;  
   wire mux_cond_55 ;  
   wire mux_cond_56 ;  
   wire mux_cond_57 ;  
   wire mux_cond_58 ;  
   wire mux_cond_59 ;  
   wire mux_cond_60 ;  
   wire mux_cond_61 ;  
   wire mux_cond_62 ;  
   wire mux_cond_63 ;  
   wire mux_cond_64 ;  
   wire mux_cond_65 ;  
   wire mux_cond_66 ;  
   wire mux_cond_67 ;  
   wire mux_cond_68 ;  
   wire r_sectored_hit_shl ;  
   wire [19:0] r_sectored_hit_pad ;  
   wire [9:0] r_sectored_repl_addr_shl ;  
   wire [19:0] r_sectored_repl_addr_pad ;  
   wire [19:0] r_superpage_repl_addr_shl ;  
   wire [19:0] r_superpage_repl_addr_pad ;  
   wire [7:0] special_entry_valid_0_shl ;  
   wire [19:0] special_entry_valid_0_pad ;  
   wire [19:0] special_entry_level_shl ;  
   wire [19:0] special_entry_level_pad ;  
   wire [7:0] state_shl ;  
   wire [19:0] state_pad ;  
   wire [14:0] r_sectored_hit_addr_shl ;  
   wire [19:0] r_sectored_hit_addr_pad ;  
   wire [5:0] mux_cond_0_shl ;  
   wire [19:0] mux_cond_0_pad ;  
   wire [11:0] mux_cond_1_shl ;  
   wire [19:0] mux_cond_1_pad ;  
   wire [2:0] mux_cond_2_shl ;  
   wire [19:0] mux_cond_2_pad ;  
   wire [12:0] mux_cond_3_shl ;  
   wire [19:0] mux_cond_3_pad ;  
   wire [11:0] mux_cond_4_shl ;  
   wire [19:0] mux_cond_4_pad ;  
   wire [1:0] mux_cond_5_shl ;  
   wire [19:0] mux_cond_5_pad ;  
   wire [13:0] mux_cond_6_shl ;  
   wire [19:0] mux_cond_6_pad ;  
   wire [6:0] mux_cond_7_shl ;  
   wire [19:0] mux_cond_7_pad ;  
   wire [4:0] mux_cond_8_shl ;  
   wire [19:0] mux_cond_8_pad ;  
   wire [17:0] mux_cond_9_shl ;  
   wire [19:0] mux_cond_9_pad ;  
   wire [5:0] mux_cond_10_shl ;  
   wire [19:0] mux_cond_10_pad ;  
   wire [9:0] mux_cond_11_shl ;  
   wire [19:0] mux_cond_11_pad ;  
   wire [1:0] mux_cond_12_shl ;  
   wire [19:0] mux_cond_12_pad ;  
   wire [9:0] mux_cond_13_shl ;  
   wire [19:0] mux_cond_13_pad ;  
   wire [12:0] mux_cond_14_shl ;  
   wire [19:0] mux_cond_14_pad ;  
   wire [7:0] mux_cond_15_shl ;  
   wire [19:0] mux_cond_15_pad ;  
   wire [6:0] mux_cond_16_shl ;  
   wire [19:0] mux_cond_16_pad ;  
   wire [7:0] mux_cond_17_shl ;  
   wire [19:0] mux_cond_17_pad ;  
   wire [16:0] mux_cond_18_shl ;  
   wire [19:0] mux_cond_18_pad ;  
   wire [8:0] mux_cond_19_shl ;  
   wire [19:0] mux_cond_19_pad ;  
   wire [1:0] mux_cond_20_shl ;  
   wire [19:0] mux_cond_20_pad ;  
   wire [5:0] mux_cond_21_shl ;  
   wire [19:0] mux_cond_21_pad ;  
   wire [11:0] mux_cond_22_shl ;  
   wire [19:0] mux_cond_22_pad ;  
   wire [2:0] mux_cond_23_shl ;  
   wire [19:0] mux_cond_23_pad ;  
   wire [14:0] mux_cond_24_shl ;  
   wire [19:0] mux_cond_24_pad ;  
   wire [3:0] mux_cond_25_shl ;  
   wire [19:0] mux_cond_25_pad ;  
   wire [11:0] mux_cond_26_shl ;  
   wire [19:0] mux_cond_26_pad ;  
   wire mux_cond_27_shl ;  
   wire [19:0] mux_cond_27_pad ;  
   wire [18:0] mux_cond_28_shl ;  
   wire [19:0] mux_cond_28_pad ;  
   wire [14:0] mux_cond_29_shl ;  
   wire [19:0] mux_cond_29_pad ;  
   wire [8:0] mux_cond_30_shl ;  
   wire [19:0] mux_cond_30_pad ;  
   wire [3:0] mux_cond_31_shl ;  
   wire [19:0] mux_cond_31_pad ;  
   wire [2:0] mux_cond_32_shl ;  
   wire [19:0] mux_cond_32_pad ;  
   wire mux_cond_33_shl ;  
   wire [19:0] mux_cond_33_pad ;  
   wire [7:0] mux_cond_34_shl ;  
   wire [19:0] mux_cond_34_pad ;  
   wire [4:0] mux_cond_35_shl ;  
   wire [19:0] mux_cond_35_pad ;  
   wire [3:0] mux_cond_36_shl ;  
   wire [19:0] mux_cond_36_pad ;  
   wire [4:0] mux_cond_37_shl ;  
   wire [19:0] mux_cond_37_pad ;  
   wire [12:0] mux_cond_38_shl ;  
   wire [19:0] mux_cond_38_pad ;  
   wire [9:0] mux_cond_39_shl ;  
   wire [19:0] mux_cond_39_pad ;  
   wire mux_cond_40_shl ;  
   wire [19:0] mux_cond_40_pad ;  
   wire [16:0] mux_cond_41_shl ;  
   wire [19:0] mux_cond_41_pad ;  
   wire [4:0] mux_cond_42_shl ;  
   wire [19:0] mux_cond_42_pad ;  
   wire [18:0] mux_cond_43_shl ;  
   wire [19:0] mux_cond_43_pad ;  
   wire [8:0] mux_cond_44_shl ;  
   wire [19:0] mux_cond_44_pad ;  
   wire [17:0] mux_cond_45_shl ;  
   wire [19:0] mux_cond_45_pad ;  
   wire [5:0] mux_cond_46_shl ;  
   wire [19:0] mux_cond_46_pad ;  
   wire [8:0] mux_cond_47_shl ;  
   wire [19:0] mux_cond_47_pad ;  
   wire [7:0] mux_cond_48_shl ;  
   wire [19:0] mux_cond_48_pad ;  
   wire [16:0] mux_cond_49_shl ;  
   wire [19:0] mux_cond_49_pad ;  
   wire [8:0] mux_cond_50_shl ;  
   wire [19:0] mux_cond_50_pad ;  
   wire [4:0] mux_cond_51_shl ;  
   wire [19:0] mux_cond_51_pad ;  
   wire [3:0] mux_cond_52_shl ;  
   wire [19:0] mux_cond_52_pad ;  
   wire [6:0] mux_cond_53_shl ;  
   wire [19:0] mux_cond_53_pad ;  
   wire [18:0] mux_cond_54_shl ;  
   wire [19:0] mux_cond_54_pad ;  
   wire [15:0] mux_cond_55_shl ;  
   wire [19:0] mux_cond_55_pad ;  
   wire [16:0] mux_cond_56_shl ;  
   wire [19:0] mux_cond_56_pad ;  
   wire [7:0] mux_cond_57_shl ;  
   wire [19:0] mux_cond_57_pad ;  
   wire [11:0] mux_cond_58_shl ;  
   wire [19:0] mux_cond_58_pad ;  
   wire [14:0] mux_cond_59_shl ;  
   wire [19:0] mux_cond_59_pad ;  
   wire [13:0] mux_cond_60_shl ;  
   wire [19:0] mux_cond_60_pad ;  
   wire [8:0] mux_cond_61_shl ;  
   wire [19:0] mux_cond_61_pad ;  
   wire [7:0] mux_cond_62_shl ;  
   wire [19:0] mux_cond_62_pad ;  
   wire [6:0] mux_cond_63_shl ;  
   wire [19:0] mux_cond_63_pad ;  
   wire [19:0] mux_cond_64_shl ;  
   wire [19:0] mux_cond_64_pad ;  
   wire [11:0] mux_cond_65_shl ;  
   wire [19:0] mux_cond_65_pad ;  
   wire [6:0] mux_cond_66_shl ;  
   wire [19:0] mux_cond_66_pad ;  
   wire [10:0] mux_cond_67_shl ;  
   wire [19:0] mux_cond_67_pad ;  
   wire [13:0] mux_cond_68_shl ;  
   wire [19:0] mux_cond_68_pad ;  
   wire [16:0] sectored_entries_0_0_valid_3_shl ;  
   wire [19:0] sectored_entries_0_0_valid_3_pad ;  
   wire [8:0] sectored_entries_0_0_valid_2_shl ;  
   wire [19:0] sectored_entries_0_0_valid_2_pad ;  
   wire [8:0] sectored_entries_0_2_valid_0_shl ;  
   wire [19:0] sectored_entries_0_2_valid_0_pad ;  
   wire [8:0] sectored_entries_0_3_valid_0_shl ;  
   wire [19:0] sectored_entries_0_3_valid_0_pad ;  
   wire [1:0] superpage_entries_2_level_shl ;  
   wire [19:0] superpage_entries_2_level_pad ;  
   wire sectored_entries_0_7_valid_1_shl ;  
   wire [19:0] sectored_entries_0_7_valid_1_pad ;  
   wire [8:0] sectored_entries_0_4_valid_0_shl ;  
   wire [19:0] sectored_entries_0_4_valid_0_pad ;  
   wire [16:0] sectored_entries_0_1_valid_3_shl ;  
   wire [19:0] sectored_entries_0_1_valid_3_pad ;  
   wire sectored_entries_0_1_valid_1_shl ;  
   wire [19:0] sectored_entries_0_1_valid_1_pad ;  
   wire [16:0] sectored_entries_0_2_valid_3_shl ;  
   wire [19:0] sectored_entries_0_2_valid_3_pad ;  
   wire sectored_entries_0_2_valid_1_shl ;  
   wire [19:0] sectored_entries_0_2_valid_1_pad ;  
   wire [11:0] superpage_entries_1_valid_0_shl ;  
   wire [19:0] superpage_entries_1_valid_0_pad ;  
   wire [8:0] sectored_entries_0_7_valid_0_shl ;  
   wire [19:0] sectored_entries_0_7_valid_0_pad ;  
   wire [11:0] superpage_entries_3_valid_0_shl ;  
   wire [19:0] superpage_entries_3_valid_0_pad ;  
   wire [16:0] sectored_entries_0_5_valid_3_shl ;  
   wire [19:0] sectored_entries_0_5_valid_3_pad ;  
   wire sectored_entries_0_5_valid_1_shl ;  
   wire [19:0] sectored_entries_0_5_valid_1_pad ;  
   wire [16:0] sectored_entries_0_4_valid_3_shl ;  
   wire [19:0] sectored_entries_0_4_valid_3_pad ;  
   wire [8:0] sectored_entries_0_5_valid_2_shl ;  
   wire [19:0] sectored_entries_0_5_valid_2_pad ;  
   wire [8:0] sectored_entries_0_1_valid_2_shl ;  
   wire [19:0] sectored_entries_0_1_valid_2_pad ;  
   wire sectored_entries_0_3_valid_1_shl ;  
   wire [19:0] sectored_entries_0_3_valid_1_pad ;  
   wire [8:0] sectored_entries_0_1_valid_0_shl ;  
   wire [19:0] sectored_entries_0_1_valid_0_pad ;  
   wire [8:0] sectored_entries_0_4_valid_2_shl ;  
   wire [19:0] sectored_entries_0_4_valid_2_pad ;  
   wire sectored_entries_0_4_valid_1_shl ;  
   wire [19:0] sectored_entries_0_4_valid_1_pad ;  
   wire [1:0] superpage_entries_3_level_shl ;  
   wire [19:0] superpage_entries_3_level_pad ;  
   wire sectored_entries_0_0_valid_1_shl ;  
   wire [19:0] sectored_entries_0_0_valid_1_pad ;  
   wire [8:0] sectored_entries_0_3_valid_2_shl ;  
   wire [19:0] sectored_entries_0_3_valid_2_pad ;  
   wire sectored_entries_0_6_valid_1_shl ;  
   wire [19:0] sectored_entries_0_6_valid_1_pad ;  
   wire [16:0] sectored_entries_0_7_valid_3_shl ;  
   wire [19:0] sectored_entries_0_7_valid_3_pad ;  
   wire [16:0] sectored_entries_0_3_valid_3_shl ;  
   wire [19:0] sectored_entries_0_3_valid_3_pad ;  
   wire [8:0] sectored_entries_0_0_valid_0_shl ;  
   wire [19:0] sectored_entries_0_0_valid_0_pad ;  
   wire [11:0] superpage_entries_0_valid_0_shl ;  
   wire [19:0] superpage_entries_0_valid_0_pad ;  
   wire [8:0] sectored_entries_0_2_valid_2_shl ;  
   wire [19:0] sectored_entries_0_2_valid_2_pad ;  
   wire [8:0] sectored_entries_0_6_valid_2_shl ;  
   wire [19:0] sectored_entries_0_6_valid_2_pad ;  
   wire [11:0] superpage_entries_2_valid_0_shl ;  
   wire [19:0] superpage_entries_2_valid_0_pad ;  
   wire [16:0] sectored_entries_0_6_valid_3_shl ;  
   wire [19:0] sectored_entries_0_6_valid_3_pad ;  
   wire [8:0] sectored_entries_0_6_valid_0_shl ;  
   wire [19:0] sectored_entries_0_6_valid_0_pad ;  
   wire [8:0] sectored_entries_0_7_valid_2_shl ;  
   wire [19:0] sectored_entries_0_7_valid_2_pad ;  
   wire [1:0] superpage_entries_0_level_shl ;  
   wire [19:0] superpage_entries_0_level_pad ;  
   wire [1:0] superpage_entries_1_level_shl ;  
   wire [19:0] superpage_entries_1_level_pad ;  
   wire [8:0] sectored_entries_0_5_valid_0_shl ;  
   wire [19:0] sectored_entries_0_5_valid_0_pad ;  
   wire [19:0] TLB_xor64 ;  
   wire [19:0] TLB_xor31 ;  
   wire [19:0] TLB_xor65 ;  
   wire [19:0] TLB_xor66 ;  
   wire [19:0] TLB_xor32 ;  
   wire [19:0] TLB_xor15 ;  
   wire [19:0] TLB_xor68 ;  
   wire [19:0] TLB_xor33 ;  
   wire [19:0] TLB_xor69 ;  
   wire [19:0] TLB_xor70 ;  
   wire [19:0] TLB_xor34 ;  
   wire [19:0] TLB_xor16 ;  
   wire [19:0] TLB_xor7 ;  
   wire [19:0] TLB_xor72 ;  
   wire [19:0] TLB_xor35 ;  
   wire [19:0] TLB_xor73 ;  
   wire [19:0] TLB_xor74 ;  
   wire [19:0] TLB_xor36 ;  
   wire [19:0] TLB_xor17 ;  
   wire [19:0] TLB_xor75 ;  
   wire [19:0] TLB_xor76 ;  
   wire [19:0] TLB_xor37 ;  
   wire [19:0] TLB_xor77 ;  
   wire [19:0] TLB_xor78 ;  
   wire [19:0] TLB_xor38 ;  
   wire [19:0] TLB_xor18 ;  
   wire [19:0] TLB_xor8 ;  
   wire [19:0] TLB_xor3 ;  
   wire [19:0] TLB_xor80 ;  
   wire [19:0] TLB_xor39 ;  
   wire [19:0] TLB_xor81 ;  
   wire [19:0] TLB_xor82 ;  
   wire [19:0] TLB_xor40 ;  
   wire [19:0] TLB_xor19 ;  
   wire [19:0] TLB_xor84 ;  
   wire [19:0] TLB_xor41 ;  
   wire [19:0] TLB_xor85 ;  
   wire [19:0] TLB_xor86 ;  
   wire [19:0] TLB_xor42 ;  
   wire [19:0] TLB_xor20 ;  
   wire [19:0] TLB_xor9 ;  
   wire [19:0] TLB_xor88 ;  
   wire [19:0] TLB_xor43 ;  
   wire [19:0] TLB_xor89 ;  
   wire [19:0] TLB_xor90 ;  
   wire [19:0] TLB_xor44 ;  
   wire [19:0] TLB_xor21 ;  
   wire [19:0] TLB_xor91 ;  
   wire [19:0] TLB_xor92 ;  
   wire [19:0] TLB_xor45 ;  
   wire [19:0] TLB_xor93 ;  
   wire [19:0] TLB_xor94 ;  
   wire [19:0] TLB_xor46 ;  
   wire [19:0] TLB_xor22 ;  
   wire [19:0] TLB_xor10 ;  
   wire [19:0] TLB_xor4 ;  
   wire [19:0] TLB_xor1 ;  
   wire [19:0] TLB_xor96 ;  
   wire [19:0] TLB_xor47 ;  
   wire [19:0] TLB_xor97 ;  
   wire [19:0] TLB_xor98 ;  
   wire [19:0] TLB_xor48 ;  
   wire [19:0] TLB_xor23 ;  
   wire [19:0] TLB_xor100 ;  
   wire [19:0] TLB_xor49 ;  
   wire [19:0] TLB_xor101 ;  
   wire [19:0] TLB_xor102 ;  
   wire [19:0] TLB_xor50 ;  
   wire [19:0] TLB_xor24 ;  
   wire [19:0] TLB_xor11 ;  
   wire [19:0] TLB_xor104 ;  
   wire [19:0] TLB_xor51 ;  
   wire [19:0] TLB_xor105 ;  
   wire [19:0] TLB_xor106 ;  
   wire [19:0] TLB_xor52 ;  
   wire [19:0] TLB_xor25 ;  
   wire [19:0] TLB_xor107 ;  
   wire [19:0] TLB_xor108 ;  
   wire [19:0] TLB_xor53 ;  
   wire [19:0] TLB_xor109 ;  
   wire [19:0] TLB_xor110 ;  
   wire [19:0] TLB_xor54 ;  
   wire [19:0] TLB_xor26 ;  
   wire [19:0] TLB_xor12 ;  
   wire [19:0] TLB_xor5 ;  
   wire [19:0] TLB_xor112 ;  
   wire [19:0] TLB_xor55 ;  
   wire [19:0] TLB_xor113 ;  
   wire [19:0] TLB_xor114 ;  
   wire [19:0] TLB_xor56 ;  
   wire [19:0] TLB_xor27 ;  
   wire [19:0] TLB_xor116 ;  
   wire [19:0] TLB_xor57 ;  
   wire [19:0] TLB_xor117 ;  
   wire [19:0] TLB_xor118 ;  
   wire [19:0] TLB_xor58 ;  
   wire [19:0] TLB_xor28 ;  
   wire [19:0] TLB_xor13 ;  
   wire [19:0] TLB_xor120 ;  
   wire [19:0] TLB_xor59 ;  
   wire [19:0] TLB_xor121 ;  
   wire [19:0] TLB_xor122 ;  
   wire [19:0] TLB_xor60 ;  
   wire [19:0] TLB_xor29 ;  
   wire [19:0] TLB_xor123 ;  
   wire [19:0] TLB_xor124 ;  
   wire [19:0] TLB_xor61 ;  
   wire [19:0] TLB_xor125 ;  
   wire [19:0] TLB_xor126 ;  
   wire [19:0] TLB_xor62 ;  
   wire [19:0] TLB_xor30 ;  
   wire [19:0] TLB_xor14 ;  
   wire [19:0] TLB_xor6 ;  
   wire [19:0] TLB_xor2 ;  
   wire [19:0] TLB_xor0 ;  
   wire [29:0] mpu_ppn_barrier_sum ;  
   wire [29:0] entries_barrier_10_sum ;  
   wire [29:0] entries_barrier_9_sum ;  
   wire [29:0] entries_barrier_7_sum ;  
   wire [29:0] entries_barrier_sum ;  
   wire [29:0] entries_barrier_6_sum ;  
   wire [29:0] entries_barrier_12_sum ;  
   wire [29:0] entries_barrier_1_sum ;  
   wire [29:0] entries_barrier_11_sum ;  
   wire [29:0] entries_barrier_8_sum ;  
   wire [29:0] pmp_sum ;  
   wire [29:0] entries_barrier_2_sum ;  
   wire [29:0] entries_barrier_4_sum ;  
   wire [29:0] entries_barrier_5_sum ;  
   wire [29:0] entries_barrier_3_sum ;  
   wire stopEn0 ;  
   wire entries_barrier_11_metaAssert_wire ;  
   wire entries_barrier_8_metaAssert_wire ;  
   wire entries_barrier_3_metaAssert_wire ;  
   wire pmp_metaAssert_wire ;  
   wire entries_barrier_6_metaAssert_wire ;  
   wire entries_barrier_12_metaAssert_wire ;  
   wire entries_barrier_9_metaAssert_wire ;  
   wire mpu_ppn_barrier_metaAssert_wire ;  
   wire entries_barrier_7_metaAssert_wire ;  
   wire entries_barrier_metaAssert_wire ;  
   wire entries_barrier_5_metaAssert_wire ;  
   wire entries_barrier_2_metaAssert_wire ;  
   wire entries_barrier_4_metaAssert_wire ;  
   wire entries_barrier_1_metaAssert_wire ;  
   wire entries_barrier_10_metaAssert_wire ;  
   wire TLB_or7 ;  
   wire TLB_or8 ;  
   wire TLB_or3 ;  
   wire TLB_or9 ;  
   wire TLB_or10 ;  
   wire TLB_or4 ;  
   wire TLB_or1 ;  
   wire TLB_or11 ;  
   wire TLB_or12 ;  
   wire TLB_or5 ;  
   wire TLB_or13 ;  
   wire TLB_or14 ;  
   wire TLB_or6 ;  
   wire TLB_or2 ;  
   wire TLB_or0 ;  
   reg TLB_metaAssert ;  
   reg [31:0] _RAND_103 ;  
  OptimizationBarrier mpu_ppn_barrier(.io_x_ppn(mpu_ppn_barrier_io_x_ppn),.io_x_u(mpu_ppn_barrier_io_x_u),.io_x_ae(mpu_ppn_barrier_io_x_ae),.io_x_sw(mpu_ppn_barrier_io_x_sw),.io_x_sx(mpu_ppn_barrier_io_x_sx),.io_x_sr(mpu_ppn_barrier_io_x_sr),.io_x_pw(mpu_ppn_barrier_io_x_pw),.io_x_px(mpu_ppn_barrier_io_x_px),.io_x_pr(mpu_ppn_barrier_io_x_pr),.io_x_ppp(mpu_ppn_barrier_io_x_ppp),.io_x_pal(mpu_ppn_barrier_io_x_pal),.io_x_paa(mpu_ppn_barrier_io_x_paa),.io_x_eff(mpu_ppn_barrier_io_x_eff),.io_x_c(mpu_ppn_barrier_io_x_c),.io_y_ppn(mpu_ppn_barrier_io_y_ppn),.io_y_u(mpu_ppn_barrier_io_y_u),.io_y_ae(mpu_ppn_barrier_io_y_ae),.io_y_sw(mpu_ppn_barrier_io_y_sw),.io_y_sx(mpu_ppn_barrier_io_y_sx),.io_y_sr(mpu_ppn_barrier_io_y_sr),.io_y_pw(mpu_ppn_barrier_io_y_pw),.io_y_px(mpu_ppn_barrier_io_y_px),.io_y_pr(mpu_ppn_barrier_io_y_pr),.io_y_ppp(mpu_ppn_barrier_io_y_ppp),.io_y_pal(mpu_ppn_barrier_io_y_pal),.io_y_paa(mpu_ppn_barrier_io_y_paa),.io_y_eff(mpu_ppn_barrier_io_y_eff),.io_y_c(mpu_ppn_barrier_io_y_c),.io_covSum(mpu_ppn_barrier_io_covSum),.metaAssert(mpu_ppn_barrier_metaAssert)); 
  PMPChecker pmp(.io_prv(pmp_io_prv),.io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),.io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),.io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),.io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),.io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),.io_pmp_0_addr(pmp_io_pmp_0_addr),.io_pmp_0_mask(pmp_io_pmp_0_mask),.io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),.io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),.io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),.io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),.io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),.io_pmp_1_addr(pmp_io_pmp_1_addr),.io_pmp_1_mask(pmp_io_pmp_1_mask),.io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),.io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),.io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),.io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),.io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),.io_pmp_2_addr(pmp_io_pmp_2_addr),.io_pmp_2_mask(pmp_io_pmp_2_mask),.io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),.io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),.io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),.io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),.io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),.io_pmp_3_addr(pmp_io_pmp_3_addr),.io_pmp_3_mask(pmp_io_pmp_3_mask),.io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),.io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),.io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),.io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),.io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),.io_pmp_4_addr(pmp_io_pmp_4_addr),.io_pmp_4_mask(pmp_io_pmp_4_mask),.io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),.io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),.io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),.io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),.io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),.io_pmp_5_addr(pmp_io_pmp_5_addr),.io_pmp_5_mask(pmp_io_pmp_5_mask),.io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),.io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),.io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),.io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),.io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),.io_pmp_6_addr(pmp_io_pmp_6_addr),.io_pmp_6_mask(pmp_io_pmp_6_mask),.io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),.io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),.io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),.io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),.io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),.io_pmp_7_addr(pmp_io_pmp_7_addr),.io_pmp_7_mask(pmp_io_pmp_7_mask),.io_addr(pmp_io_addr),.io_size(pmp_io_size),.io_r(pmp_io_r),.io_w(pmp_io_w),.io_x(pmp_io_x),.io_covSum(pmp_io_covSum),.metaAssert(pmp_metaAssert)); 
  OptimizationBarrier entries_barrier(.io_x_ppn(entries_barrier_io_x_ppn),.io_x_u(entries_barrier_io_x_u),.io_x_ae(entries_barrier_io_x_ae),.io_x_sw(entries_barrier_io_x_sw),.io_x_sx(entries_barrier_io_x_sx),.io_x_sr(entries_barrier_io_x_sr),.io_x_pw(entries_barrier_io_x_pw),.io_x_px(entries_barrier_io_x_px),.io_x_pr(entries_barrier_io_x_pr),.io_x_ppp(entries_barrier_io_x_ppp),.io_x_pal(entries_barrier_io_x_pal),.io_x_paa(entries_barrier_io_x_paa),.io_x_eff(entries_barrier_io_x_eff),.io_x_c(entries_barrier_io_x_c),.io_y_ppn(entries_barrier_io_y_ppn),.io_y_u(entries_barrier_io_y_u),.io_y_ae(entries_barrier_io_y_ae),.io_y_sw(entries_barrier_io_y_sw),.io_y_sx(entries_barrier_io_y_sx),.io_y_sr(entries_barrier_io_y_sr),.io_y_pw(entries_barrier_io_y_pw),.io_y_px(entries_barrier_io_y_px),.io_y_pr(entries_barrier_io_y_pr),.io_y_ppp(entries_barrier_io_y_ppp),.io_y_pal(entries_barrier_io_y_pal),.io_y_paa(entries_barrier_io_y_paa),.io_y_eff(entries_barrier_io_y_eff),.io_y_c(entries_barrier_io_y_c),.io_covSum(entries_barrier_io_covSum),.metaAssert(entries_barrier_metaAssert)); 
  OptimizationBarrier entries_barrier_1(.io_x_ppn(entries_barrier_1_io_x_ppn),.io_x_u(entries_barrier_1_io_x_u),.io_x_ae(entries_barrier_1_io_x_ae),.io_x_sw(entries_barrier_1_io_x_sw),.io_x_sx(entries_barrier_1_io_x_sx),.io_x_sr(entries_barrier_1_io_x_sr),.io_x_pw(entries_barrier_1_io_x_pw),.io_x_px(entries_barrier_1_io_x_px),.io_x_pr(entries_barrier_1_io_x_pr),.io_x_ppp(entries_barrier_1_io_x_ppp),.io_x_pal(entries_barrier_1_io_x_pal),.io_x_paa(entries_barrier_1_io_x_paa),.io_x_eff(entries_barrier_1_io_x_eff),.io_x_c(entries_barrier_1_io_x_c),.io_y_ppn(entries_barrier_1_io_y_ppn),.io_y_u(entries_barrier_1_io_y_u),.io_y_ae(entries_barrier_1_io_y_ae),.io_y_sw(entries_barrier_1_io_y_sw),.io_y_sx(entries_barrier_1_io_y_sx),.io_y_sr(entries_barrier_1_io_y_sr),.io_y_pw(entries_barrier_1_io_y_pw),.io_y_px(entries_barrier_1_io_y_px),.io_y_pr(entries_barrier_1_io_y_pr),.io_y_ppp(entries_barrier_1_io_y_ppp),.io_y_pal(entries_barrier_1_io_y_pal),.io_y_paa(entries_barrier_1_io_y_paa),.io_y_eff(entries_barrier_1_io_y_eff),.io_y_c(entries_barrier_1_io_y_c),.io_covSum(entries_barrier_1_io_covSum),.metaAssert(entries_barrier_1_metaAssert)); 
  OptimizationBarrier entries_barrier_2(.io_x_ppn(entries_barrier_2_io_x_ppn),.io_x_u(entries_barrier_2_io_x_u),.io_x_ae(entries_barrier_2_io_x_ae),.io_x_sw(entries_barrier_2_io_x_sw),.io_x_sx(entries_barrier_2_io_x_sx),.io_x_sr(entries_barrier_2_io_x_sr),.io_x_pw(entries_barrier_2_io_x_pw),.io_x_px(entries_barrier_2_io_x_px),.io_x_pr(entries_barrier_2_io_x_pr),.io_x_ppp(entries_barrier_2_io_x_ppp),.io_x_pal(entries_barrier_2_io_x_pal),.io_x_paa(entries_barrier_2_io_x_paa),.io_x_eff(entries_barrier_2_io_x_eff),.io_x_c(entries_barrier_2_io_x_c),.io_y_ppn(entries_barrier_2_io_y_ppn),.io_y_u(entries_barrier_2_io_y_u),.io_y_ae(entries_barrier_2_io_y_ae),.io_y_sw(entries_barrier_2_io_y_sw),.io_y_sx(entries_barrier_2_io_y_sx),.io_y_sr(entries_barrier_2_io_y_sr),.io_y_pw(entries_barrier_2_io_y_pw),.io_y_px(entries_barrier_2_io_y_px),.io_y_pr(entries_barrier_2_io_y_pr),.io_y_ppp(entries_barrier_2_io_y_ppp),.io_y_pal(entries_barrier_2_io_y_pal),.io_y_paa(entries_barrier_2_io_y_paa),.io_y_eff(entries_barrier_2_io_y_eff),.io_y_c(entries_barrier_2_io_y_c),.io_covSum(entries_barrier_2_io_covSum),.metaAssert(entries_barrier_2_metaAssert)); 
  OptimizationBarrier entries_barrier_3(.io_x_ppn(entries_barrier_3_io_x_ppn),.io_x_u(entries_barrier_3_io_x_u),.io_x_ae(entries_barrier_3_io_x_ae),.io_x_sw(entries_barrier_3_io_x_sw),.io_x_sx(entries_barrier_3_io_x_sx),.io_x_sr(entries_barrier_3_io_x_sr),.io_x_pw(entries_barrier_3_io_x_pw),.io_x_px(entries_barrier_3_io_x_px),.io_x_pr(entries_barrier_3_io_x_pr),.io_x_ppp(entries_barrier_3_io_x_ppp),.io_x_pal(entries_barrier_3_io_x_pal),.io_x_paa(entries_barrier_3_io_x_paa),.io_x_eff(entries_barrier_3_io_x_eff),.io_x_c(entries_barrier_3_io_x_c),.io_y_ppn(entries_barrier_3_io_y_ppn),.io_y_u(entries_barrier_3_io_y_u),.io_y_ae(entries_barrier_3_io_y_ae),.io_y_sw(entries_barrier_3_io_y_sw),.io_y_sx(entries_barrier_3_io_y_sx),.io_y_sr(entries_barrier_3_io_y_sr),.io_y_pw(entries_barrier_3_io_y_pw),.io_y_px(entries_barrier_3_io_y_px),.io_y_pr(entries_barrier_3_io_y_pr),.io_y_ppp(entries_barrier_3_io_y_ppp),.io_y_pal(entries_barrier_3_io_y_pal),.io_y_paa(entries_barrier_3_io_y_paa),.io_y_eff(entries_barrier_3_io_y_eff),.io_y_c(entries_barrier_3_io_y_c),.io_covSum(entries_barrier_3_io_covSum),.metaAssert(entries_barrier_3_metaAssert)); 
  OptimizationBarrier entries_barrier_4(.io_x_ppn(entries_barrier_4_io_x_ppn),.io_x_u(entries_barrier_4_io_x_u),.io_x_ae(entries_barrier_4_io_x_ae),.io_x_sw(entries_barrier_4_io_x_sw),.io_x_sx(entries_barrier_4_io_x_sx),.io_x_sr(entries_barrier_4_io_x_sr),.io_x_pw(entries_barrier_4_io_x_pw),.io_x_px(entries_barrier_4_io_x_px),.io_x_pr(entries_barrier_4_io_x_pr),.io_x_ppp(entries_barrier_4_io_x_ppp),.io_x_pal(entries_barrier_4_io_x_pal),.io_x_paa(entries_barrier_4_io_x_paa),.io_x_eff(entries_barrier_4_io_x_eff),.io_x_c(entries_barrier_4_io_x_c),.io_y_ppn(entries_barrier_4_io_y_ppn),.io_y_u(entries_barrier_4_io_y_u),.io_y_ae(entries_barrier_4_io_y_ae),.io_y_sw(entries_barrier_4_io_y_sw),.io_y_sx(entries_barrier_4_io_y_sx),.io_y_sr(entries_barrier_4_io_y_sr),.io_y_pw(entries_barrier_4_io_y_pw),.io_y_px(entries_barrier_4_io_y_px),.io_y_pr(entries_barrier_4_io_y_pr),.io_y_ppp(entries_barrier_4_io_y_ppp),.io_y_pal(entries_barrier_4_io_y_pal),.io_y_paa(entries_barrier_4_io_y_paa),.io_y_eff(entries_barrier_4_io_y_eff),.io_y_c(entries_barrier_4_io_y_c),.io_covSum(entries_barrier_4_io_covSum),.metaAssert(entries_barrier_4_metaAssert)); 
  OptimizationBarrier entries_barrier_5(.io_x_ppn(entries_barrier_5_io_x_ppn),.io_x_u(entries_barrier_5_io_x_u),.io_x_ae(entries_barrier_5_io_x_ae),.io_x_sw(entries_barrier_5_io_x_sw),.io_x_sx(entries_barrier_5_io_x_sx),.io_x_sr(entries_barrier_5_io_x_sr),.io_x_pw(entries_barrier_5_io_x_pw),.io_x_px(entries_barrier_5_io_x_px),.io_x_pr(entries_barrier_5_io_x_pr),.io_x_ppp(entries_barrier_5_io_x_ppp),.io_x_pal(entries_barrier_5_io_x_pal),.io_x_paa(entries_barrier_5_io_x_paa),.io_x_eff(entries_barrier_5_io_x_eff),.io_x_c(entries_barrier_5_io_x_c),.io_y_ppn(entries_barrier_5_io_y_ppn),.io_y_u(entries_barrier_5_io_y_u),.io_y_ae(entries_barrier_5_io_y_ae),.io_y_sw(entries_barrier_5_io_y_sw),.io_y_sx(entries_barrier_5_io_y_sx),.io_y_sr(entries_barrier_5_io_y_sr),.io_y_pw(entries_barrier_5_io_y_pw),.io_y_px(entries_barrier_5_io_y_px),.io_y_pr(entries_barrier_5_io_y_pr),.io_y_ppp(entries_barrier_5_io_y_ppp),.io_y_pal(entries_barrier_5_io_y_pal),.io_y_paa(entries_barrier_5_io_y_paa),.io_y_eff(entries_barrier_5_io_y_eff),.io_y_c(entries_barrier_5_io_y_c),.io_covSum(entries_barrier_5_io_covSum),.metaAssert(entries_barrier_5_metaAssert)); 
  OptimizationBarrier entries_barrier_6(.io_x_ppn(entries_barrier_6_io_x_ppn),.io_x_u(entries_barrier_6_io_x_u),.io_x_ae(entries_barrier_6_io_x_ae),.io_x_sw(entries_barrier_6_io_x_sw),.io_x_sx(entries_barrier_6_io_x_sx),.io_x_sr(entries_barrier_6_io_x_sr),.io_x_pw(entries_barrier_6_io_x_pw),.io_x_px(entries_barrier_6_io_x_px),.io_x_pr(entries_barrier_6_io_x_pr),.io_x_ppp(entries_barrier_6_io_x_ppp),.io_x_pal(entries_barrier_6_io_x_pal),.io_x_paa(entries_barrier_6_io_x_paa),.io_x_eff(entries_barrier_6_io_x_eff),.io_x_c(entries_barrier_6_io_x_c),.io_y_ppn(entries_barrier_6_io_y_ppn),.io_y_u(entries_barrier_6_io_y_u),.io_y_ae(entries_barrier_6_io_y_ae),.io_y_sw(entries_barrier_6_io_y_sw),.io_y_sx(entries_barrier_6_io_y_sx),.io_y_sr(entries_barrier_6_io_y_sr),.io_y_pw(entries_barrier_6_io_y_pw),.io_y_px(entries_barrier_6_io_y_px),.io_y_pr(entries_barrier_6_io_y_pr),.io_y_ppp(entries_barrier_6_io_y_ppp),.io_y_pal(entries_barrier_6_io_y_pal),.io_y_paa(entries_barrier_6_io_y_paa),.io_y_eff(entries_barrier_6_io_y_eff),.io_y_c(entries_barrier_6_io_y_c),.io_covSum(entries_barrier_6_io_covSum),.metaAssert(entries_barrier_6_metaAssert)); 
  OptimizationBarrier entries_barrier_7(.io_x_ppn(entries_barrier_7_io_x_ppn),.io_x_u(entries_barrier_7_io_x_u),.io_x_ae(entries_barrier_7_io_x_ae),.io_x_sw(entries_barrier_7_io_x_sw),.io_x_sx(entries_barrier_7_io_x_sx),.io_x_sr(entries_barrier_7_io_x_sr),.io_x_pw(entries_barrier_7_io_x_pw),.io_x_px(entries_barrier_7_io_x_px),.io_x_pr(entries_barrier_7_io_x_pr),.io_x_ppp(entries_barrier_7_io_x_ppp),.io_x_pal(entries_barrier_7_io_x_pal),.io_x_paa(entries_barrier_7_io_x_paa),.io_x_eff(entries_barrier_7_io_x_eff),.io_x_c(entries_barrier_7_io_x_c),.io_y_ppn(entries_barrier_7_io_y_ppn),.io_y_u(entries_barrier_7_io_y_u),.io_y_ae(entries_barrier_7_io_y_ae),.io_y_sw(entries_barrier_7_io_y_sw),.io_y_sx(entries_barrier_7_io_y_sx),.io_y_sr(entries_barrier_7_io_y_sr),.io_y_pw(entries_barrier_7_io_y_pw),.io_y_px(entries_barrier_7_io_y_px),.io_y_pr(entries_barrier_7_io_y_pr),.io_y_ppp(entries_barrier_7_io_y_ppp),.io_y_pal(entries_barrier_7_io_y_pal),.io_y_paa(entries_barrier_7_io_y_paa),.io_y_eff(entries_barrier_7_io_y_eff),.io_y_c(entries_barrier_7_io_y_c),.io_covSum(entries_barrier_7_io_covSum),.metaAssert(entries_barrier_7_metaAssert)); 
  OptimizationBarrier entries_barrier_8(.io_x_ppn(entries_barrier_8_io_x_ppn),.io_x_u(entries_barrier_8_io_x_u),.io_x_ae(entries_barrier_8_io_x_ae),.io_x_sw(entries_barrier_8_io_x_sw),.io_x_sx(entries_barrier_8_io_x_sx),.io_x_sr(entries_barrier_8_io_x_sr),.io_x_pw(entries_barrier_8_io_x_pw),.io_x_px(entries_barrier_8_io_x_px),.io_x_pr(entries_barrier_8_io_x_pr),.io_x_ppp(entries_barrier_8_io_x_ppp),.io_x_pal(entries_barrier_8_io_x_pal),.io_x_paa(entries_barrier_8_io_x_paa),.io_x_eff(entries_barrier_8_io_x_eff),.io_x_c(entries_barrier_8_io_x_c),.io_y_ppn(entries_barrier_8_io_y_ppn),.io_y_u(entries_barrier_8_io_y_u),.io_y_ae(entries_barrier_8_io_y_ae),.io_y_sw(entries_barrier_8_io_y_sw),.io_y_sx(entries_barrier_8_io_y_sx),.io_y_sr(entries_barrier_8_io_y_sr),.io_y_pw(entries_barrier_8_io_y_pw),.io_y_px(entries_barrier_8_io_y_px),.io_y_pr(entries_barrier_8_io_y_pr),.io_y_ppp(entries_barrier_8_io_y_ppp),.io_y_pal(entries_barrier_8_io_y_pal),.io_y_paa(entries_barrier_8_io_y_paa),.io_y_eff(entries_barrier_8_io_y_eff),.io_y_c(entries_barrier_8_io_y_c),.io_covSum(entries_barrier_8_io_covSum),.metaAssert(entries_barrier_8_metaAssert)); 
  OptimizationBarrier entries_barrier_9(.io_x_ppn(entries_barrier_9_io_x_ppn),.io_x_u(entries_barrier_9_io_x_u),.io_x_ae(entries_barrier_9_io_x_ae),.io_x_sw(entries_barrier_9_io_x_sw),.io_x_sx(entries_barrier_9_io_x_sx),.io_x_sr(entries_barrier_9_io_x_sr),.io_x_pw(entries_barrier_9_io_x_pw),.io_x_px(entries_barrier_9_io_x_px),.io_x_pr(entries_barrier_9_io_x_pr),.io_x_ppp(entries_barrier_9_io_x_ppp),.io_x_pal(entries_barrier_9_io_x_pal),.io_x_paa(entries_barrier_9_io_x_paa),.io_x_eff(entries_barrier_9_io_x_eff),.io_x_c(entries_barrier_9_io_x_c),.io_y_ppn(entries_barrier_9_io_y_ppn),.io_y_u(entries_barrier_9_io_y_u),.io_y_ae(entries_barrier_9_io_y_ae),.io_y_sw(entries_barrier_9_io_y_sw),.io_y_sx(entries_barrier_9_io_y_sx),.io_y_sr(entries_barrier_9_io_y_sr),.io_y_pw(entries_barrier_9_io_y_pw),.io_y_px(entries_barrier_9_io_y_px),.io_y_pr(entries_barrier_9_io_y_pr),.io_y_ppp(entries_barrier_9_io_y_ppp),.io_y_pal(entries_barrier_9_io_y_pal),.io_y_paa(entries_barrier_9_io_y_paa),.io_y_eff(entries_barrier_9_io_y_eff),.io_y_c(entries_barrier_9_io_y_c),.io_covSum(entries_barrier_9_io_covSum),.metaAssert(entries_barrier_9_metaAssert)); 
  OptimizationBarrier entries_barrier_10(.io_x_ppn(entries_barrier_10_io_x_ppn),.io_x_u(entries_barrier_10_io_x_u),.io_x_ae(entries_barrier_10_io_x_ae),.io_x_sw(entries_barrier_10_io_x_sw),.io_x_sx(entries_barrier_10_io_x_sx),.io_x_sr(entries_barrier_10_io_x_sr),.io_x_pw(entries_barrier_10_io_x_pw),.io_x_px(entries_barrier_10_io_x_px),.io_x_pr(entries_barrier_10_io_x_pr),.io_x_ppp(entries_barrier_10_io_x_ppp),.io_x_pal(entries_barrier_10_io_x_pal),.io_x_paa(entries_barrier_10_io_x_paa),.io_x_eff(entries_barrier_10_io_x_eff),.io_x_c(entries_barrier_10_io_x_c),.io_y_ppn(entries_barrier_10_io_y_ppn),.io_y_u(entries_barrier_10_io_y_u),.io_y_ae(entries_barrier_10_io_y_ae),.io_y_sw(entries_barrier_10_io_y_sw),.io_y_sx(entries_barrier_10_io_y_sx),.io_y_sr(entries_barrier_10_io_y_sr),.io_y_pw(entries_barrier_10_io_y_pw),.io_y_px(entries_barrier_10_io_y_px),.io_y_pr(entries_barrier_10_io_y_pr),.io_y_ppp(entries_barrier_10_io_y_ppp),.io_y_pal(entries_barrier_10_io_y_pal),.io_y_paa(entries_barrier_10_io_y_paa),.io_y_eff(entries_barrier_10_io_y_eff),.io_y_c(entries_barrier_10_io_y_c),.io_covSum(entries_barrier_10_io_covSum),.metaAssert(entries_barrier_10_metaAssert)); 
  OptimizationBarrier entries_barrier_11(.io_x_ppn(entries_barrier_11_io_x_ppn),.io_x_u(entries_barrier_11_io_x_u),.io_x_ae(entries_barrier_11_io_x_ae),.io_x_sw(entries_barrier_11_io_x_sw),.io_x_sx(entries_barrier_11_io_x_sx),.io_x_sr(entries_barrier_11_io_x_sr),.io_x_pw(entries_barrier_11_io_x_pw),.io_x_px(entries_barrier_11_io_x_px),.io_x_pr(entries_barrier_11_io_x_pr),.io_x_ppp(entries_barrier_11_io_x_ppp),.io_x_pal(entries_barrier_11_io_x_pal),.io_x_paa(entries_barrier_11_io_x_paa),.io_x_eff(entries_barrier_11_io_x_eff),.io_x_c(entries_barrier_11_io_x_c),.io_y_ppn(entries_barrier_11_io_y_ppn),.io_y_u(entries_barrier_11_io_y_u),.io_y_ae(entries_barrier_11_io_y_ae),.io_y_sw(entries_barrier_11_io_y_sw),.io_y_sx(entries_barrier_11_io_y_sx),.io_y_sr(entries_barrier_11_io_y_sr),.io_y_pw(entries_barrier_11_io_y_pw),.io_y_px(entries_barrier_11_io_y_px),.io_y_pr(entries_barrier_11_io_y_pr),.io_y_ppp(entries_barrier_11_io_y_ppp),.io_y_pal(entries_barrier_11_io_y_pal),.io_y_paa(entries_barrier_11_io_y_paa),.io_y_eff(entries_barrier_11_io_y_eff),.io_y_c(entries_barrier_11_io_y_c),.io_covSum(entries_barrier_11_io_covSum),.metaAssert(entries_barrier_11_metaAssert)); 
  OptimizationBarrier entries_barrier_12(.io_x_ppn(entries_barrier_12_io_x_ppn),.io_x_u(entries_barrier_12_io_x_u),.io_x_ae(entries_barrier_12_io_x_ae),.io_x_sw(entries_barrier_12_io_x_sw),.io_x_sx(entries_barrier_12_io_x_sx),.io_x_sr(entries_barrier_12_io_x_sr),.io_x_pw(entries_barrier_12_io_x_pw),.io_x_px(entries_barrier_12_io_x_px),.io_x_pr(entries_barrier_12_io_x_pr),.io_x_ppp(entries_barrier_12_io_x_ppp),.io_x_pal(entries_barrier_12_io_x_pal),.io_x_paa(entries_barrier_12_io_x_paa),.io_x_eff(entries_barrier_12_io_x_eff),.io_x_c(entries_barrier_12_io_x_c),.io_y_ppn(entries_barrier_12_io_y_ppn),.io_y_u(entries_barrier_12_io_y_u),.io_y_ae(entries_barrier_12_io_y_ae),.io_y_sw(entries_barrier_12_io_y_sw),.io_y_sx(entries_barrier_12_io_y_sx),.io_y_sr(entries_barrier_12_io_y_sr),.io_y_pw(entries_barrier_12_io_y_pw),.io_y_px(entries_barrier_12_io_y_px),.io_y_pr(entries_barrier_12_io_y_pr),.io_y_ppp(entries_barrier_12_io_y_ppp),.io_y_pal(entries_barrier_12_io_y_pal),.io_y_paa(entries_barrier_12_io_y_paa),.io_y_eff(entries_barrier_12_io_y_eff),.io_y_c(entries_barrier_12_io_y_c),.io_covSum(entries_barrier_12_io_covSum),.metaAssert(entries_barrier_12_metaAssert)); 
  assign vpn=io_req_bits_vaddr[38:12]; 
  assign priv_s=io_ptw_status_dprv[0]; 
  assign priv_uses_vm=io_ptw_status_dprv<=2'h1; 
  assign _vm_enabled_T_2=io_ptw_ptbr_mode[3]&priv_uses_vm; 
  assign vm_enabled=_vm_enabled_T_2&~io_req_bits_passthrough; 
  assign refill_ppn=io_ptw_resp_bits_pte_ppn[19:0]; 
  assign _invalidate_refill_T=state==2'h1; 
  assign _invalidate_refill_T_1=state==2'h3; 
  assign _invalidate_refill_T_2=_invalidate_refill_T|_invalidate_refill_T_1; 
  assign invalidate_refill=_invalidate_refill_T_2|io_sfence_valid; 
  assign mpu_ppn_hi=mpu_ppn_barrier_io_y_ppn[19:18]; 
  assign mpu_ppn_ignore=special_entry_level<2'h1; 
  assign _mpu_ppn_T_17=mpu_ppn_ignore ? vpn:27'h0; 
  assign _GEN_919={7'b0,mpu_ppn_barrier_io_y_ppn}; 
  assign _mpu_ppn_T_18=_mpu_ppn_T_17|_GEN_919; 
  assign mpu_ppn_lo=_mpu_ppn_T_18[17:9]; 
  assign mpu_ppn_ignore_1=special_entry_level<2'h2; 
  assign _mpu_ppn_T_19=mpu_ppn_ignore_1 ? vpn:27'h0; 
  assign _mpu_ppn_T_20=_mpu_ppn_T_19|_GEN_919; 
  assign mpu_ppn_lo_1=_mpu_ppn_T_20[8:0]; 
  assign _mpu_ppn_T_21={mpu_ppn_hi,mpu_ppn_lo,mpu_ppn_lo_1}; 
  assign _mpu_ppn_T_23=vm_enabled ? {8'b0,_mpu_ppn_T_21}:io_req_bits_vaddr[39:12]; 
  assign mpu_ppn=io_ptw_resp_valid ? {8'b0,refill_ppn}:_mpu_ppn_T_23; 
  assign mpu_physaddr_lo=io_req_bits_vaddr[11:0]; 
  assign mpu_physaddr={mpu_ppn,mpu_physaddr_lo}; 
  assign _mpu_priv_T=io_ptw_resp_valid|io_req_bits_passthrough; 
  assign _mpu_priv_T_2={io_ptw_status_debug,io_ptw_status_dprv}; 
  assign mpu_priv=_mpu_priv_T ? 3'h1:_mpu_priv_T_2; 
  assign _legal_address_T=mpu_physaddr^40'h3000; 
  assign _legal_address_T_1={1'b0,$signed(_legal_address_T)}; 
  assign _legal_address_T_3=$signed(_legal_address_T_1)&-41'sh1000; 
  assign _legal_address_T_4=$signed(_legal_address_T_3)==41'sh0; 
  assign _legal_address_T_5=mpu_physaddr^40'hc000000; 
  assign _legal_address_T_6={1'b0,$signed(_legal_address_T_5)}; 
  assign _legal_address_T_8=$signed(_legal_address_T_6)&-41'sh4000000; 
  assign _legal_address_T_9=$signed(_legal_address_T_8)==41'sh0; 
  assign _legal_address_T_10=mpu_physaddr^40'h2000000; 
  assign _legal_address_T_11={1'b0,$signed(_legal_address_T_10)}; 
  assign _legal_address_T_13=$signed(_legal_address_T_11)&-41'sh10000; 
  assign _legal_address_T_14=$signed(_legal_address_T_13)==41'sh0; 
  assign _legal_address_T_16={1'b0,$signed(mpu_physaddr)}; 
  assign _legal_address_T_18=$signed(_legal_address_T_16)&-41'sh1000; 
  assign _legal_address_T_19=$signed(_legal_address_T_18)==41'sh0; 
  assign _legal_address_T_20=mpu_physaddr^40'h10000; 
  assign _legal_address_T_21={1'b0,$signed(_legal_address_T_20)}; 
  assign _legal_address_T_23=$signed(_legal_address_T_21)&-41'sh10000; 
  assign _legal_address_T_24=$signed(_legal_address_T_23)==41'sh0; 
  assign _legal_address_T_25=mpu_physaddr^40'h80000000; 
  assign _legal_address_T_26={1'b0,$signed(_legal_address_T_25)}; 
  assign _legal_address_T_28=$signed(_legal_address_T_26)&-41'sh10000000; 
  assign _legal_address_T_29=$signed(_legal_address_T_28)==41'sh0; 
  assign _legal_address_T_30=mpu_physaddr^40'h60000000; 
  assign _legal_address_T_31={1'b0,$signed(_legal_address_T_30)}; 
  assign _legal_address_T_33=$signed(_legal_address_T_31)&-41'sh20000000; 
  assign _legal_address_T_34=$signed(_legal_address_T_33)==41'sh0; 
  assign _legal_address_T_35=_legal_address_T_4|_legal_address_T_9; 
  assign _legal_address_T_36=_legal_address_T_35|_legal_address_T_14; 
  assign _legal_address_T_37=_legal_address_T_36|_legal_address_T_19; 
  assign _legal_address_T_38=_legal_address_T_37|_legal_address_T_24; 
  assign _legal_address_T_39=_legal_address_T_38|_legal_address_T_29; 
  assign legal_address=_legal_address_T_39|_legal_address_T_34; 
  assign _cacheable_T_8=$signed(_legal_address_T_26)&41'sh80000000; 
  assign _cacheable_T_9=$signed(_cacheable_T_8)==41'sh0; 
  assign cacheable=legal_address&_cacheable_T_9; 
  assign _homogeneous_T_54=mpu_physaddr^40'h8000000; 
  assign _homogeneous_T_55={1'b0,$signed(_homogeneous_T_54)}; 
  assign _homogeneous_T_57=$signed(_homogeneous_T_55)&41'shc8000000; 
  assign _homogeneous_T_58=$signed(_homogeneous_T_57)==41'sh0; 
  assign _homogeneous_T_71=$signed(_legal_address_T_16)&41'shc8010000; 
  assign _homogeneous_T_72=$signed(_homogeneous_T_71)==41'sh0; 
  assign _homogeneous_T_79=_homogeneous_T_72|_homogeneous_T_58; 
  assign _deny_access_to_debug_T=mpu_priv<=3'h3; 
  assign deny_access_to_debug=_deny_access_to_debug_T&_legal_address_T_19; 
  assign _prot_r_T_7=legal_address&~deny_access_to_debug; 
  assign prot_r=_prot_r_T_7&pmp_io_r; 
  assign _prot_w_T_10=mpu_physaddr^40'h40000000; 
  assign _prot_w_T_11={1'b0,$signed(_prot_w_T_10)}; 
  assign _prot_w_T_13=$signed(_prot_w_T_11)&41'shc0000000; 
  assign _prot_w_T_14=$signed(_prot_w_T_13)==41'sh0; 
  assign _prot_w_T_18=$signed(_legal_address_T_26)&41'shc0000000; 
  assign _prot_w_T_19=$signed(_prot_w_T_18)==41'sh0; 
  assign _prot_w_T_21=_homogeneous_T_79|_prot_w_T_14; 
  assign _prot_w_T_22=_prot_w_T_21|_prot_w_T_19; 
  assign _prot_w_T_31=legal_address&_prot_w_T_22; 
  assign _prot_w_T_33=_prot_w_T_31&~deny_access_to_debug; 
  assign prot_w=_prot_w_T_33&pmp_io_w; 
  assign prot_al=legal_address&_homogeneous_T_79; 
  assign _prot_x_T_3=$signed(_legal_address_T_16)&41'shca000000; 
  assign _prot_x_T_4=$signed(_prot_x_T_3)==41'sh0; 
  assign _prot_x_T_15=_prot_x_T_4|_prot_w_T_14; 
  assign _prot_x_T_16=_prot_x_T_15|_prot_w_T_19; 
  assign _prot_x_T_31=legal_address&_prot_x_T_16; 
  assign _prot_x_T_33=_prot_x_T_31&~deny_access_to_debug; 
  assign prot_x=_prot_x_T_33&pmp_io_x; 
  assign _prot_eff_T_20=$signed(_legal_address_T_16)&41'shca012000; 
  assign _prot_eff_T_21=$signed(_prot_eff_T_20)==41'sh0; 
  assign _prot_eff_T_25=$signed(_legal_address_T_11)&41'shca010000; 
  assign _prot_eff_T_26=$signed(_prot_eff_T_25)==41'sh0; 
  assign _prot_eff_T_37=_prot_eff_T_21|_prot_eff_T_26; 
  assign _prot_eff_T_38=_prot_eff_T_37|_homogeneous_T_58; 
  assign _prot_eff_T_39=_prot_eff_T_38|_prot_w_T_14; 
  assign prot_eff=legal_address&_prot_eff_T_39; 
  assign _sector_hits_T=sectored_entries_0_0_valid_0|sectored_entries_0_0_valid_1; 
  assign _sector_hits_T_1=_sector_hits_T|sectored_entries_0_0_valid_2; 
  assign _sector_hits_T_2=_sector_hits_T_1|sectored_entries_0_0_valid_3; 
  assign _sector_hits_T_3=sectored_entries_0_0_tag^vpn; 
  assign _sector_hits_T_5=_sector_hits_T_3[26:2]==25'h0; 
  assign sector_hits_0=_sector_hits_T_2&_sector_hits_T_5; 
  assign _sector_hits_T_6=sectored_entries_0_1_valid_0|sectored_entries_0_1_valid_1; 
  assign _sector_hits_T_7=_sector_hits_T_6|sectored_entries_0_1_valid_2; 
  assign _sector_hits_T_8=_sector_hits_T_7|sectored_entries_0_1_valid_3; 
  assign _sector_hits_T_9=sectored_entries_0_1_tag^vpn; 
  assign _sector_hits_T_11=_sector_hits_T_9[26:2]==25'h0; 
  assign sector_hits_1=_sector_hits_T_8&_sector_hits_T_11; 
  assign _sector_hits_T_12=sectored_entries_0_2_valid_0|sectored_entries_0_2_valid_1; 
  assign _sector_hits_T_13=_sector_hits_T_12|sectored_entries_0_2_valid_2; 
  assign _sector_hits_T_14=_sector_hits_T_13|sectored_entries_0_2_valid_3; 
  assign _sector_hits_T_15=sectored_entries_0_2_tag^vpn; 
  assign _sector_hits_T_17=_sector_hits_T_15[26:2]==25'h0; 
  assign sector_hits_2=_sector_hits_T_14&_sector_hits_T_17; 
  assign _sector_hits_T_18=sectored_entries_0_3_valid_0|sectored_entries_0_3_valid_1; 
  assign _sector_hits_T_19=_sector_hits_T_18|sectored_entries_0_3_valid_2; 
  assign _sector_hits_T_20=_sector_hits_T_19|sectored_entries_0_3_valid_3; 
  assign _sector_hits_T_21=sectored_entries_0_3_tag^vpn; 
  assign _sector_hits_T_23=_sector_hits_T_21[26:2]==25'h0; 
  assign sector_hits_3=_sector_hits_T_20&_sector_hits_T_23; 
  assign _sector_hits_T_24=sectored_entries_0_4_valid_0|sectored_entries_0_4_valid_1; 
  assign _sector_hits_T_25=_sector_hits_T_24|sectored_entries_0_4_valid_2; 
  assign _sector_hits_T_26=_sector_hits_T_25|sectored_entries_0_4_valid_3; 
  assign _sector_hits_T_27=sectored_entries_0_4_tag^vpn; 
  assign _sector_hits_T_29=_sector_hits_T_27[26:2]==25'h0; 
  assign sector_hits_4=_sector_hits_T_26&_sector_hits_T_29; 
  assign _sector_hits_T_30=sectored_entries_0_5_valid_0|sectored_entries_0_5_valid_1; 
  assign _sector_hits_T_31=_sector_hits_T_30|sectored_entries_0_5_valid_2; 
  assign _sector_hits_T_32=_sector_hits_T_31|sectored_entries_0_5_valid_3; 
  assign _sector_hits_T_33=sectored_entries_0_5_tag^vpn; 
  assign _sector_hits_T_35=_sector_hits_T_33[26:2]==25'h0; 
  assign sector_hits_5=_sector_hits_T_32&_sector_hits_T_35; 
  assign _sector_hits_T_36=sectored_entries_0_6_valid_0|sectored_entries_0_6_valid_1; 
  assign _sector_hits_T_37=_sector_hits_T_36|sectored_entries_0_6_valid_2; 
  assign _sector_hits_T_38=_sector_hits_T_37|sectored_entries_0_6_valid_3; 
  assign _sector_hits_T_39=sectored_entries_0_6_tag^vpn; 
  assign _sector_hits_T_41=_sector_hits_T_39[26:2]==25'h0; 
  assign sector_hits_6=_sector_hits_T_38&_sector_hits_T_41; 
  assign _sector_hits_T_42=sectored_entries_0_7_valid_0|sectored_entries_0_7_valid_1; 
  assign _sector_hits_T_43=_sector_hits_T_42|sectored_entries_0_7_valid_2; 
  assign _sector_hits_T_44=_sector_hits_T_43|sectored_entries_0_7_valid_3; 
  assign _sector_hits_T_45=sectored_entries_0_7_tag^vpn; 
  assign _sector_hits_T_47=_sector_hits_T_45[26:2]==25'h0; 
  assign sector_hits_7=_sector_hits_T_44&_sector_hits_T_47; 
  assign _superpage_hits_T_2=superpage_entries_0_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_4=superpage_entries_0_valid_0&_superpage_hits_T_2; 
  assign superpage_hits_ignore_1=superpage_entries_0_level<2'h1; 
  assign _superpage_hits_T_7=superpage_entries_0_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_8=superpage_hits_ignore_1|_superpage_hits_T_7; 
  assign superpage_hits_0=_superpage_hits_T_4&_superpage_hits_T_8; 
  assign _superpage_hits_T_16=superpage_entries_1_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_18=superpage_entries_1_valid_0&_superpage_hits_T_16; 
  assign superpage_hits_ignore_4=superpage_entries_1_level<2'h1; 
  assign _superpage_hits_T_21=superpage_entries_1_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_22=superpage_hits_ignore_4|_superpage_hits_T_21; 
  assign superpage_hits_1=_superpage_hits_T_18&_superpage_hits_T_22; 
  assign _superpage_hits_T_30=superpage_entries_2_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_32=superpage_entries_2_valid_0&_superpage_hits_T_30; 
  assign superpage_hits_ignore_7=superpage_entries_2_level<2'h1; 
  assign _superpage_hits_T_35=superpage_entries_2_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_36=superpage_hits_ignore_7|_superpage_hits_T_35; 
  assign superpage_hits_2=_superpage_hits_T_32&_superpage_hits_T_36; 
  assign _superpage_hits_T_44=superpage_entries_3_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_46=superpage_entries_3_valid_0&_superpage_hits_T_44; 
  assign superpage_hits_ignore_10=superpage_entries_3_level<2'h1; 
  assign _superpage_hits_T_49=superpage_entries_3_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_50=superpage_hits_ignore_10|_superpage_hits_T_49; 
  assign superpage_hits_3=_superpage_hits_T_46&_superpage_hits_T_50; 
  assign hitsVec_idx=vpn[1:0]; 
  assign _GEN_1=2'h1==hitsVec_idx ? sectored_entries_0_0_valid_1:sectored_entries_0_0_valid_0; 
  assign _GEN_2=2'h2==hitsVec_idx ? sectored_entries_0_0_valid_2:_GEN_1; 
  assign _GEN_3=2'h3==hitsVec_idx ? sectored_entries_0_0_valid_3:_GEN_2; 
  assign _hitsVec_T_3=_GEN_3&_sector_hits_T_5; 
  assign hitsVec_0=vm_enabled&_hitsVec_T_3; 
  assign _GEN_5=2'h1==hitsVec_idx ? sectored_entries_0_1_valid_1:sectored_entries_0_1_valid_0; 
  assign _GEN_6=2'h2==hitsVec_idx ? sectored_entries_0_1_valid_2:_GEN_5; 
  assign _GEN_7=2'h3==hitsVec_idx ? sectored_entries_0_1_valid_3:_GEN_6; 
  assign _hitsVec_T_7=_GEN_7&_sector_hits_T_11; 
  assign hitsVec_1=vm_enabled&_hitsVec_T_7; 
  assign _GEN_9=2'h1==hitsVec_idx ? sectored_entries_0_2_valid_1:sectored_entries_0_2_valid_0; 
  assign _GEN_10=2'h2==hitsVec_idx ? sectored_entries_0_2_valid_2:_GEN_9; 
  assign _GEN_11=2'h3==hitsVec_idx ? sectored_entries_0_2_valid_3:_GEN_10; 
  assign _hitsVec_T_11=_GEN_11&_sector_hits_T_17; 
  assign hitsVec_2=vm_enabled&_hitsVec_T_11; 
  assign _GEN_13=2'h1==hitsVec_idx ? sectored_entries_0_3_valid_1:sectored_entries_0_3_valid_0; 
  assign _GEN_14=2'h2==hitsVec_idx ? sectored_entries_0_3_valid_2:_GEN_13; 
  assign _GEN_15=2'h3==hitsVec_idx ? sectored_entries_0_3_valid_3:_GEN_14; 
  assign _hitsVec_T_15=_GEN_15&_sector_hits_T_23; 
  assign hitsVec_3=vm_enabled&_hitsVec_T_15; 
  assign _GEN_17=2'h1==hitsVec_idx ? sectored_entries_0_4_valid_1:sectored_entries_0_4_valid_0; 
  assign _GEN_18=2'h2==hitsVec_idx ? sectored_entries_0_4_valid_2:_GEN_17; 
  assign _GEN_19=2'h3==hitsVec_idx ? sectored_entries_0_4_valid_3:_GEN_18; 
  assign _hitsVec_T_19=_GEN_19&_sector_hits_T_29; 
  assign hitsVec_4=vm_enabled&_hitsVec_T_19; 
  assign _GEN_21=2'h1==hitsVec_idx ? sectored_entries_0_5_valid_1:sectored_entries_0_5_valid_0; 
  assign _GEN_22=2'h2==hitsVec_idx ? sectored_entries_0_5_valid_2:_GEN_21; 
  assign _GEN_23=2'h3==hitsVec_idx ? sectored_entries_0_5_valid_3:_GEN_22; 
  assign _hitsVec_T_23=_GEN_23&_sector_hits_T_35; 
  assign hitsVec_5=vm_enabled&_hitsVec_T_23; 
  assign _GEN_25=2'h1==hitsVec_idx ? sectored_entries_0_6_valid_1:sectored_entries_0_6_valid_0; 
  assign _GEN_26=2'h2==hitsVec_idx ? sectored_entries_0_6_valid_2:_GEN_25; 
  assign _GEN_27=2'h3==hitsVec_idx ? sectored_entries_0_6_valid_3:_GEN_26; 
  assign _hitsVec_T_27=_GEN_27&_sector_hits_T_41; 
  assign hitsVec_6=vm_enabled&_hitsVec_T_27; 
  assign _GEN_29=2'h1==hitsVec_idx ? sectored_entries_0_7_valid_1:sectored_entries_0_7_valid_0; 
  assign _GEN_30=2'h2==hitsVec_idx ? sectored_entries_0_7_valid_2:_GEN_29; 
  assign _GEN_31=2'h3==hitsVec_idx ? sectored_entries_0_7_valid_3:_GEN_30; 
  assign _hitsVec_T_31=_GEN_31&_sector_hits_T_47; 
  assign hitsVec_7=vm_enabled&_hitsVec_T_31; 
  assign hitsVec_8=vm_enabled&superpage_hits_0; 
  assign hitsVec_9=vm_enabled&superpage_hits_1; 
  assign hitsVec_10=vm_enabled&superpage_hits_2; 
  assign hitsVec_11=vm_enabled&superpage_hits_3; 
  assign _hitsVec_T_94=special_entry_tag[26:18]==vpn[26:18]; 
  assign _hitsVec_T_96=special_entry_valid_0&_hitsVec_T_94; 
  assign _hitsVec_T_99=special_entry_tag[17:9]==vpn[17:9]; 
  assign _hitsVec_T_100=mpu_ppn_ignore|_hitsVec_T_99; 
  assign _hitsVec_T_101=_hitsVec_T_96&_hitsVec_T_100; 
  assign _hitsVec_T_104=special_entry_tag[8:0]==vpn[8:0]; 
  assign _hitsVec_T_105=mpu_ppn_ignore_1|_hitsVec_T_104; 
  assign _hitsVec_T_106=_hitsVec_T_101&_hitsVec_T_105; 
  assign hitsVec_12=vm_enabled&_hitsVec_T_106; 
  assign real_hits_lo={hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; 
  assign real_hits={hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; 
  assign hits_hi=~vm_enabled; 
  assign hits={hits_hi,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; 
  assign newEntry_g=io_ptw_resp_bits_pte_g&io_ptw_resp_bits_pte_v; 
  assign _newEntry_sr_T_1=io_ptw_resp_bits_pte_x&~io_ptw_resp_bits_pte_w; 
  assign _newEntry_sr_T_2=io_ptw_resp_bits_pte_r|_newEntry_sr_T_1; 
  assign _newEntry_sr_T_3=io_ptw_resp_bits_pte_v&_newEntry_sr_T_2; 
  assign _newEntry_sr_T_4=_newEntry_sr_T_3&io_ptw_resp_bits_pte_a; 
  assign newEntry_sr=_newEntry_sr_T_4&io_ptw_resp_bits_pte_r; 
  assign _newEntry_sw_T_5=_newEntry_sr_T_4&io_ptw_resp_bits_pte_w; 
  assign newEntry_sw=_newEntry_sw_T_5&io_ptw_resp_bits_pte_d; 
  assign newEntry_sx=_newEntry_sr_T_4&io_ptw_resp_bits_pte_x; 
  assign special_entry_data_0_lo={prot_x,prot_r,_prot_w_T_31,prot_al,prot_al,prot_eff,cacheable,1'h0}; 
  assign _special_entry_data_0_T={refill_ppn,io_ptw_resp_bits_pte_u,newEntry_g,io_ptw_resp_bits_ae,newEntry_sw,newEntry_sx,newEntry_sr,prot_w,special_entry_data_0_lo}; 
  assign _GEN_32=invalidate_refill ? 1'h0:1'h1; 
  assign _T_2=io_ptw_resp_bits_level<2'h2; 
  assign _T_3=r_superpage_repl_addr==2'h0; 
  assign _GEN_35=_T_3 ? _GEN_32:superpage_entries_0_valid_0; 
  assign _T_4=r_superpage_repl_addr==2'h1; 
  assign _GEN_39=_T_4 ? _GEN_32:superpage_entries_1_valid_0; 
  assign _T_5=r_superpage_repl_addr==2'h2; 
  assign _GEN_43=_T_5 ? _GEN_32:superpage_entries_2_valid_0; 
  assign _T_6=r_superpage_repl_addr==2'h3; 
  assign _GEN_47=_T_6 ? _GEN_32:superpage_entries_3_valid_0; 
  assign waddr=r_sectored_hit ? r_sectored_hit_addr:r_sectored_repl_addr; 
  assign _T_7=waddr==3'h0; 
  assign _GEN_49=r_sectored_hit ? sectored_entries_0_0_valid_0:1'h0; 
  assign _GEN_50=r_sectored_hit ? sectored_entries_0_0_valid_1:1'h0; 
  assign _GEN_51=r_sectored_hit ? sectored_entries_0_0_valid_2:1'h0; 
  assign _GEN_52=r_sectored_hit ? sectored_entries_0_0_valid_3:1'h0; 
  assign idx=r_refill_tag[1:0]; 
  assign _GEN_921=2'h0==idx; 
  assign _GEN_53=_GEN_921|_GEN_49; 
  assign _GEN_922=2'h1==idx; 
  assign _GEN_54=_GEN_922|_GEN_50; 
  assign _GEN_923=2'h2==idx; 
  assign _GEN_55=_GEN_923|_GEN_51; 
  assign _GEN_924=2'h3==idx; 
  assign _GEN_56=_GEN_924|_GEN_52; 
  assign _GEN_61=invalidate_refill ? 1'h0:_GEN_53; 
  assign _GEN_62=invalidate_refill ? 1'h0:_GEN_54; 
  assign _GEN_63=invalidate_refill ? 1'h0:_GEN_55; 
  assign _GEN_64=invalidate_refill ? 1'h0:_GEN_56; 
  assign _GEN_65=_T_7 ? _GEN_61:sectored_entries_0_0_valid_0; 
  assign _GEN_66=_T_7 ? _GEN_62:sectored_entries_0_0_valid_1; 
  assign _GEN_67=_T_7 ? _GEN_63:sectored_entries_0_0_valid_2; 
  assign _GEN_68=_T_7 ? _GEN_64:sectored_entries_0_0_valid_3; 
  assign _T_9=waddr==3'h1; 
  assign _GEN_75=r_sectored_hit ? sectored_entries_0_1_valid_0:1'h0; 
  assign _GEN_76=r_sectored_hit ? sectored_entries_0_1_valid_1:1'h0; 
  assign _GEN_77=r_sectored_hit ? sectored_entries_0_1_valid_2:1'h0; 
  assign _GEN_78=r_sectored_hit ? sectored_entries_0_1_valid_3:1'h0; 
  assign _GEN_79=_GEN_921|_GEN_75; 
  assign _GEN_80=_GEN_922|_GEN_76; 
  assign _GEN_81=_GEN_923|_GEN_77; 
  assign _GEN_82=_GEN_924|_GEN_78; 
  assign _GEN_87=invalidate_refill ? 1'h0:_GEN_79; 
  assign _GEN_88=invalidate_refill ? 1'h0:_GEN_80; 
  assign _GEN_89=invalidate_refill ? 1'h0:_GEN_81; 
  assign _GEN_90=invalidate_refill ? 1'h0:_GEN_82; 
  assign _GEN_91=_T_9 ? _GEN_87:sectored_entries_0_1_valid_0; 
  assign _GEN_92=_T_9 ? _GEN_88:sectored_entries_0_1_valid_1; 
  assign _GEN_93=_T_9 ? _GEN_89:sectored_entries_0_1_valid_2; 
  assign _GEN_94=_T_9 ? _GEN_90:sectored_entries_0_1_valid_3; 
  assign _T_11=waddr==3'h2; 
  assign _GEN_101=r_sectored_hit ? sectored_entries_0_2_valid_0:1'h0; 
  assign _GEN_102=r_sectored_hit ? sectored_entries_0_2_valid_1:1'h0; 
  assign _GEN_103=r_sectored_hit ? sectored_entries_0_2_valid_2:1'h0; 
  assign _GEN_104=r_sectored_hit ? sectored_entries_0_2_valid_3:1'h0; 
  assign _GEN_105=_GEN_921|_GEN_101; 
  assign _GEN_106=_GEN_922|_GEN_102; 
  assign _GEN_107=_GEN_923|_GEN_103; 
  assign _GEN_108=_GEN_924|_GEN_104; 
  assign _GEN_113=invalidate_refill ? 1'h0:_GEN_105; 
  assign _GEN_114=invalidate_refill ? 1'h0:_GEN_106; 
  assign _GEN_115=invalidate_refill ? 1'h0:_GEN_107; 
  assign _GEN_116=invalidate_refill ? 1'h0:_GEN_108; 
  assign _GEN_117=_T_11 ? _GEN_113:sectored_entries_0_2_valid_0; 
  assign _GEN_118=_T_11 ? _GEN_114:sectored_entries_0_2_valid_1; 
  assign _GEN_119=_T_11 ? _GEN_115:sectored_entries_0_2_valid_2; 
  assign _GEN_120=_T_11 ? _GEN_116:sectored_entries_0_2_valid_3; 
  assign _T_13=waddr==3'h3; 
  assign _GEN_127=r_sectored_hit ? sectored_entries_0_3_valid_0:1'h0; 
  assign _GEN_128=r_sectored_hit ? sectored_entries_0_3_valid_1:1'h0; 
  assign _GEN_129=r_sectored_hit ? sectored_entries_0_3_valid_2:1'h0; 
  assign _GEN_130=r_sectored_hit ? sectored_entries_0_3_valid_3:1'h0; 
  assign _GEN_131=_GEN_921|_GEN_127; 
  assign _GEN_132=_GEN_922|_GEN_128; 
  assign _GEN_133=_GEN_923|_GEN_129; 
  assign _GEN_134=_GEN_924|_GEN_130; 
  assign _GEN_139=invalidate_refill ? 1'h0:_GEN_131; 
  assign _GEN_140=invalidate_refill ? 1'h0:_GEN_132; 
  assign _GEN_141=invalidate_refill ? 1'h0:_GEN_133; 
  assign _GEN_142=invalidate_refill ? 1'h0:_GEN_134; 
  assign _GEN_143=_T_13 ? _GEN_139:sectored_entries_0_3_valid_0; 
  assign _GEN_144=_T_13 ? _GEN_140:sectored_entries_0_3_valid_1; 
  assign _GEN_145=_T_13 ? _GEN_141:sectored_entries_0_3_valid_2; 
  assign _GEN_146=_T_13 ? _GEN_142:sectored_entries_0_3_valid_3; 
  assign _T_15=waddr==3'h4; 
  assign _GEN_153=r_sectored_hit ? sectored_entries_0_4_valid_0:1'h0; 
  assign _GEN_154=r_sectored_hit ? sectored_entries_0_4_valid_1:1'h0; 
  assign _GEN_155=r_sectored_hit ? sectored_entries_0_4_valid_2:1'h0; 
  assign _GEN_156=r_sectored_hit ? sectored_entries_0_4_valid_3:1'h0; 
  assign _GEN_157=_GEN_921|_GEN_153; 
  assign _GEN_158=_GEN_922|_GEN_154; 
  assign _GEN_159=_GEN_923|_GEN_155; 
  assign _GEN_160=_GEN_924|_GEN_156; 
  assign _GEN_165=invalidate_refill ? 1'h0:_GEN_157; 
  assign _GEN_166=invalidate_refill ? 1'h0:_GEN_158; 
  assign _GEN_167=invalidate_refill ? 1'h0:_GEN_159; 
  assign _GEN_168=invalidate_refill ? 1'h0:_GEN_160; 
  assign _GEN_169=_T_15 ? _GEN_165:sectored_entries_0_4_valid_0; 
  assign _GEN_170=_T_15 ? _GEN_166:sectored_entries_0_4_valid_1; 
  assign _GEN_171=_T_15 ? _GEN_167:sectored_entries_0_4_valid_2; 
  assign _GEN_172=_T_15 ? _GEN_168:sectored_entries_0_4_valid_3; 
  assign _T_17=waddr==3'h5; 
  assign _GEN_179=r_sectored_hit ? sectored_entries_0_5_valid_0:1'h0; 
  assign _GEN_180=r_sectored_hit ? sectored_entries_0_5_valid_1:1'h0; 
  assign _GEN_181=r_sectored_hit ? sectored_entries_0_5_valid_2:1'h0; 
  assign _GEN_182=r_sectored_hit ? sectored_entries_0_5_valid_3:1'h0; 
  assign _GEN_183=_GEN_921|_GEN_179; 
  assign _GEN_184=_GEN_922|_GEN_180; 
  assign _GEN_185=_GEN_923|_GEN_181; 
  assign _GEN_186=_GEN_924|_GEN_182; 
  assign _GEN_191=invalidate_refill ? 1'h0:_GEN_183; 
  assign _GEN_192=invalidate_refill ? 1'h0:_GEN_184; 
  assign _GEN_193=invalidate_refill ? 1'h0:_GEN_185; 
  assign _GEN_194=invalidate_refill ? 1'h0:_GEN_186; 
  assign _GEN_195=_T_17 ? _GEN_191:sectored_entries_0_5_valid_0; 
  assign _GEN_196=_T_17 ? _GEN_192:sectored_entries_0_5_valid_1; 
  assign _GEN_197=_T_17 ? _GEN_193:sectored_entries_0_5_valid_2; 
  assign _GEN_198=_T_17 ? _GEN_194:sectored_entries_0_5_valid_3; 
  assign _T_19=waddr==3'h6; 
  assign _GEN_205=r_sectored_hit ? sectored_entries_0_6_valid_0:1'h0; 
  assign _GEN_206=r_sectored_hit ? sectored_entries_0_6_valid_1:1'h0; 
  assign _GEN_207=r_sectored_hit ? sectored_entries_0_6_valid_2:1'h0; 
  assign _GEN_208=r_sectored_hit ? sectored_entries_0_6_valid_3:1'h0; 
  assign _GEN_209=_GEN_921|_GEN_205; 
  assign _GEN_210=_GEN_922|_GEN_206; 
  assign _GEN_211=_GEN_923|_GEN_207; 
  assign _GEN_212=_GEN_924|_GEN_208; 
  assign _GEN_217=invalidate_refill ? 1'h0:_GEN_209; 
  assign _GEN_218=invalidate_refill ? 1'h0:_GEN_210; 
  assign _GEN_219=invalidate_refill ? 1'h0:_GEN_211; 
  assign _GEN_220=invalidate_refill ? 1'h0:_GEN_212; 
  assign _GEN_221=_T_19 ? _GEN_217:sectored_entries_0_6_valid_0; 
  assign _GEN_222=_T_19 ? _GEN_218:sectored_entries_0_6_valid_1; 
  assign _GEN_223=_T_19 ? _GEN_219:sectored_entries_0_6_valid_2; 
  assign _GEN_224=_T_19 ? _GEN_220:sectored_entries_0_6_valid_3; 
  assign _T_21=waddr==3'h7; 
  assign _GEN_231=r_sectored_hit ? sectored_entries_0_7_valid_0:1'h0; 
  assign _GEN_232=r_sectored_hit ? sectored_entries_0_7_valid_1:1'h0; 
  assign _GEN_233=r_sectored_hit ? sectored_entries_0_7_valid_2:1'h0; 
  assign _GEN_234=r_sectored_hit ? sectored_entries_0_7_valid_3:1'h0; 
  assign _GEN_235=_GEN_921|_GEN_231; 
  assign _GEN_236=_GEN_922|_GEN_232; 
  assign _GEN_237=_GEN_923|_GEN_233; 
  assign _GEN_238=_GEN_924|_GEN_234; 
  assign _GEN_243=invalidate_refill ? 1'h0:_GEN_235; 
  assign _GEN_244=invalidate_refill ? 1'h0:_GEN_236; 
  assign _GEN_245=invalidate_refill ? 1'h0:_GEN_237; 
  assign _GEN_246=invalidate_refill ? 1'h0:_GEN_238; 
  assign _GEN_247=_T_21 ? _GEN_243:sectored_entries_0_7_valid_0; 
  assign _GEN_248=_T_21 ? _GEN_244:sectored_entries_0_7_valid_1; 
  assign _GEN_249=_T_21 ? _GEN_245:sectored_entries_0_7_valid_2; 
  assign _GEN_250=_T_21 ? _GEN_246:sectored_entries_0_7_valid_3; 
  assign _GEN_259=_T_2 ? _GEN_35:superpage_entries_0_valid_0; 
  assign _GEN_263=_T_2 ? _GEN_39:superpage_entries_1_valid_0; 
  assign _GEN_267=_T_2 ? _GEN_43:superpage_entries_2_valid_0; 
  assign _GEN_271=_T_2 ? _GEN_47:superpage_entries_3_valid_0; 
  assign _GEN_273=_T_2 ? sectored_entries_0_0_valid_0:_GEN_65; 
  assign _GEN_274=_T_2 ? sectored_entries_0_0_valid_1:_GEN_66; 
  assign _GEN_275=_T_2 ? sectored_entries_0_0_valid_2:_GEN_67; 
  assign _GEN_276=_T_2 ? sectored_entries_0_0_valid_3:_GEN_68; 
  assign _GEN_283=_T_2 ? sectored_entries_0_1_valid_0:_GEN_91; 
  assign _GEN_284=_T_2 ? sectored_entries_0_1_valid_1:_GEN_92; 
  assign _GEN_285=_T_2 ? sectored_entries_0_1_valid_2:_GEN_93; 
  assign _GEN_286=_T_2 ? sectored_entries_0_1_valid_3:_GEN_94; 
  assign _GEN_293=_T_2 ? sectored_entries_0_2_valid_0:_GEN_117; 
  assign _GEN_294=_T_2 ? sectored_entries_0_2_valid_1:_GEN_118; 
  assign _GEN_295=_T_2 ? sectored_entries_0_2_valid_2:_GEN_119; 
  assign _GEN_296=_T_2 ? sectored_entries_0_2_valid_3:_GEN_120; 
  assign _GEN_303=_T_2 ? sectored_entries_0_3_valid_0:_GEN_143; 
  assign _GEN_304=_T_2 ? sectored_entries_0_3_valid_1:_GEN_144; 
  assign _GEN_305=_T_2 ? sectored_entries_0_3_valid_2:_GEN_145; 
  assign _GEN_306=_T_2 ? sectored_entries_0_3_valid_3:_GEN_146; 
  assign _GEN_313=_T_2 ? sectored_entries_0_4_valid_0:_GEN_169; 
  assign _GEN_314=_T_2 ? sectored_entries_0_4_valid_1:_GEN_170; 
  assign _GEN_315=_T_2 ? sectored_entries_0_4_valid_2:_GEN_171; 
  assign _GEN_316=_T_2 ? sectored_entries_0_4_valid_3:_GEN_172; 
  assign _GEN_323=_T_2 ? sectored_entries_0_5_valid_0:_GEN_195; 
  assign _GEN_324=_T_2 ? sectored_entries_0_5_valid_1:_GEN_196; 
  assign _GEN_325=_T_2 ? sectored_entries_0_5_valid_2:_GEN_197; 
  assign _GEN_326=_T_2 ? sectored_entries_0_5_valid_3:_GEN_198; 
  assign _GEN_333=_T_2 ? sectored_entries_0_6_valid_0:_GEN_221; 
  assign _GEN_334=_T_2 ? sectored_entries_0_6_valid_1:_GEN_222; 
  assign _GEN_335=_T_2 ? sectored_entries_0_6_valid_2:_GEN_223; 
  assign _GEN_336=_T_2 ? sectored_entries_0_6_valid_3:_GEN_224; 
  assign _GEN_343=_T_2 ? sectored_entries_0_7_valid_0:_GEN_247; 
  assign _GEN_344=_T_2 ? sectored_entries_0_7_valid_1:_GEN_248; 
  assign _GEN_345=_T_2 ? sectored_entries_0_7_valid_2:_GEN_249; 
  assign _GEN_346=_T_2 ? sectored_entries_0_7_valid_3:_GEN_250; 
  assign _GEN_355=io_ptw_resp_bits_homogeneous ? special_entry_valid_0:_GEN_32; 
  assign _GEN_359=io_ptw_resp_bits_homogeneous ? _GEN_259:superpage_entries_0_valid_0; 
  assign _GEN_363=io_ptw_resp_bits_homogeneous ? _GEN_263:superpage_entries_1_valid_0; 
  assign _GEN_367=io_ptw_resp_bits_homogeneous ? _GEN_267:superpage_entries_2_valid_0; 
  assign _GEN_371=io_ptw_resp_bits_homogeneous ? _GEN_271:superpage_entries_3_valid_0; 
  assign _GEN_373=io_ptw_resp_bits_homogeneous ? _GEN_273:sectored_entries_0_0_valid_0; 
  assign _GEN_374=io_ptw_resp_bits_homogeneous ? _GEN_274:sectored_entries_0_0_valid_1; 
  assign _GEN_375=io_ptw_resp_bits_homogeneous ? _GEN_275:sectored_entries_0_0_valid_2; 
  assign _GEN_376=io_ptw_resp_bits_homogeneous ? _GEN_276:sectored_entries_0_0_valid_3; 
  assign _GEN_383=io_ptw_resp_bits_homogeneous ? _GEN_283:sectored_entries_0_1_valid_0; 
  assign _GEN_384=io_ptw_resp_bits_homogeneous ? _GEN_284:sectored_entries_0_1_valid_1; 
  assign _GEN_385=io_ptw_resp_bits_homogeneous ? _GEN_285:sectored_entries_0_1_valid_2; 
  assign _GEN_386=io_ptw_resp_bits_homogeneous ? _GEN_286:sectored_entries_0_1_valid_3; 
  assign _GEN_393=io_ptw_resp_bits_homogeneous ? _GEN_293:sectored_entries_0_2_valid_0; 
  assign _GEN_394=io_ptw_resp_bits_homogeneous ? _GEN_294:sectored_entries_0_2_valid_1; 
  assign _GEN_395=io_ptw_resp_bits_homogeneous ? _GEN_295:sectored_entries_0_2_valid_2; 
  assign _GEN_396=io_ptw_resp_bits_homogeneous ? _GEN_296:sectored_entries_0_2_valid_3; 
  assign _GEN_403=io_ptw_resp_bits_homogeneous ? _GEN_303:sectored_entries_0_3_valid_0; 
  assign _GEN_404=io_ptw_resp_bits_homogeneous ? _GEN_304:sectored_entries_0_3_valid_1; 
  assign _GEN_405=io_ptw_resp_bits_homogeneous ? _GEN_305:sectored_entries_0_3_valid_2; 
  assign _GEN_406=io_ptw_resp_bits_homogeneous ? _GEN_306:sectored_entries_0_3_valid_3; 
  assign _GEN_413=io_ptw_resp_bits_homogeneous ? _GEN_313:sectored_entries_0_4_valid_0; 
  assign _GEN_414=io_ptw_resp_bits_homogeneous ? _GEN_314:sectored_entries_0_4_valid_1; 
  assign _GEN_415=io_ptw_resp_bits_homogeneous ? _GEN_315:sectored_entries_0_4_valid_2; 
  assign _GEN_416=io_ptw_resp_bits_homogeneous ? _GEN_316:sectored_entries_0_4_valid_3; 
  assign _GEN_423=io_ptw_resp_bits_homogeneous ? _GEN_323:sectored_entries_0_5_valid_0; 
  assign _GEN_424=io_ptw_resp_bits_homogeneous ? _GEN_324:sectored_entries_0_5_valid_1; 
  assign _GEN_425=io_ptw_resp_bits_homogeneous ? _GEN_325:sectored_entries_0_5_valid_2; 
  assign _GEN_426=io_ptw_resp_bits_homogeneous ? _GEN_326:sectored_entries_0_5_valid_3; 
  assign _GEN_433=io_ptw_resp_bits_homogeneous ? _GEN_333:sectored_entries_0_6_valid_0; 
  assign _GEN_434=io_ptw_resp_bits_homogeneous ? _GEN_334:sectored_entries_0_6_valid_1; 
  assign _GEN_435=io_ptw_resp_bits_homogeneous ? _GEN_335:sectored_entries_0_6_valid_2; 
  assign _GEN_436=io_ptw_resp_bits_homogeneous ? _GEN_336:sectored_entries_0_6_valid_3; 
  assign _GEN_443=io_ptw_resp_bits_homogeneous ? _GEN_343:sectored_entries_0_7_valid_0; 
  assign _GEN_444=io_ptw_resp_bits_homogeneous ? _GEN_344:sectored_entries_0_7_valid_1; 
  assign _GEN_445=io_ptw_resp_bits_homogeneous ? _GEN_345:sectored_entries_0_7_valid_2; 
  assign _GEN_446=io_ptw_resp_bits_homogeneous ? _GEN_346:sectored_entries_0_7_valid_3; 
  assign _GEN_455=io_ptw_resp_valid ? _GEN_355:special_entry_valid_0; 
  assign _GEN_459=io_ptw_resp_valid ? _GEN_359:superpage_entries_0_valid_0; 
  assign _GEN_463=io_ptw_resp_valid ? _GEN_363:superpage_entries_1_valid_0; 
  assign _GEN_467=io_ptw_resp_valid ? _GEN_367:superpage_entries_2_valid_0; 
  assign _GEN_471=io_ptw_resp_valid ? _GEN_371:superpage_entries_3_valid_0; 
  assign _GEN_473=io_ptw_resp_valid ? _GEN_373:sectored_entries_0_0_valid_0; 
  assign _GEN_474=io_ptw_resp_valid ? _GEN_374:sectored_entries_0_0_valid_1; 
  assign _GEN_475=io_ptw_resp_valid ? _GEN_375:sectored_entries_0_0_valid_2; 
  assign _GEN_476=io_ptw_resp_valid ? _GEN_376:sectored_entries_0_0_valid_3; 
  assign _GEN_483=io_ptw_resp_valid ? _GEN_383:sectored_entries_0_1_valid_0; 
  assign _GEN_484=io_ptw_resp_valid ? _GEN_384:sectored_entries_0_1_valid_1; 
  assign _GEN_485=io_ptw_resp_valid ? _GEN_385:sectored_entries_0_1_valid_2; 
  assign _GEN_486=io_ptw_resp_valid ? _GEN_386:sectored_entries_0_1_valid_3; 
  assign _GEN_493=io_ptw_resp_valid ? _GEN_393:sectored_entries_0_2_valid_0; 
  assign _GEN_494=io_ptw_resp_valid ? _GEN_394:sectored_entries_0_2_valid_1; 
  assign _GEN_495=io_ptw_resp_valid ? _GEN_395:sectored_entries_0_2_valid_2; 
  assign _GEN_496=io_ptw_resp_valid ? _GEN_396:sectored_entries_0_2_valid_3; 
  assign _GEN_503=io_ptw_resp_valid ? _GEN_403:sectored_entries_0_3_valid_0; 
  assign _GEN_504=io_ptw_resp_valid ? _GEN_404:sectored_entries_0_3_valid_1; 
  assign _GEN_505=io_ptw_resp_valid ? _GEN_405:sectored_entries_0_3_valid_2; 
  assign _GEN_506=io_ptw_resp_valid ? _GEN_406:sectored_entries_0_3_valid_3; 
  assign _GEN_513=io_ptw_resp_valid ? _GEN_413:sectored_entries_0_4_valid_0; 
  assign _GEN_514=io_ptw_resp_valid ? _GEN_414:sectored_entries_0_4_valid_1; 
  assign _GEN_515=io_ptw_resp_valid ? _GEN_415:sectored_entries_0_4_valid_2; 
  assign _GEN_516=io_ptw_resp_valid ? _GEN_416:sectored_entries_0_4_valid_3; 
  assign _GEN_523=io_ptw_resp_valid ? _GEN_423:sectored_entries_0_5_valid_0; 
  assign _GEN_524=io_ptw_resp_valid ? _GEN_424:sectored_entries_0_5_valid_1; 
  assign _GEN_525=io_ptw_resp_valid ? _GEN_425:sectored_entries_0_5_valid_2; 
  assign _GEN_526=io_ptw_resp_valid ? _GEN_426:sectored_entries_0_5_valid_3; 
  assign _GEN_533=io_ptw_resp_valid ? _GEN_433:sectored_entries_0_6_valid_0; 
  assign _GEN_534=io_ptw_resp_valid ? _GEN_434:sectored_entries_0_6_valid_1; 
  assign _GEN_535=io_ptw_resp_valid ? _GEN_435:sectored_entries_0_6_valid_2; 
  assign _GEN_536=io_ptw_resp_valid ? _GEN_436:sectored_entries_0_6_valid_3; 
  assign _GEN_543=io_ptw_resp_valid ? _GEN_443:sectored_entries_0_7_valid_0; 
  assign _GEN_544=io_ptw_resp_valid ? _GEN_444:sectored_entries_0_7_valid_1; 
  assign _GEN_545=io_ptw_resp_valid ? _GEN_445:sectored_entries_0_7_valid_2; 
  assign _GEN_546=io_ptw_resp_valid ? _GEN_446:sectored_entries_0_7_valid_3; 
  assign _GEN_554=2'h1==hitsVec_idx ? sectored_entries_0_0_data_1:sectored_entries_0_0_data_0; 
  assign _GEN_555=2'h2==hitsVec_idx ? sectored_entries_0_0_data_2:_GEN_554; 
  assign _GEN_556=2'h3==hitsVec_idx ? sectored_entries_0_0_data_3:_GEN_555; 
  assign _GEN_558=2'h1==hitsVec_idx ? sectored_entries_0_1_data_1:sectored_entries_0_1_data_0; 
  assign _GEN_559=2'h2==hitsVec_idx ? sectored_entries_0_1_data_2:_GEN_558; 
  assign _GEN_560=2'h3==hitsVec_idx ? sectored_entries_0_1_data_3:_GEN_559; 
  assign _GEN_562=2'h1==hitsVec_idx ? sectored_entries_0_2_data_1:sectored_entries_0_2_data_0; 
  assign _GEN_563=2'h2==hitsVec_idx ? sectored_entries_0_2_data_2:_GEN_562; 
  assign _GEN_564=2'h3==hitsVec_idx ? sectored_entries_0_2_data_3:_GEN_563; 
  assign _GEN_566=2'h1==hitsVec_idx ? sectored_entries_0_3_data_1:sectored_entries_0_3_data_0; 
  assign _GEN_567=2'h2==hitsVec_idx ? sectored_entries_0_3_data_2:_GEN_566; 
  assign _GEN_568=2'h3==hitsVec_idx ? sectored_entries_0_3_data_3:_GEN_567; 
  assign _GEN_570=2'h1==hitsVec_idx ? sectored_entries_0_4_data_1:sectored_entries_0_4_data_0; 
  assign _GEN_571=2'h2==hitsVec_idx ? sectored_entries_0_4_data_2:_GEN_570; 
  assign _GEN_572=2'h3==hitsVec_idx ? sectored_entries_0_4_data_3:_GEN_571; 
  assign _GEN_574=2'h1==hitsVec_idx ? sectored_entries_0_5_data_1:sectored_entries_0_5_data_0; 
  assign _GEN_575=2'h2==hitsVec_idx ? sectored_entries_0_5_data_2:_GEN_574; 
  assign _GEN_576=2'h3==hitsVec_idx ? sectored_entries_0_5_data_3:_GEN_575; 
  assign _GEN_578=2'h1==hitsVec_idx ? sectored_entries_0_6_data_1:sectored_entries_0_6_data_0; 
  assign _GEN_579=2'h2==hitsVec_idx ? sectored_entries_0_6_data_2:_GEN_578; 
  assign _GEN_580=2'h3==hitsVec_idx ? sectored_entries_0_6_data_3:_GEN_579; 
  assign _GEN_582=2'h1==hitsVec_idx ? sectored_entries_0_7_data_1:sectored_entries_0_7_data_0; 
  assign _GEN_583=2'h2==hitsVec_idx ? sectored_entries_0_7_data_2:_GEN_582; 
  assign _GEN_584=2'h3==hitsVec_idx ? sectored_entries_0_7_data_3:_GEN_583; 
  assign ppn_hi=entries_barrier_8_io_y_ppn[19:18]; 
  assign _ppn_T_1=superpage_hits_ignore_1 ? vpn:27'h0; 
  assign _GEN_953={7'b0,entries_barrier_8_io_y_ppn}; 
  assign _ppn_T_2=_ppn_T_1|_GEN_953; 
  assign ppn_lo=_ppn_T_2[17:9]; 
  assign _ppn_T_4=vpn|_GEN_953; 
  assign ppn_lo_1=_ppn_T_4[8:0]; 
  assign _ppn_T_5={ppn_hi,ppn_lo,ppn_lo_1}; 
  assign ppn_hi_2=entries_barrier_9_io_y_ppn[19:18]; 
  assign _ppn_T_6=superpage_hits_ignore_4 ? vpn:27'h0; 
  assign _GEN_955={7'b0,entries_barrier_9_io_y_ppn}; 
  assign _ppn_T_7=_ppn_T_6|_GEN_955; 
  assign ppn_lo_2=_ppn_T_7[17:9]; 
  assign _ppn_T_9=vpn|_GEN_955; 
  assign ppn_lo_3=_ppn_T_9[8:0]; 
  assign _ppn_T_10={ppn_hi_2,ppn_lo_2,ppn_lo_3}; 
  assign ppn_hi_4=entries_barrier_10_io_y_ppn[19:18]; 
  assign _ppn_T_11=superpage_hits_ignore_7 ? vpn:27'h0; 
  assign _GEN_957={7'b0,entries_barrier_10_io_y_ppn}; 
  assign _ppn_T_12=_ppn_T_11|_GEN_957; 
  assign ppn_lo_4=_ppn_T_12[17:9]; 
  assign _ppn_T_14=vpn|_GEN_957; 
  assign ppn_lo_5=_ppn_T_14[8:0]; 
  assign _ppn_T_15={ppn_hi_4,ppn_lo_4,ppn_lo_5}; 
  assign ppn_hi_6=entries_barrier_11_io_y_ppn[19:18]; 
  assign _ppn_T_16=superpage_hits_ignore_10 ? vpn:27'h0; 
  assign _GEN_959={7'b0,entries_barrier_11_io_y_ppn}; 
  assign _ppn_T_17=_ppn_T_16|_GEN_959; 
  assign ppn_lo_6=_ppn_T_17[17:9]; 
  assign _ppn_T_19=vpn|_GEN_959; 
  assign ppn_lo_7=_ppn_T_19[8:0]; 
  assign _ppn_T_20={ppn_hi_6,ppn_lo_6,ppn_lo_7}; 
  assign ppn_hi_8=entries_barrier_12_io_y_ppn[19:18]; 
  assign _GEN_961={7'b0,entries_barrier_12_io_y_ppn}; 
  assign _ppn_T_22=_mpu_ppn_T_17|_GEN_961; 
  assign ppn_lo_8=_ppn_T_22[17:9]; 
  assign _ppn_T_24=_mpu_ppn_T_19|_GEN_961; 
  assign ppn_lo_9=_ppn_T_24[8:0]; 
  assign _ppn_T_25={ppn_hi_8,ppn_lo_8,ppn_lo_9}; 
  assign _ppn_T_27=hitsVec_0 ? entries_barrier_io_y_ppn:20'h0; 
  assign _ppn_T_28=hitsVec_1 ? entries_barrier_1_io_y_ppn:20'h0; 
  assign _ppn_T_29=hitsVec_2 ? entries_barrier_2_io_y_ppn:20'h0; 
  assign _ppn_T_30=hitsVec_3 ? entries_barrier_3_io_y_ppn:20'h0; 
  assign _ppn_T_31=hitsVec_4 ? entries_barrier_4_io_y_ppn:20'h0; 
  assign _ppn_T_32=hitsVec_5 ? entries_barrier_5_io_y_ppn:20'h0; 
  assign _ppn_T_33=hitsVec_6 ? entries_barrier_6_io_y_ppn:20'h0; 
  assign _ppn_T_34=hitsVec_7 ? entries_barrier_7_io_y_ppn:20'h0; 
  assign _ppn_T_35=hitsVec_8 ? _ppn_T_5:20'h0; 
  assign _ppn_T_36=hitsVec_9 ? _ppn_T_10:20'h0; 
  assign _ppn_T_37=hitsVec_10 ? _ppn_T_15:20'h0; 
  assign _ppn_T_38=hitsVec_11 ? _ppn_T_20:20'h0; 
  assign _ppn_T_39=hitsVec_12 ? _ppn_T_25:20'h0; 
  assign _ppn_T_40=hits_hi ? vpn[19:0]:20'h0; 
  assign _ppn_T_41=_ppn_T_27|_ppn_T_28; 
  assign _ppn_T_42=_ppn_T_41|_ppn_T_29; 
  assign _ppn_T_43=_ppn_T_42|_ppn_T_30; 
  assign _ppn_T_44=_ppn_T_43|_ppn_T_31; 
  assign _ppn_T_45=_ppn_T_44|_ppn_T_32; 
  assign _ppn_T_46=_ppn_T_45|_ppn_T_33; 
  assign _ppn_T_47=_ppn_T_46|_ppn_T_34; 
  assign _ppn_T_48=_ppn_T_47|_ppn_T_35; 
  assign _ppn_T_49=_ppn_T_48|_ppn_T_36; 
  assign _ppn_T_50=_ppn_T_49|_ppn_T_37; 
  assign _ppn_T_51=_ppn_T_50|_ppn_T_38; 
  assign _ppn_T_52=_ppn_T_51|_ppn_T_39; 
  assign ppn=_ppn_T_52|_ppn_T_40; 
  assign ptw_ae_array_lo={entries_barrier_5_io_y_ae,entries_barrier_4_io_y_ae,entries_barrier_3_io_y_ae,entries_barrier_2_io_y_ae,entries_barrier_1_io_y_ae,entries_barrier_io_y_ae}; 
  assign ptw_ae_array={1'h0,entries_barrier_12_io_y_ae,entries_barrier_11_io_y_ae,entries_barrier_10_io_y_ae,entries_barrier_9_io_y_ae,entries_barrier_8_io_y_ae,entries_barrier_7_io_y_ae,entries_barrier_6_io_y_ae,ptw_ae_array_lo}; 
  assign _priv_rw_ok_T_1=~priv_s|io_ptw_status_sum; 
  assign priv_rw_ok_lo={entries_barrier_5_io_y_u,entries_barrier_4_io_y_u,entries_barrier_3_io_y_u,entries_barrier_2_io_y_u,entries_barrier_1_io_y_u,entries_barrier_io_y_u}; 
  assign _priv_rw_ok_T_2={entries_barrier_12_io_y_u,entries_barrier_11_io_y_u,entries_barrier_10_io_y_u,entries_barrier_9_io_y_u,entries_barrier_8_io_y_u,entries_barrier_7_io_y_u,entries_barrier_6_io_y_u,priv_rw_ok_lo}; 
  assign _priv_rw_ok_T_3=_priv_rw_ok_T_1 ? _priv_rw_ok_T_2:13'h0; 
  assign _priv_rw_ok_T_6=priv_s ? ~_priv_rw_ok_T_2:13'h0; 
  assign priv_rw_ok=_priv_rw_ok_T_3|_priv_rw_ok_T_6; 
  assign r_array_lo={entries_barrier_5_io_y_sr,entries_barrier_4_io_y_sr,entries_barrier_3_io_y_sr,entries_barrier_2_io_y_sr,entries_barrier_1_io_y_sr,entries_barrier_io_y_sr}; 
  assign _r_array_T={entries_barrier_12_io_y_sr,entries_barrier_11_io_y_sr,entries_barrier_10_io_y_sr,entries_barrier_9_io_y_sr,entries_barrier_8_io_y_sr,entries_barrier_7_io_y_sr,entries_barrier_6_io_y_sr,r_array_lo}; 
  assign r_array_lo_1={entries_barrier_5_io_y_sx,entries_barrier_4_io_y_sx,entries_barrier_3_io_y_sx,entries_barrier_2_io_y_sx,entries_barrier_1_io_y_sx,entries_barrier_io_y_sx}; 
  assign _r_array_T_1={entries_barrier_12_io_y_sx,entries_barrier_11_io_y_sx,entries_barrier_10_io_y_sx,entries_barrier_9_io_y_sx,entries_barrier_8_io_y_sx,entries_barrier_7_io_y_sx,entries_barrier_6_io_y_sx,r_array_lo_1}; 
  assign _r_array_T_2=io_ptw_status_mxr ? _r_array_T_1:13'h0; 
  assign _r_array_T_3=_r_array_T|_r_array_T_2; 
  assign r_array_lo_2=priv_rw_ok&_r_array_T_3; 
  assign r_array={1'h1,r_array_lo_2}; 
  assign w_array_lo={entries_barrier_5_io_y_sw,entries_barrier_4_io_y_sw,entries_barrier_3_io_y_sw,entries_barrier_2_io_y_sw,entries_barrier_1_io_y_sw,entries_barrier_io_y_sw}; 
  assign _w_array_T={entries_barrier_12_io_y_sw,entries_barrier_11_io_y_sw,entries_barrier_10_io_y_sw,entries_barrier_9_io_y_sw,entries_barrier_8_io_y_sw,entries_barrier_7_io_y_sw,entries_barrier_6_io_y_sw,w_array_lo}; 
  assign w_array_lo_1=priv_rw_ok&_w_array_T; 
  assign w_array={1'h1,w_array_lo_1}; 
  assign pr_array_hi=prot_r ? 2'h3:2'h0; 
  assign pr_array_lo={entries_barrier_5_io_y_pr,entries_barrier_4_io_y_pr,entries_barrier_3_io_y_pr,entries_barrier_2_io_y_pr,entries_barrier_1_io_y_pr,entries_barrier_io_y_pr}; 
  assign _pr_array_T_1={pr_array_hi,entries_barrier_11_io_y_pr,entries_barrier_10_io_y_pr,entries_barrier_9_io_y_pr,entries_barrier_8_io_y_pr,entries_barrier_7_io_y_pr,entries_barrier_6_io_y_pr,pr_array_lo}; 
  assign pr_array=_pr_array_T_1&~ptw_ae_array; 
  assign pw_array_hi=prot_w ? 2'h3:2'h0; 
  assign pw_array_lo={entries_barrier_5_io_y_pw,entries_barrier_4_io_y_pw,entries_barrier_3_io_y_pw,entries_barrier_2_io_y_pw,entries_barrier_1_io_y_pw,entries_barrier_io_y_pw}; 
  assign _pw_array_T_1={pw_array_hi,entries_barrier_11_io_y_pw,entries_barrier_10_io_y_pw,entries_barrier_9_io_y_pw,entries_barrier_8_io_y_pw,entries_barrier_7_io_y_pw,entries_barrier_6_io_y_pw,pw_array_lo}; 
  assign pw_array=_pw_array_T_1&~ptw_ae_array; 
  assign eff_array_hi=prot_eff ? 2'h3:2'h0; 
  assign eff_array_lo={entries_barrier_5_io_y_eff,entries_barrier_4_io_y_eff,entries_barrier_3_io_y_eff,entries_barrier_2_io_y_eff,entries_barrier_1_io_y_eff,entries_barrier_io_y_eff}; 
  assign eff_array={eff_array_hi,entries_barrier_11_io_y_eff,entries_barrier_10_io_y_eff,entries_barrier_9_io_y_eff,entries_barrier_8_io_y_eff,entries_barrier_7_io_y_eff,entries_barrier_6_io_y_eff,eff_array_lo}; 
  assign c_array_hi=cacheable ? 2'h3:2'h0; 
  assign c_array_lo={entries_barrier_5_io_y_c,entries_barrier_4_io_y_c,entries_barrier_3_io_y_c,entries_barrier_2_io_y_c,entries_barrier_1_io_y_c,entries_barrier_io_y_c}; 
  assign c_array={c_array_hi,entries_barrier_11_io_y_c,entries_barrier_10_io_y_c,entries_barrier_9_io_y_c,entries_barrier_8_io_y_c,entries_barrier_7_io_y_c,entries_barrier_6_io_y_c,c_array_lo}; 
  assign ppp_array_hi=_prot_w_T_31 ? 2'h3:2'h0; 
  assign ppp_array_lo={entries_barrier_5_io_y_ppp,entries_barrier_4_io_y_ppp,entries_barrier_3_io_y_ppp,entries_barrier_2_io_y_ppp,entries_barrier_1_io_y_ppp,entries_barrier_io_y_ppp}; 
  assign ppp_array={ppp_array_hi,entries_barrier_11_io_y_ppp,entries_barrier_10_io_y_ppp,entries_barrier_9_io_y_ppp,entries_barrier_8_io_y_ppp,entries_barrier_7_io_y_ppp,entries_barrier_6_io_y_ppp,ppp_array_lo}; 
  assign paa_array_hi=prot_al ? 2'h3:2'h0; 
  assign paa_array_lo={entries_barrier_5_io_y_paa,entries_barrier_4_io_y_paa,entries_barrier_3_io_y_paa,entries_barrier_2_io_y_paa,entries_barrier_1_io_y_paa,entries_barrier_io_y_paa}; 
  assign paa_array={paa_array_hi,entries_barrier_11_io_y_paa,entries_barrier_10_io_y_paa,entries_barrier_9_io_y_paa,entries_barrier_8_io_y_paa,entries_barrier_7_io_y_paa,entries_barrier_6_io_y_paa,paa_array_lo}; 
  assign pal_array_lo={entries_barrier_5_io_y_pal,entries_barrier_4_io_y_pal,entries_barrier_3_io_y_pal,entries_barrier_2_io_y_pal,entries_barrier_1_io_y_pal,entries_barrier_io_y_pal}; 
  assign pal_array={paa_array_hi,entries_barrier_11_io_y_pal,entries_barrier_10_io_y_pal,entries_barrier_9_io_y_pal,entries_barrier_8_io_y_pal,entries_barrier_7_io_y_pal,entries_barrier_6_io_y_pal,pal_array_lo}; 
  assign ppp_array_if_cached=ppp_array|c_array; 
  assign paa_array_if_cached=paa_array|c_array; 
  assign pal_array_if_cached=pal_array|c_array; 
  assign _misaligned_T=4'h1<<io_req_bits_size; 
  assign _misaligned_T_2=_misaligned_T-4'h1; 
  assign _GEN_963={36'b0,_misaligned_T_2}; 
  assign _misaligned_T_3=io_req_bits_vaddr&_GEN_963; 
  assign misaligned=|_misaligned_T_3; 
  assign bad_va_maskedVAddr=io_req_bits_vaddr&40'hc000000000; 
  assign _bad_va_T_1=bad_va_maskedVAddr==40'h0; 
  assign _bad_va_T_2=bad_va_maskedVAddr==40'hc000000000; 
  assign _bad_va_T_3=_bad_va_T_1|_bad_va_T_2; 
  assign bad_va=vm_enabled&~_bad_va_T_3; 
  assign _cmd_lrsc_T=io_req_bits_cmd==5'h6; 
  assign _cmd_lrsc_T_1=io_req_bits_cmd==5'h7; 
  assign cmd_lrsc=_cmd_lrsc_T|_cmd_lrsc_T_1; 
  assign _cmd_amo_logical_T=io_req_bits_cmd==5'h4; 
  assign _cmd_amo_logical_T_1=io_req_bits_cmd==5'h9; 
  assign _cmd_amo_logical_T_2=io_req_bits_cmd==5'ha; 
  assign _cmd_amo_logical_T_3=io_req_bits_cmd==5'hb; 
  assign _cmd_amo_logical_T_4=_cmd_amo_logical_T|_cmd_amo_logical_T_1; 
  assign _cmd_amo_logical_T_5=_cmd_amo_logical_T_4|_cmd_amo_logical_T_2; 
  assign cmd_amo_logical=_cmd_amo_logical_T_5|_cmd_amo_logical_T_3; 
  assign _cmd_amo_arithmetic_T=io_req_bits_cmd==5'h8; 
  assign _cmd_amo_arithmetic_T_1=io_req_bits_cmd==5'hc; 
  assign _cmd_amo_arithmetic_T_2=io_req_bits_cmd==5'hd; 
  assign _cmd_amo_arithmetic_T_3=io_req_bits_cmd==5'he; 
  assign _cmd_amo_arithmetic_T_4=io_req_bits_cmd==5'hf; 
  assign _cmd_amo_arithmetic_T_5=_cmd_amo_arithmetic_T|_cmd_amo_arithmetic_T_1; 
  assign _cmd_amo_arithmetic_T_6=_cmd_amo_arithmetic_T_5|_cmd_amo_arithmetic_T_2; 
  assign _cmd_amo_arithmetic_T_7=_cmd_amo_arithmetic_T_6|_cmd_amo_arithmetic_T_3; 
  assign cmd_amo_arithmetic=_cmd_amo_arithmetic_T_7|_cmd_amo_arithmetic_T_4; 
  assign cmd_put_partial=io_req_bits_cmd==5'h11; 
  assign _cmd_read_T=io_req_bits_cmd==5'h0; 
  assign _cmd_read_T_2=_cmd_read_T|_cmd_lrsc_T; 
  assign _cmd_read_T_4=_cmd_read_T_2|_cmd_lrsc_T_1; 
  assign _cmd_read_T_21=cmd_amo_logical|cmd_amo_arithmetic; 
  assign cmd_read=_cmd_read_T_4|_cmd_read_T_21; 
  assign _cmd_write_T=io_req_bits_cmd==5'h1; 
  assign _cmd_write_T_2=_cmd_write_T|cmd_put_partial; 
  assign _cmd_write_T_4=_cmd_write_T_2|_cmd_lrsc_T_1; 
  assign cmd_write=_cmd_write_T_4|_cmd_read_T_21; 
  assign _cmd_write_perms_T=io_req_bits_cmd==5'h5; 
  assign _cmd_write_perms_T_1=io_req_bits_cmd==5'h17; 
  assign _cmd_write_perms_T_2=_cmd_write_perms_T|_cmd_write_perms_T_1; 
  assign cmd_write_perms=cmd_write|_cmd_write_perms_T_2; 
  assign _ae_array_T=misaligned ? eff_array:14'h0; 
  assign _ae_array_T_2=cmd_lrsc ? ~c_array:14'h0; 
  assign ae_array=_ae_array_T|_ae_array_T_2; 
  assign _ae_ld_array_T_1=ae_array|~pr_array; 
  assign ae_ld_array=cmd_read ? _ae_ld_array_T_1:14'h0; 
  assign _ae_st_array_T_1=ae_array|~pw_array; 
  assign _ae_st_array_T_2=cmd_write_perms ? _ae_st_array_T_1:14'h0; 
  assign _ae_st_array_T_4=cmd_put_partial ? ~ppp_array_if_cached:14'h0; 
  assign _ae_st_array_T_5=_ae_st_array_T_2|_ae_st_array_T_4; 
  assign _ae_st_array_T_7=cmd_amo_logical ? ~pal_array_if_cached:14'h0; 
  assign _ae_st_array_T_8=_ae_st_array_T_5|_ae_st_array_T_7; 
  assign _ae_st_array_T_10=cmd_amo_arithmetic ? ~paa_array_if_cached:14'h0; 
  assign ae_st_array=_ae_st_array_T_8|_ae_st_array_T_10; 
  assign _ma_ld_array_T=misaligned&cmd_read; 
  assign ma_ld_array=_ma_ld_array_T ? ~eff_array:14'h0; 
  assign _ma_st_array_T=misaligned&cmd_write; 
  assign ma_st_array=_ma_st_array_T ? ~eff_array:14'h0; 
  assign _pf_ld_array_T=r_array|ptw_ae_array; 
  assign pf_ld_array=cmd_read ? ~_pf_ld_array_T:14'h0; 
  assign _pf_st_array_T=w_array|ptw_ae_array; 
  assign pf_st_array=cmd_write_perms ? ~_pf_st_array_T:14'h0; 
  assign tlb_hit=|real_hits; 
  assign _tlb_miss_T_1=vm_enabled&~bad_va; 
  assign tlb_miss=_tlb_miss_T_1&~tlb_hit; 
  assign _T_23=io_req_valid&vm_enabled; 
  assign _T_24=sector_hits_0|sector_hits_1; 
  assign _T_25=_T_24|sector_hits_2; 
  assign _T_26=_T_25|sector_hits_3; 
  assign _T_27=_T_26|sector_hits_4; 
  assign _T_28=_T_27|sector_hits_5; 
  assign _T_29=_T_28|sector_hits_6; 
  assign _T_30=_T_29|sector_hits_7; 
  assign _T_31={sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; 
  assign hi_1=_T_31[7:4]; 
  assign lo_1=_T_31[3:0]; 
  assign hi_2=|hi_1; 
  assign _T_32=hi_1|lo_1; 
  assign hi_3=_T_32[3:2]; 
  assign lo_2=_T_32[1:0]; 
  assign hi_4=|hi_3; 
  assign _T_33=hi_3|lo_2; 
  assign lo_3=_T_33[1]; 
  assign state_vec_0_touch_way_sized={hi_2,hi_4,lo_3}; 
  assign state_vec_0_hi_hi=~state_vec_0_touch_way_sized[2]; 
  assign state_vec_0_left_subtree_state=state_vec_0[5:3]; 
  assign state_vec_0_right_subtree_state=state_vec_0[2:0]; 
  assign state_vec_0_hi_hi_1=~state_vec_0_touch_way_sized[1]; 
  assign state_vec_0_left_subtree_state_1=state_vec_0_left_subtree_state[1]; 
  assign state_vec_0_right_subtree_state_1=state_vec_0_left_subtree_state[0]; 
  assign state_vec_0_hi_lo=state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_1:~state_vec_0_touch_way_sized[0]; 
  assign state_vec_0_lo=state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0]:state_vec_0_right_subtree_state_1; 
  assign _state_vec_0_T_7={state_vec_0_hi_hi_1,state_vec_0_hi_lo,state_vec_0_lo}; 
  assign state_vec_0_hi_lo_1=state_vec_0_hi_hi ? state_vec_0_left_subtree_state:_state_vec_0_T_7; 
  assign state_vec_0_left_subtree_state_2=state_vec_0_right_subtree_state[1]; 
  assign state_vec_0_right_subtree_state_2=state_vec_0_right_subtree_state[0]; 
  assign state_vec_0_hi_lo_2=state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_2:~state_vec_0_touch_way_sized[0]; 
  assign state_vec_0_lo_1=state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0]:state_vec_0_right_subtree_state_2; 
  assign _state_vec_0_T_15={state_vec_0_hi_hi_1,state_vec_0_hi_lo_2,state_vec_0_lo_1}; 
  assign state_vec_0_lo_2=state_vec_0_hi_hi ? _state_vec_0_T_15:state_vec_0_right_subtree_state; 
  assign _state_vec_0_T_16={state_vec_0_hi_hi,state_vec_0_hi_lo_1,state_vec_0_lo_2}; 
  assign _T_35=superpage_hits_0|superpage_hits_1; 
  assign _T_36=_T_35|superpage_hits_2; 
  assign _T_37=_T_36|superpage_hits_3; 
  assign _T_38={superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; 
  assign hi_6=_T_38[3:2]; 
  assign lo_6=_T_38[1:0]; 
  assign hi_7=|hi_6; 
  assign _T_39=hi_6|lo_6; 
  assign lo_7=_T_39[1]; 
  assign state_reg_touch_way_sized={hi_7,lo_7}; 
  assign state_reg_hi_hi=~state_reg_touch_way_sized[1]; 
  assign state_reg_left_subtree_state=state_reg_1[1]; 
  assign state_reg_right_subtree_state=state_reg_1[0]; 
  assign state_reg_hi_lo=state_reg_hi_hi ? state_reg_left_subtree_state:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo=state_reg_hi_hi ? ~state_reg_touch_way_sized[0]:state_reg_right_subtree_state; 
  assign _state_reg_T_6={state_reg_hi_hi,state_reg_hi_lo,state_reg_lo}; 
  assign multipleHits_leftOne=real_hits[0]; 
  assign multipleHits_leftOne_1=real_hits[1]; 
  assign multipleHits_rightOne=real_hits[2]; 
  assign multipleHits_rightOne_1=multipleHits_leftOne_1|multipleHits_rightOne; 
  assign multipleHits_rightTwo=multipleHits_leftOne_1&multipleHits_rightOne; 
  assign multipleHits_leftOne_2=multipleHits_leftOne|multipleHits_rightOne_1; 
  assign _multipleHits_T_9=multipleHits_leftOne&multipleHits_rightOne_1; 
  assign multipleHits_leftTwo=multipleHits_rightTwo|_multipleHits_T_9; 
  assign multipleHits_leftOne_3=real_hits[3]; 
  assign multipleHits_leftOne_4=real_hits[4]; 
  assign multipleHits_rightOne_2=real_hits[5]; 
  assign multipleHits_rightOne_3=multipleHits_leftOne_4|multipleHits_rightOne_2; 
  assign multipleHits_rightTwo_1=multipleHits_leftOne_4&multipleHits_rightOne_2; 
  assign multipleHits_rightOne_4=multipleHits_leftOne_3|multipleHits_rightOne_3; 
  assign _multipleHits_T_18=multipleHits_leftOne_3&multipleHits_rightOne_3; 
  assign multipleHits_rightTwo_2=multipleHits_rightTwo_1|_multipleHits_T_18; 
  assign multipleHits_leftOne_5=multipleHits_leftOne_2|multipleHits_rightOne_4; 
  assign _multipleHits_T_19=multipleHits_leftTwo|multipleHits_rightTwo_2; 
  assign _multipleHits_T_20=multipleHits_leftOne_2&multipleHits_rightOne_4; 
  assign multipleHits_leftTwo_1=_multipleHits_T_19|_multipleHits_T_20; 
  assign multipleHits_leftOne_6=real_hits[6]; 
  assign multipleHits_leftOne_7=real_hits[7]; 
  assign multipleHits_rightOne_5=real_hits[8]; 
  assign multipleHits_rightOne_6=multipleHits_leftOne_7|multipleHits_rightOne_5; 
  assign multipleHits_rightTwo_3=multipleHits_leftOne_7&multipleHits_rightOne_5; 
  assign multipleHits_leftOne_8=multipleHits_leftOne_6|multipleHits_rightOne_6; 
  assign _multipleHits_T_30=multipleHits_leftOne_6&multipleHits_rightOne_6; 
  assign multipleHits_leftTwo_2=multipleHits_rightTwo_3|_multipleHits_T_30; 
  assign multipleHits_leftOne_9=real_hits[9]; 
  assign multipleHits_rightOne_7=real_hits[10]; 
  assign multipleHits_leftOne_10=multipleHits_leftOne_9|multipleHits_rightOne_7; 
  assign multipleHits_leftTwo_3=multipleHits_leftOne_9&multipleHits_rightOne_7; 
  assign multipleHits_leftOne_11=real_hits[11]; 
  assign multipleHits_rightOne_8=real_hits[12]; 
  assign multipleHits_rightOne_9=multipleHits_leftOne_11|multipleHits_rightOne_8; 
  assign multipleHits_rightTwo_4=multipleHits_leftOne_11&multipleHits_rightOne_8; 
  assign multipleHits_rightOne_10=multipleHits_leftOne_10|multipleHits_rightOne_9; 
  assign _multipleHits_T_42=multipleHits_leftTwo_3|multipleHits_rightTwo_4; 
  assign _multipleHits_T_43=multipleHits_leftOne_10&multipleHits_rightOne_9; 
  assign multipleHits_rightTwo_5=_multipleHits_T_42|_multipleHits_T_43; 
  assign multipleHits_rightOne_11=multipleHits_leftOne_8|multipleHits_rightOne_10; 
  assign _multipleHits_T_44=multipleHits_leftTwo_2|multipleHits_rightTwo_5; 
  assign _multipleHits_T_45=multipleHits_leftOne_8&multipleHits_rightOne_10; 
  assign multipleHits_rightTwo_6=_multipleHits_T_44|_multipleHits_T_45; 
  assign _multipleHits_T_47=multipleHits_leftTwo_1|multipleHits_rightTwo_6; 
  assign _multipleHits_T_48=multipleHits_leftOne_5&multipleHits_rightOne_11; 
  assign multipleHits=_multipleHits_T_47|_multipleHits_T_48; 
  assign _io_resp_pf_ld_T=bad_va&cmd_read; 
  assign _io_resp_pf_ld_T_1=pf_ld_array&hits; 
  assign _io_resp_pf_ld_T_2=|_io_resp_pf_ld_T_1; 
  assign _io_resp_pf_st_T=bad_va&cmd_write_perms; 
  assign _io_resp_pf_st_T_1=pf_st_array&hits; 
  assign _io_resp_pf_st_T_2=|_io_resp_pf_st_T_1; 
  assign _io_resp_ae_ld_T=ae_ld_array&hits; 
  assign _io_resp_ae_st_T=ae_st_array&hits; 
  assign _io_resp_ma_ld_T=ma_ld_array&hits; 
  assign _io_resp_ma_st_T=ma_st_array&hits; 
  assign _io_resp_cacheable_T=c_array&hits; 
  assign _io_resp_miss_T=io_ptw_resp_valid|tlb_miss; 
  assign _T_41=io_req_ready&io_req_valid; 
  assign _T_42=_T_41&tlb_miss; 
  assign r_superpage_repl_addr_hi=state_reg_1[2]; 
  assign r_superpage_repl_addr_lo=r_superpage_repl_addr_hi ? state_reg_left_subtree_state:state_reg_right_subtree_state; 
  assign _r_superpage_repl_addr_T_2={r_superpage_repl_addr_hi,r_superpage_repl_addr_lo}; 
  assign r_superpage_repl_addr_valids={superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; 
  assign _r_superpage_repl_addr_T_3=&r_superpage_repl_addr_valids; 
  assign _r_superpage_repl_addr_T_5=~r_superpage_repl_addr_valids[0]; 
  assign _r_superpage_repl_addr_T_6=~r_superpage_repl_addr_valids[1]; 
  assign _r_superpage_repl_addr_T_7=~r_superpage_repl_addr_valids[2]; 
  assign r_sectored_repl_addr_hi=state_vec_0[6]; 
  assign r_sectored_repl_addr_hi_1=state_vec_0_left_subtree_state[2]; 
  assign r_sectored_repl_addr_lo=r_sectored_repl_addr_hi_1 ? state_vec_0_left_subtree_state_1:state_vec_0_right_subtree_state_1; 
  assign _r_sectored_repl_addr_T_2={r_sectored_repl_addr_hi_1,r_sectored_repl_addr_lo}; 
  assign r_sectored_repl_addr_hi_2=state_vec_0_right_subtree_state[2]; 
  assign r_sectored_repl_addr_lo_1=r_sectored_repl_addr_hi_2 ? state_vec_0_left_subtree_state_2:state_vec_0_right_subtree_state_2; 
  assign _r_sectored_repl_addr_T_5={r_sectored_repl_addr_hi_2,r_sectored_repl_addr_lo_1}; 
  assign r_sectored_repl_addr_lo_2=r_sectored_repl_addr_hi ? _r_sectored_repl_addr_T_2:_r_sectored_repl_addr_T_5; 
  assign _r_sectored_repl_addr_T_6={r_sectored_repl_addr_hi,r_sectored_repl_addr_lo_2}; 
  assign r_sectored_repl_addr_valids={_sector_hits_T_44,_sector_hits_T_38,_sector_hits_T_32,_sector_hits_T_26,_sector_hits_T_20,_sector_hits_T_14,_sector_hits_T_8,_sector_hits_T_2}; 
  assign _r_sectored_repl_addr_T_7=&r_sectored_repl_addr_valids; 
  assign _r_sectored_repl_addr_T_9=~r_sectored_repl_addr_valids[0]; 
  assign _r_sectored_repl_addr_T_10=~r_sectored_repl_addr_valids[1]; 
  assign _r_sectored_repl_addr_T_11=~r_sectored_repl_addr_valids[2]; 
  assign _r_sectored_repl_addr_T_12=~r_sectored_repl_addr_valids[3]; 
  assign _r_sectored_repl_addr_T_13=~r_sectored_repl_addr_valids[4]; 
  assign _r_sectored_repl_addr_T_14=~r_sectored_repl_addr_valids[5]; 
  assign _r_sectored_repl_addr_T_15=~r_sectored_repl_addr_valids[6]; 
  assign _T_44=state==2'h2; 
  assign _T_45=_T_44&io_sfence_valid; 
  assign _T_48=io_sfence_bits_addr[38:12]==vpn; 
  assign _T_49=~io_sfence_bits_rs1|_T_48; 
  assign _T_51=_T_49|reset; 
  assign _T_59=_sector_hits_T_3[26:18]==9'h0; 
  assign _GEN_617=sectored_entries_0_0_data_0[13] ? _GEN_473:1'h0; 
  assign _GEN_618=sectored_entries_0_0_data_1[13] ? _GEN_474:1'h0; 
  assign _GEN_619=sectored_entries_0_0_data_2[13] ? _GEN_475:1'h0; 
  assign _GEN_620=sectored_entries_0_0_data_3[13] ? _GEN_476:1'h0; 
  assign _GEN_621=io_sfence_bits_rs2&_GEN_617; 
  assign _GEN_622=io_sfence_bits_rs2&_GEN_618; 
  assign _GEN_623=io_sfence_bits_rs2&_GEN_619; 
  assign _GEN_624=io_sfence_bits_rs2&_GEN_620; 
  assign _T_198=_sector_hits_T_9[26:18]==9'h0; 
  assign _GEN_645=sectored_entries_0_1_data_0[13] ? _GEN_483:1'h0; 
  assign _GEN_646=sectored_entries_0_1_data_1[13] ? _GEN_484:1'h0; 
  assign _GEN_647=sectored_entries_0_1_data_2[13] ? _GEN_485:1'h0; 
  assign _GEN_648=sectored_entries_0_1_data_3[13] ? _GEN_486:1'h0; 
  assign _GEN_649=io_sfence_bits_rs2&_GEN_645; 
  assign _GEN_650=io_sfence_bits_rs2&_GEN_646; 
  assign _GEN_651=io_sfence_bits_rs2&_GEN_647; 
  assign _GEN_652=io_sfence_bits_rs2&_GEN_648; 
  assign _T_337=_sector_hits_T_15[26:18]==9'h0; 
  assign _GEN_673=sectored_entries_0_2_data_0[13] ? _GEN_493:1'h0; 
  assign _GEN_674=sectored_entries_0_2_data_1[13] ? _GEN_494:1'h0; 
  assign _GEN_675=sectored_entries_0_2_data_2[13] ? _GEN_495:1'h0; 
  assign _GEN_676=sectored_entries_0_2_data_3[13] ? _GEN_496:1'h0; 
  assign _GEN_677=io_sfence_bits_rs2&_GEN_673; 
  assign _GEN_678=io_sfence_bits_rs2&_GEN_674; 
  assign _GEN_679=io_sfence_bits_rs2&_GEN_675; 
  assign _GEN_680=io_sfence_bits_rs2&_GEN_676; 
  assign _T_476=_sector_hits_T_21[26:18]==9'h0; 
  assign _GEN_701=sectored_entries_0_3_data_0[13] ? _GEN_503:1'h0; 
  assign _GEN_702=sectored_entries_0_3_data_1[13] ? _GEN_504:1'h0; 
  assign _GEN_703=sectored_entries_0_3_data_2[13] ? _GEN_505:1'h0; 
  assign _GEN_704=sectored_entries_0_3_data_3[13] ? _GEN_506:1'h0; 
  assign _GEN_705=io_sfence_bits_rs2&_GEN_701; 
  assign _GEN_706=io_sfence_bits_rs2&_GEN_702; 
  assign _GEN_707=io_sfence_bits_rs2&_GEN_703; 
  assign _GEN_708=io_sfence_bits_rs2&_GEN_704; 
  assign _T_615=_sector_hits_T_27[26:18]==9'h0; 
  assign _GEN_729=sectored_entries_0_4_data_0[13] ? _GEN_513:1'h0; 
  assign _GEN_730=sectored_entries_0_4_data_1[13] ? _GEN_514:1'h0; 
  assign _GEN_731=sectored_entries_0_4_data_2[13] ? _GEN_515:1'h0; 
  assign _GEN_732=sectored_entries_0_4_data_3[13] ? _GEN_516:1'h0; 
  assign _GEN_733=io_sfence_bits_rs2&_GEN_729; 
  assign _GEN_734=io_sfence_bits_rs2&_GEN_730; 
  assign _GEN_735=io_sfence_bits_rs2&_GEN_731; 
  assign _GEN_736=io_sfence_bits_rs2&_GEN_732; 
  assign _T_754=_sector_hits_T_33[26:18]==9'h0; 
  assign _GEN_757=sectored_entries_0_5_data_0[13] ? _GEN_523:1'h0; 
  assign _GEN_758=sectored_entries_0_5_data_1[13] ? _GEN_524:1'h0; 
  assign _GEN_759=sectored_entries_0_5_data_2[13] ? _GEN_525:1'h0; 
  assign _GEN_760=sectored_entries_0_5_data_3[13] ? _GEN_526:1'h0; 
  assign _GEN_761=io_sfence_bits_rs2&_GEN_757; 
  assign _GEN_762=io_sfence_bits_rs2&_GEN_758; 
  assign _GEN_763=io_sfence_bits_rs2&_GEN_759; 
  assign _GEN_764=io_sfence_bits_rs2&_GEN_760; 
  assign _T_893=_sector_hits_T_39[26:18]==9'h0; 
  assign _GEN_785=sectored_entries_0_6_data_0[13] ? _GEN_533:1'h0; 
  assign _GEN_786=sectored_entries_0_6_data_1[13] ? _GEN_534:1'h0; 
  assign _GEN_787=sectored_entries_0_6_data_2[13] ? _GEN_535:1'h0; 
  assign _GEN_788=sectored_entries_0_6_data_3[13] ? _GEN_536:1'h0; 
  assign _GEN_789=io_sfence_bits_rs2&_GEN_785; 
  assign _GEN_790=io_sfence_bits_rs2&_GEN_786; 
  assign _GEN_791=io_sfence_bits_rs2&_GEN_787; 
  assign _GEN_792=io_sfence_bits_rs2&_GEN_788; 
  assign _T_1032=_sector_hits_T_45[26:18]==9'h0; 
  assign _GEN_813=sectored_entries_0_7_data_0[13] ? _GEN_543:1'h0; 
  assign _GEN_814=sectored_entries_0_7_data_1[13] ? _GEN_544:1'h0; 
  assign _GEN_815=sectored_entries_0_7_data_2[13] ? _GEN_545:1'h0; 
  assign _GEN_816=sectored_entries_0_7_data_3[13] ? _GEN_546:1'h0; 
  assign _GEN_817=io_sfence_bits_rs2&_GEN_813; 
  assign _GEN_818=io_sfence_bits_rs2&_GEN_814; 
  assign _GEN_819=io_sfence_bits_rs2&_GEN_815; 
  assign _GEN_820=io_sfence_bits_rs2&_GEN_816; 
  assign _GEN_826=superpage_entries_0_data_0[13] ? _GEN_459:1'h0; 
  assign _GEN_827=io_sfence_bits_rs2&_GEN_826; 
  assign _GEN_830=superpage_entries_1_data_0[13] ? _GEN_463:1'h0; 
  assign _GEN_831=io_sfence_bits_rs2&_GEN_830; 
  assign _GEN_834=superpage_entries_2_data_0[13] ? _GEN_467:1'h0; 
  assign _GEN_835=io_sfence_bits_rs2&_GEN_834; 
  assign _GEN_838=superpage_entries_3_data_0[13] ? _GEN_471:1'h0; 
  assign _GEN_839=io_sfence_bits_rs2&_GEN_838; 
  assign _GEN_842=special_entry_data_0[13] ? _GEN_455:1'h0; 
  assign _GEN_843=io_sfence_bits_rs2&_GEN_842; 
  assign _T_1326=multipleHits|reset; 
  assign io_req_ready=state==2'h0; 
  assign io_resp_miss=_io_resp_miss_T|multipleHits; 
  assign io_resp_paddr={ppn,mpu_physaddr_lo}; 
  assign io_resp_pf_ld=_io_resp_pf_ld_T|_io_resp_pf_ld_T_2; 
  assign io_resp_pf_st=_io_resp_pf_st_T|_io_resp_pf_st_T_2; 
  assign io_resp_ae_ld=|_io_resp_ae_ld_T; 
  assign io_resp_ae_st=|_io_resp_ae_st_T; 
  assign io_resp_ma_ld=|_io_resp_ma_ld_T; 
  assign io_resp_ma_st=|_io_resp_ma_st_T; 
  assign io_resp_cacheable=|_io_resp_cacheable_T; 
  assign io_ptw_req_valid=state==2'h1; 
  assign io_ptw_req_bits_bits_addr=r_refill_tag; 
  assign mpu_ppn_barrier_io_x_ppn=special_entry_data_0[34:15]; 
  assign mpu_ppn_barrier_io_x_u=special_entry_data_0[14]; 
  assign mpu_ppn_barrier_io_x_ae=special_entry_data_0[12]; 
  assign mpu_ppn_barrier_io_x_sw=special_entry_data_0[11]; 
  assign mpu_ppn_barrier_io_x_sx=special_entry_data_0[10]; 
  assign mpu_ppn_barrier_io_x_sr=special_entry_data_0[9]; 
  assign mpu_ppn_barrier_io_x_pw=special_entry_data_0[8]; 
  assign mpu_ppn_barrier_io_x_px=special_entry_data_0[7]; 
  assign mpu_ppn_barrier_io_x_pr=special_entry_data_0[6]; 
  assign mpu_ppn_barrier_io_x_ppp=special_entry_data_0[5]; 
  assign mpu_ppn_barrier_io_x_pal=special_entry_data_0[4]; 
  assign mpu_ppn_barrier_io_x_paa=special_entry_data_0[3]; 
  assign mpu_ppn_barrier_io_x_eff=special_entry_data_0[2]; 
  assign mpu_ppn_barrier_io_x_c=special_entry_data_0[1]; 
  assign pmp_io_prv=mpu_priv[1:0]; 
  assign pmp_io_pmp_0_cfg_l=io_ptw_pmp_0_cfg_l; 
  assign pmp_io_pmp_0_cfg_a=io_ptw_pmp_0_cfg_a; 
  assign pmp_io_pmp_0_cfg_x=io_ptw_pmp_0_cfg_x; 
  assign pmp_io_pmp_0_cfg_w=io_ptw_pmp_0_cfg_w; 
  assign pmp_io_pmp_0_cfg_r=io_ptw_pmp_0_cfg_r; 
  assign pmp_io_pmp_0_addr=io_ptw_pmp_0_addr; 
  assign pmp_io_pmp_0_mask=io_ptw_pmp_0_mask; 
  assign pmp_io_pmp_1_cfg_l=io_ptw_pmp_1_cfg_l; 
  assign pmp_io_pmp_1_cfg_a=io_ptw_pmp_1_cfg_a; 
  assign pmp_io_pmp_1_cfg_x=io_ptw_pmp_1_cfg_x; 
  assign pmp_io_pmp_1_cfg_w=io_ptw_pmp_1_cfg_w; 
  assign pmp_io_pmp_1_cfg_r=io_ptw_pmp_1_cfg_r; 
  assign pmp_io_pmp_1_addr=io_ptw_pmp_1_addr; 
  assign pmp_io_pmp_1_mask=io_ptw_pmp_1_mask; 
  assign pmp_io_pmp_2_cfg_l=io_ptw_pmp_2_cfg_l; 
  assign pmp_io_pmp_2_cfg_a=io_ptw_pmp_2_cfg_a; 
  assign pmp_io_pmp_2_cfg_x=io_ptw_pmp_2_cfg_x; 
  assign pmp_io_pmp_2_cfg_w=io_ptw_pmp_2_cfg_w; 
  assign pmp_io_pmp_2_cfg_r=io_ptw_pmp_2_cfg_r; 
  assign pmp_io_pmp_2_addr=io_ptw_pmp_2_addr; 
  assign pmp_io_pmp_2_mask=io_ptw_pmp_2_mask; 
  assign pmp_io_pmp_3_cfg_l=io_ptw_pmp_3_cfg_l; 
  assign pmp_io_pmp_3_cfg_a=io_ptw_pmp_3_cfg_a; 
  assign pmp_io_pmp_3_cfg_x=io_ptw_pmp_3_cfg_x; 
  assign pmp_io_pmp_3_cfg_w=io_ptw_pmp_3_cfg_w; 
  assign pmp_io_pmp_3_cfg_r=io_ptw_pmp_3_cfg_r; 
  assign pmp_io_pmp_3_addr=io_ptw_pmp_3_addr; 
  assign pmp_io_pmp_3_mask=io_ptw_pmp_3_mask; 
  assign pmp_io_pmp_4_cfg_l=io_ptw_pmp_4_cfg_l; 
  assign pmp_io_pmp_4_cfg_a=io_ptw_pmp_4_cfg_a; 
  assign pmp_io_pmp_4_cfg_x=io_ptw_pmp_4_cfg_x; 
  assign pmp_io_pmp_4_cfg_w=io_ptw_pmp_4_cfg_w; 
  assign pmp_io_pmp_4_cfg_r=io_ptw_pmp_4_cfg_r; 
  assign pmp_io_pmp_4_addr=io_ptw_pmp_4_addr; 
  assign pmp_io_pmp_4_mask=io_ptw_pmp_4_mask; 
  assign pmp_io_pmp_5_cfg_l=io_ptw_pmp_5_cfg_l; 
  assign pmp_io_pmp_5_cfg_a=io_ptw_pmp_5_cfg_a; 
  assign pmp_io_pmp_5_cfg_x=io_ptw_pmp_5_cfg_x; 
  assign pmp_io_pmp_5_cfg_w=io_ptw_pmp_5_cfg_w; 
  assign pmp_io_pmp_5_cfg_r=io_ptw_pmp_5_cfg_r; 
  assign pmp_io_pmp_5_addr=io_ptw_pmp_5_addr; 
  assign pmp_io_pmp_5_mask=io_ptw_pmp_5_mask; 
  assign pmp_io_pmp_6_cfg_l=io_ptw_pmp_6_cfg_l; 
  assign pmp_io_pmp_6_cfg_a=io_ptw_pmp_6_cfg_a; 
  assign pmp_io_pmp_6_cfg_x=io_ptw_pmp_6_cfg_x; 
  assign pmp_io_pmp_6_cfg_w=io_ptw_pmp_6_cfg_w; 
  assign pmp_io_pmp_6_cfg_r=io_ptw_pmp_6_cfg_r; 
  assign pmp_io_pmp_6_addr=io_ptw_pmp_6_addr; 
  assign pmp_io_pmp_6_mask=io_ptw_pmp_6_mask; 
  assign pmp_io_pmp_7_cfg_l=io_ptw_pmp_7_cfg_l; 
  assign pmp_io_pmp_7_cfg_a=io_ptw_pmp_7_cfg_a; 
  assign pmp_io_pmp_7_cfg_x=io_ptw_pmp_7_cfg_x; 
  assign pmp_io_pmp_7_cfg_w=io_ptw_pmp_7_cfg_w; 
  assign pmp_io_pmp_7_cfg_r=io_ptw_pmp_7_cfg_r; 
  assign pmp_io_pmp_7_addr=io_ptw_pmp_7_addr; 
  assign pmp_io_pmp_7_mask=io_ptw_pmp_7_mask; 
  assign pmp_io_addr=mpu_physaddr[31:0]; 
  assign pmp_io_size=io_req_bits_size; 
  assign entries_barrier_io_x_ppn=_GEN_556[34:15]; 
  assign entries_barrier_io_x_u=_GEN_556[14]; 
  assign entries_barrier_io_x_ae=_GEN_556[12]; 
  assign entries_barrier_io_x_sw=_GEN_556[11]; 
  assign entries_barrier_io_x_sx=_GEN_556[10]; 
  assign entries_barrier_io_x_sr=_GEN_556[9]; 
  assign entries_barrier_io_x_pw=_GEN_556[8]; 
  assign entries_barrier_io_x_px=_GEN_556[7]; 
  assign entries_barrier_io_x_pr=_GEN_556[6]; 
  assign entries_barrier_io_x_ppp=_GEN_556[5]; 
  assign entries_barrier_io_x_pal=_GEN_556[4]; 
  assign entries_barrier_io_x_paa=_GEN_556[3]; 
  assign entries_barrier_io_x_eff=_GEN_556[2]; 
  assign entries_barrier_io_x_c=_GEN_556[1]; 
  assign entries_barrier_1_io_x_ppn=_GEN_560[34:15]; 
  assign entries_barrier_1_io_x_u=_GEN_560[14]; 
  assign entries_barrier_1_io_x_ae=_GEN_560[12]; 
  assign entries_barrier_1_io_x_sw=_GEN_560[11]; 
  assign entries_barrier_1_io_x_sx=_GEN_560[10]; 
  assign entries_barrier_1_io_x_sr=_GEN_560[9]; 
  assign entries_barrier_1_io_x_pw=_GEN_560[8]; 
  assign entries_barrier_1_io_x_px=_GEN_560[7]; 
  assign entries_barrier_1_io_x_pr=_GEN_560[6]; 
  assign entries_barrier_1_io_x_ppp=_GEN_560[5]; 
  assign entries_barrier_1_io_x_pal=_GEN_560[4]; 
  assign entries_barrier_1_io_x_paa=_GEN_560[3]; 
  assign entries_barrier_1_io_x_eff=_GEN_560[2]; 
  assign entries_barrier_1_io_x_c=_GEN_560[1]; 
  assign entries_barrier_2_io_x_ppn=_GEN_564[34:15]; 
  assign entries_barrier_2_io_x_u=_GEN_564[14]; 
  assign entries_barrier_2_io_x_ae=_GEN_564[12]; 
  assign entries_barrier_2_io_x_sw=_GEN_564[11]; 
  assign entries_barrier_2_io_x_sx=_GEN_564[10]; 
  assign entries_barrier_2_io_x_sr=_GEN_564[9]; 
  assign entries_barrier_2_io_x_pw=_GEN_564[8]; 
  assign entries_barrier_2_io_x_px=_GEN_564[7]; 
  assign entries_barrier_2_io_x_pr=_GEN_564[6]; 
  assign entries_barrier_2_io_x_ppp=_GEN_564[5]; 
  assign entries_barrier_2_io_x_pal=_GEN_564[4]; 
  assign entries_barrier_2_io_x_paa=_GEN_564[3]; 
  assign entries_barrier_2_io_x_eff=_GEN_564[2]; 
  assign entries_barrier_2_io_x_c=_GEN_564[1]; 
  assign entries_barrier_3_io_x_ppn=_GEN_568[34:15]; 
  assign entries_barrier_3_io_x_u=_GEN_568[14]; 
  assign entries_barrier_3_io_x_ae=_GEN_568[12]; 
  assign entries_barrier_3_io_x_sw=_GEN_568[11]; 
  assign entries_barrier_3_io_x_sx=_GEN_568[10]; 
  assign entries_barrier_3_io_x_sr=_GEN_568[9]; 
  assign entries_barrier_3_io_x_pw=_GEN_568[8]; 
  assign entries_barrier_3_io_x_px=_GEN_568[7]; 
  assign entries_barrier_3_io_x_pr=_GEN_568[6]; 
  assign entries_barrier_3_io_x_ppp=_GEN_568[5]; 
  assign entries_barrier_3_io_x_pal=_GEN_568[4]; 
  assign entries_barrier_3_io_x_paa=_GEN_568[3]; 
  assign entries_barrier_3_io_x_eff=_GEN_568[2]; 
  assign entries_barrier_3_io_x_c=_GEN_568[1]; 
  assign entries_barrier_4_io_x_ppn=_GEN_572[34:15]; 
  assign entries_barrier_4_io_x_u=_GEN_572[14]; 
  assign entries_barrier_4_io_x_ae=_GEN_572[12]; 
  assign entries_barrier_4_io_x_sw=_GEN_572[11]; 
  assign entries_barrier_4_io_x_sx=_GEN_572[10]; 
  assign entries_barrier_4_io_x_sr=_GEN_572[9]; 
  assign entries_barrier_4_io_x_pw=_GEN_572[8]; 
  assign entries_barrier_4_io_x_px=_GEN_572[7]; 
  assign entries_barrier_4_io_x_pr=_GEN_572[6]; 
  assign entries_barrier_4_io_x_ppp=_GEN_572[5]; 
  assign entries_barrier_4_io_x_pal=_GEN_572[4]; 
  assign entries_barrier_4_io_x_paa=_GEN_572[3]; 
  assign entries_barrier_4_io_x_eff=_GEN_572[2]; 
  assign entries_barrier_4_io_x_c=_GEN_572[1]; 
  assign entries_barrier_5_io_x_ppn=_GEN_576[34:15]; 
  assign entries_barrier_5_io_x_u=_GEN_576[14]; 
  assign entries_barrier_5_io_x_ae=_GEN_576[12]; 
  assign entries_barrier_5_io_x_sw=_GEN_576[11]; 
  assign entries_barrier_5_io_x_sx=_GEN_576[10]; 
  assign entries_barrier_5_io_x_sr=_GEN_576[9]; 
  assign entries_barrier_5_io_x_pw=_GEN_576[8]; 
  assign entries_barrier_5_io_x_px=_GEN_576[7]; 
  assign entries_barrier_5_io_x_pr=_GEN_576[6]; 
  assign entries_barrier_5_io_x_ppp=_GEN_576[5]; 
  assign entries_barrier_5_io_x_pal=_GEN_576[4]; 
  assign entries_barrier_5_io_x_paa=_GEN_576[3]; 
  assign entries_barrier_5_io_x_eff=_GEN_576[2]; 
  assign entries_barrier_5_io_x_c=_GEN_576[1]; 
  assign entries_barrier_6_io_x_ppn=_GEN_580[34:15]; 
  assign entries_barrier_6_io_x_u=_GEN_580[14]; 
  assign entries_barrier_6_io_x_ae=_GEN_580[12]; 
  assign entries_barrier_6_io_x_sw=_GEN_580[11]; 
  assign entries_barrier_6_io_x_sx=_GEN_580[10]; 
  assign entries_barrier_6_io_x_sr=_GEN_580[9]; 
  assign entries_barrier_6_io_x_pw=_GEN_580[8]; 
  assign entries_barrier_6_io_x_px=_GEN_580[7]; 
  assign entries_barrier_6_io_x_pr=_GEN_580[6]; 
  assign entries_barrier_6_io_x_ppp=_GEN_580[5]; 
  assign entries_barrier_6_io_x_pal=_GEN_580[4]; 
  assign entries_barrier_6_io_x_paa=_GEN_580[3]; 
  assign entries_barrier_6_io_x_eff=_GEN_580[2]; 
  assign entries_barrier_6_io_x_c=_GEN_580[1]; 
  assign entries_barrier_7_io_x_ppn=_GEN_584[34:15]; 
  assign entries_barrier_7_io_x_u=_GEN_584[14]; 
  assign entries_barrier_7_io_x_ae=_GEN_584[12]; 
  assign entries_barrier_7_io_x_sw=_GEN_584[11]; 
  assign entries_barrier_7_io_x_sx=_GEN_584[10]; 
  assign entries_barrier_7_io_x_sr=_GEN_584[9]; 
  assign entries_barrier_7_io_x_pw=_GEN_584[8]; 
  assign entries_barrier_7_io_x_px=_GEN_584[7]; 
  assign entries_barrier_7_io_x_pr=_GEN_584[6]; 
  assign entries_barrier_7_io_x_ppp=_GEN_584[5]; 
  assign entries_barrier_7_io_x_pal=_GEN_584[4]; 
  assign entries_barrier_7_io_x_paa=_GEN_584[3]; 
  assign entries_barrier_7_io_x_eff=_GEN_584[2]; 
  assign entries_barrier_7_io_x_c=_GEN_584[1]; 
  assign entries_barrier_8_io_x_ppn=superpage_entries_0_data_0[34:15]; 
  assign entries_barrier_8_io_x_u=superpage_entries_0_data_0[14]; 
  assign entries_barrier_8_io_x_ae=superpage_entries_0_data_0[12]; 
  assign entries_barrier_8_io_x_sw=superpage_entries_0_data_0[11]; 
  assign entries_barrier_8_io_x_sx=superpage_entries_0_data_0[10]; 
  assign entries_barrier_8_io_x_sr=superpage_entries_0_data_0[9]; 
  assign entries_barrier_8_io_x_pw=superpage_entries_0_data_0[8]; 
  assign entries_barrier_8_io_x_px=superpage_entries_0_data_0[7]; 
  assign entries_barrier_8_io_x_pr=superpage_entries_0_data_0[6]; 
  assign entries_barrier_8_io_x_ppp=superpage_entries_0_data_0[5]; 
  assign entries_barrier_8_io_x_pal=superpage_entries_0_data_0[4]; 
  assign entries_barrier_8_io_x_paa=superpage_entries_0_data_0[3]; 
  assign entries_barrier_8_io_x_eff=superpage_entries_0_data_0[2]; 
  assign entries_barrier_8_io_x_c=superpage_entries_0_data_0[1]; 
  assign entries_barrier_9_io_x_ppn=superpage_entries_1_data_0[34:15]; 
  assign entries_barrier_9_io_x_u=superpage_entries_1_data_0[14]; 
  assign entries_barrier_9_io_x_ae=superpage_entries_1_data_0[12]; 
  assign entries_barrier_9_io_x_sw=superpage_entries_1_data_0[11]; 
  assign entries_barrier_9_io_x_sx=superpage_entries_1_data_0[10]; 
  assign entries_barrier_9_io_x_sr=superpage_entries_1_data_0[9]; 
  assign entries_barrier_9_io_x_pw=superpage_entries_1_data_0[8]; 
  assign entries_barrier_9_io_x_px=superpage_entries_1_data_0[7]; 
  assign entries_barrier_9_io_x_pr=superpage_entries_1_data_0[6]; 
  assign entries_barrier_9_io_x_ppp=superpage_entries_1_data_0[5]; 
  assign entries_barrier_9_io_x_pal=superpage_entries_1_data_0[4]; 
  assign entries_barrier_9_io_x_paa=superpage_entries_1_data_0[3]; 
  assign entries_barrier_9_io_x_eff=superpage_entries_1_data_0[2]; 
  assign entries_barrier_9_io_x_c=superpage_entries_1_data_0[1]; 
  assign entries_barrier_10_io_x_ppn=superpage_entries_2_data_0[34:15]; 
  assign entries_barrier_10_io_x_u=superpage_entries_2_data_0[14]; 
  assign entries_barrier_10_io_x_ae=superpage_entries_2_data_0[12]; 
  assign entries_barrier_10_io_x_sw=superpage_entries_2_data_0[11]; 
  assign entries_barrier_10_io_x_sx=superpage_entries_2_data_0[10]; 
  assign entries_barrier_10_io_x_sr=superpage_entries_2_data_0[9]; 
  assign entries_barrier_10_io_x_pw=superpage_entries_2_data_0[8]; 
  assign entries_barrier_10_io_x_px=superpage_entries_2_data_0[7]; 
  assign entries_barrier_10_io_x_pr=superpage_entries_2_data_0[6]; 
  assign entries_barrier_10_io_x_ppp=superpage_entries_2_data_0[5]; 
  assign entries_barrier_10_io_x_pal=superpage_entries_2_data_0[4]; 
  assign entries_barrier_10_io_x_paa=superpage_entries_2_data_0[3]; 
  assign entries_barrier_10_io_x_eff=superpage_entries_2_data_0[2]; 
  assign entries_barrier_10_io_x_c=superpage_entries_2_data_0[1]; 
  assign entries_barrier_11_io_x_ppn=superpage_entries_3_data_0[34:15]; 
  assign entries_barrier_11_io_x_u=superpage_entries_3_data_0[14]; 
  assign entries_barrier_11_io_x_ae=superpage_entries_3_data_0[12]; 
  assign entries_barrier_11_io_x_sw=superpage_entries_3_data_0[11]; 
  assign entries_barrier_11_io_x_sx=superpage_entries_3_data_0[10]; 
  assign entries_barrier_11_io_x_sr=superpage_entries_3_data_0[9]; 
  assign entries_barrier_11_io_x_pw=superpage_entries_3_data_0[8]; 
  assign entries_barrier_11_io_x_px=superpage_entries_3_data_0[7]; 
  assign entries_barrier_11_io_x_pr=superpage_entries_3_data_0[6]; 
  assign entries_barrier_11_io_x_ppp=superpage_entries_3_data_0[5]; 
  assign entries_barrier_11_io_x_pal=superpage_entries_3_data_0[4]; 
  assign entries_barrier_11_io_x_paa=superpage_entries_3_data_0[3]; 
  assign entries_barrier_11_io_x_eff=superpage_entries_3_data_0[2]; 
  assign entries_barrier_11_io_x_c=superpage_entries_3_data_0[1]; 
  assign entries_barrier_12_io_x_ppn=special_entry_data_0[34:15]; 
  assign entries_barrier_12_io_x_u=special_entry_data_0[14]; 
  assign entries_barrier_12_io_x_ae=special_entry_data_0[12]; 
  assign entries_barrier_12_io_x_sw=special_entry_data_0[11]; 
  assign entries_barrier_12_io_x_sx=special_entry_data_0[10]; 
  assign entries_barrier_12_io_x_sr=special_entry_data_0[9]; 
  assign entries_barrier_12_io_x_pw=special_entry_data_0[8]; 
  assign entries_barrier_12_io_x_px=special_entry_data_0[7]; 
  assign entries_barrier_12_io_x_pr=special_entry_data_0[6]; 
  assign entries_barrier_12_io_x_ppp=special_entry_data_0[5]; 
  assign entries_barrier_12_io_x_pal=special_entry_data_0[4]; 
  assign entries_barrier_12_io_x_paa=special_entry_data_0[3]; 
  assign entries_barrier_12_io_x_eff=special_entry_data_0[2]; 
  assign entries_barrier_12_io_x_c=special_entry_data_0[1]; 
  assign TLB_cov_read_addr=TLB_state; 
  assign TLB_cov_read_data=TLB_cov[TLB_cov_read_addr]; 
  assign TLB_cov_write_data=1'h1; 
  assign TLB_cov_write_addr=TLB_state; 
  assign TLB_cov_write_mask=1'h1; 
  assign TLB_cov_write_en=1'h1; 
  assign mux_cond_0=sectored_entries_0_6_data_1[0]; 
  assign mux_cond_1=sectored_entries_0_7_data_1[0]; 
  assign mux_cond_2=~sectored_entries_0_2_data_0[13]; 
  assign mux_cond_3=~sectored_entries_0_7_data_1[13]; 
  assign mux_cond_4=sectored_entries_0_7_data_3[0]; 
  assign mux_cond_5=sectored_entries_0_4_data_0[0]; 
  assign mux_cond_6=sectored_entries_0_3_data_3[0]; 
  assign mux_cond_7=sectored_entries_0_2_data_3[0]; 
  assign mux_cond_8=sectored_entries_0_2_data_0[0]; 
  assign mux_cond_9=~sectored_entries_0_6_data_1[13]; 
  assign mux_cond_10=~sectored_entries_0_2_data_2[13]; 
  assign mux_cond_11=~superpage_entries_0_data_0[13]; 
  assign mux_cond_12=sectored_entries_0_3_data_1[0]; 
  assign mux_cond_13=sectored_entries_0_4_data_3[0]; 
  assign mux_cond_14=~sectored_entries_0_3_data_3[13]; 
  assign mux_cond_15=sectored_entries_0_3_data_2[0]; 
  assign mux_cond_16=~sectored_entries_0_4_data_3[13]; 
  assign mux_cond_17=~sectored_entries_0_4_data_0[13]; 
  assign mux_cond_18=~sectored_entries_0_4_data_1[13]; 
  assign mux_cond_19=sectored_entries_0_6_data_0[0]; 
  assign mux_cond_20=sectored_entries_0_5_data_0[0]; 
  assign mux_cond_21=sectored_entries_0_6_data_2[0]; 
  assign mux_cond_22=sectored_entries_0_0_data_3[0]; 
  assign mux_cond_23=~sectored_entries_0_3_data_1[13]; 
  assign mux_cond_24=~sectored_entries_0_7_data_0[13]; 
  assign mux_cond_25=sectored_entries_0_7_data_0[0]; 
  assign mux_cond_26=~sectored_entries_0_7_data_3[13]; 
  assign mux_cond_27=~sectored_entries_0_0_data_3[13]; 
  assign mux_cond_28=~superpage_entries_1_data_0[13]; 
  assign mux_cond_29=~sectored_entries_0_7_data_2[13]; 
  assign mux_cond_30=~sectored_entries_0_6_data_0[13]; 
  assign mux_cond_31=~sectored_entries_0_6_data_3[13]; 
  assign mux_cond_32=sectored_entries_0_2_data_2[0]; 
  assign mux_cond_33=sectored_entries_0_1_data_1[0]; 
  assign mux_cond_34=~sectored_entries_0_2_data_1[13]; 
  assign mux_cond_35=~sectored_entries_0_4_data_2[13]; 
  assign mux_cond_36=~sectored_entries_0_1_data_3[13]; 
  assign mux_cond_37=~sectored_entries_0_0_data_2[13]; 
  assign mux_cond_38=~sectored_entries_0_0_data_0[13]; 
  assign mux_cond_39=~sectored_entries_0_2_data_3[13]; 
  assign mux_cond_40=sectored_entries_0_7_data_2[0]; 
  assign mux_cond_41=sectored_entries_0_0_data_0[0]; 
  assign mux_cond_42=~sectored_entries_0_5_data_0[13]; 
  assign mux_cond_43=sectored_entries_0_4_data_1[0]; 
  assign mux_cond_44=sectored_entries_0_5_data_1[0]; 
  assign mux_cond_45=~sectored_entries_0_5_data_3[13]; 
  assign mux_cond_46=sectored_entries_0_1_data_0[0]; 
  assign mux_cond_47=sectored_entries_0_5_data_3[0]; 
  assign mux_cond_48=~sectored_entries_0_0_data_1[13]; 
  assign mux_cond_49=~special_entry_data_0[13]; 
  assign mux_cond_50=~superpage_entries_2_data_0[13]; 
  assign mux_cond_51=sectored_entries_0_0_data_2[0]; 
  assign mux_cond_52=sectored_entries_0_6_data_3[0]; 
  assign mux_cond_53=~sectored_entries_0_3_data_0[13]; 
  assign mux_cond_54=~sectored_entries_0_1_data_0[13]; 
  assign mux_cond_55=sectored_entries_0_1_data_2[0]; 
  assign mux_cond_56=~sectored_entries_0_5_data_2[13]; 
  assign mux_cond_57=~sectored_entries_0_6_data_2[13]; 
  assign mux_cond_58=sectored_entries_0_1_data_3[0]; 
  assign mux_cond_59=~sectored_entries_0_3_data_2[13]; 
  assign mux_cond_60=~sectored_entries_0_1_data_1[13]; 
  assign mux_cond_61=~sectored_entries_0_1_data_2[13]; 
  assign mux_cond_62=sectored_entries_0_3_data_0[0]; 
  assign mux_cond_63=sectored_entries_0_5_data_2[0]; 
  assign mux_cond_64=sectored_entries_0_0_data_1[0]; 
  assign mux_cond_65=sectored_entries_0_2_data_1[0]; 
  assign mux_cond_66=~sectored_entries_0_5_data_1[13]; 
  assign mux_cond_67=~superpage_entries_3_data_0[13]; 
  assign mux_cond_68=sectored_entries_0_4_data_2[0]; 
  assign r_sectored_hit_shl=r_sectored_hit; 
  assign r_sectored_hit_pad={19'h0,r_sectored_hit_shl}; 
  assign r_sectored_repl_addr_shl={r_sectored_repl_addr,7'h0}; 
  assign r_sectored_repl_addr_pad={10'h0,r_sectored_repl_addr_shl}; 
  assign r_superpage_repl_addr_shl={r_superpage_repl_addr,18'h0}; 
  assign r_superpage_repl_addr_pad=r_superpage_repl_addr_shl; 
  assign special_entry_valid_0_shl={special_entry_valid_0,7'h0}; 
  assign special_entry_valid_0_pad={12'h0,special_entry_valid_0_shl}; 
  assign special_entry_level_shl={special_entry_level,18'h0}; 
  assign special_entry_level_pad=special_entry_level_shl; 
  assign state_shl={state,6'h0}; 
  assign state_pad={12'h0,state_shl}; 
  assign r_sectored_hit_addr_shl={r_sectored_hit_addr,12'h0}; 
  assign r_sectored_hit_addr_pad={5'h0,r_sectored_hit_addr_shl}; 
  assign mux_cond_0_shl={mux_cond_0,5'h0}; 
  assign mux_cond_0_pad={14'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,11'h0}; 
  assign mux_cond_1_pad={8'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl={mux_cond_2,2'h0}; 
  assign mux_cond_2_pad={17'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,12'h0}; 
  assign mux_cond_3_pad={7'h0,mux_cond_3_shl}; 
  assign mux_cond_4_shl={mux_cond_4,11'h0}; 
  assign mux_cond_4_pad={8'h0,mux_cond_4_shl}; 
  assign mux_cond_5_shl={mux_cond_5,1'h0}; 
  assign mux_cond_5_pad={18'h0,mux_cond_5_shl}; 
  assign mux_cond_6_shl={mux_cond_6,13'h0}; 
  assign mux_cond_6_pad={6'h0,mux_cond_6_shl}; 
  assign mux_cond_7_shl={mux_cond_7,6'h0}; 
  assign mux_cond_7_pad={13'h0,mux_cond_7_shl}; 
  assign mux_cond_8_shl={mux_cond_8,4'h0}; 
  assign mux_cond_8_pad={15'h0,mux_cond_8_shl}; 
  assign mux_cond_9_shl={mux_cond_9,17'h0}; 
  assign mux_cond_9_pad={2'h0,mux_cond_9_shl}; 
  assign mux_cond_10_shl={mux_cond_10,5'h0}; 
  assign mux_cond_10_pad={14'h0,mux_cond_10_shl}; 
  assign mux_cond_11_shl={mux_cond_11,9'h0}; 
  assign mux_cond_11_pad={10'h0,mux_cond_11_shl}; 
  assign mux_cond_12_shl={mux_cond_12,1'h0}; 
  assign mux_cond_12_pad={18'h0,mux_cond_12_shl}; 
  assign mux_cond_13_shl={mux_cond_13,9'h0}; 
  assign mux_cond_13_pad={10'h0,mux_cond_13_shl}; 
  assign mux_cond_14_shl={mux_cond_14,12'h0}; 
  assign mux_cond_14_pad={7'h0,mux_cond_14_shl}; 
  assign mux_cond_15_shl={mux_cond_15,7'h0}; 
  assign mux_cond_15_pad={12'h0,mux_cond_15_shl}; 
  assign mux_cond_16_shl={mux_cond_16,6'h0}; 
  assign mux_cond_16_pad={13'h0,mux_cond_16_shl}; 
  assign mux_cond_17_shl={mux_cond_17,7'h0}; 
  assign mux_cond_17_pad={12'h0,mux_cond_17_shl}; 
  assign mux_cond_18_shl={mux_cond_18,16'h0}; 
  assign mux_cond_18_pad={3'h0,mux_cond_18_shl}; 
  assign mux_cond_19_shl={mux_cond_19,8'h0}; 
  assign mux_cond_19_pad={11'h0,mux_cond_19_shl}; 
  assign mux_cond_20_shl={mux_cond_20,1'h0}; 
  assign mux_cond_20_pad={18'h0,mux_cond_20_shl}; 
  assign mux_cond_21_shl={mux_cond_21,5'h0}; 
  assign mux_cond_21_pad={14'h0,mux_cond_21_shl}; 
  assign mux_cond_22_shl={mux_cond_22,11'h0}; 
  assign mux_cond_22_pad={8'h0,mux_cond_22_shl}; 
  assign mux_cond_23_shl={mux_cond_23,2'h0}; 
  assign mux_cond_23_pad={17'h0,mux_cond_23_shl}; 
  assign mux_cond_24_shl={mux_cond_24,14'h0}; 
  assign mux_cond_24_pad={5'h0,mux_cond_24_shl}; 
  assign mux_cond_25_shl={mux_cond_25,3'h0}; 
  assign mux_cond_25_pad={16'h0,mux_cond_25_shl}; 
  assign mux_cond_26_shl={mux_cond_26,11'h0}; 
  assign mux_cond_26_pad={8'h0,mux_cond_26_shl}; 
  assign mux_cond_27_shl=mux_cond_27; 
  assign mux_cond_27_pad={19'h0,mux_cond_27_shl}; 
  assign mux_cond_28_shl={mux_cond_28,18'h0}; 
  assign mux_cond_28_pad={1'h0,mux_cond_28_shl}; 
  assign mux_cond_29_shl={mux_cond_29,14'h0}; 
  assign mux_cond_29_pad={5'h0,mux_cond_29_shl}; 
  assign mux_cond_30_shl={mux_cond_30,8'h0}; 
  assign mux_cond_30_pad={11'h0,mux_cond_30_shl}; 
  assign mux_cond_31_shl={mux_cond_31,3'h0}; 
  assign mux_cond_31_pad={16'h0,mux_cond_31_shl}; 
  assign mux_cond_32_shl={mux_cond_32,2'h0}; 
  assign mux_cond_32_pad={17'h0,mux_cond_32_shl}; 
  assign mux_cond_33_shl=mux_cond_33; 
  assign mux_cond_33_pad={19'h0,mux_cond_33_shl}; 
  assign mux_cond_34_shl={mux_cond_34,7'h0}; 
  assign mux_cond_34_pad={12'h0,mux_cond_34_shl}; 
  assign mux_cond_35_shl={mux_cond_35,4'h0}; 
  assign mux_cond_35_pad={15'h0,mux_cond_35_shl}; 
  assign mux_cond_36_shl={mux_cond_36,3'h0}; 
  assign mux_cond_36_pad={16'h0,mux_cond_36_shl}; 
  assign mux_cond_37_shl={mux_cond_37,4'h0}; 
  assign mux_cond_37_pad={15'h0,mux_cond_37_shl}; 
  assign mux_cond_38_shl={mux_cond_38,12'h0}; 
  assign mux_cond_38_pad={7'h0,mux_cond_38_shl}; 
  assign mux_cond_39_shl={mux_cond_39,9'h0}; 
  assign mux_cond_39_pad={10'h0,mux_cond_39_shl}; 
  assign mux_cond_40_shl=mux_cond_40; 
  assign mux_cond_40_pad={19'h0,mux_cond_40_shl}; 
  assign mux_cond_41_shl={mux_cond_41,16'h0}; 
  assign mux_cond_41_pad={3'h0,mux_cond_41_shl}; 
  assign mux_cond_42_shl={mux_cond_42,4'h0}; 
  assign mux_cond_42_pad={15'h0,mux_cond_42_shl}; 
  assign mux_cond_43_shl={mux_cond_43,18'h0}; 
  assign mux_cond_43_pad={1'h0,mux_cond_43_shl}; 
  assign mux_cond_44_shl={mux_cond_44,8'h0}; 
  assign mux_cond_44_pad={11'h0,mux_cond_44_shl}; 
  assign mux_cond_45_shl={mux_cond_45,17'h0}; 
  assign mux_cond_45_pad={2'h0,mux_cond_45_shl}; 
  assign mux_cond_46_shl={mux_cond_46,5'h0}; 
  assign mux_cond_46_pad={14'h0,mux_cond_46_shl}; 
  assign mux_cond_47_shl={mux_cond_47,8'h0}; 
  assign mux_cond_47_pad={11'h0,mux_cond_47_shl}; 
  assign mux_cond_48_shl={mux_cond_48,7'h0}; 
  assign mux_cond_48_pad={12'h0,mux_cond_48_shl}; 
  assign mux_cond_49_shl={mux_cond_49,16'h0}; 
  assign mux_cond_49_pad={3'h0,mux_cond_49_shl}; 
  assign mux_cond_50_shl={mux_cond_50,8'h0}; 
  assign mux_cond_50_pad={11'h0,mux_cond_50_shl}; 
  assign mux_cond_51_shl={mux_cond_51,4'h0}; 
  assign mux_cond_51_pad={15'h0,mux_cond_51_shl}; 
  assign mux_cond_52_shl={mux_cond_52,3'h0}; 
  assign mux_cond_52_pad={16'h0,mux_cond_52_shl}; 
  assign mux_cond_53_shl={mux_cond_53,6'h0}; 
  assign mux_cond_53_pad={13'h0,mux_cond_53_shl}; 
  assign mux_cond_54_shl={mux_cond_54,18'h0}; 
  assign mux_cond_54_pad={1'h0,mux_cond_54_shl}; 
  assign mux_cond_55_shl={mux_cond_55,15'h0}; 
  assign mux_cond_55_pad={4'h0,mux_cond_55_shl}; 
  assign mux_cond_56_shl={mux_cond_56,16'h0}; 
  assign mux_cond_56_pad={3'h0,mux_cond_56_shl}; 
  assign mux_cond_57_shl={mux_cond_57,7'h0}; 
  assign mux_cond_57_pad={12'h0,mux_cond_57_shl}; 
  assign mux_cond_58_shl={mux_cond_58,11'h0}; 
  assign mux_cond_58_pad={8'h0,mux_cond_58_shl}; 
  assign mux_cond_59_shl={mux_cond_59,14'h0}; 
  assign mux_cond_59_pad={5'h0,mux_cond_59_shl}; 
  assign mux_cond_60_shl={mux_cond_60,13'h0}; 
  assign mux_cond_60_pad={6'h0,mux_cond_60_shl}; 
  assign mux_cond_61_shl={mux_cond_61,8'h0}; 
  assign mux_cond_61_pad={11'h0,mux_cond_61_shl}; 
  assign mux_cond_62_shl={mux_cond_62,7'h0}; 
  assign mux_cond_62_pad={12'h0,mux_cond_62_shl}; 
  assign mux_cond_63_shl={mux_cond_63,6'h0}; 
  assign mux_cond_63_pad={13'h0,mux_cond_63_shl}; 
  assign mux_cond_64_shl={mux_cond_64,19'h0}; 
  assign mux_cond_64_pad=mux_cond_64_shl; 
  assign mux_cond_65_shl={mux_cond_65,11'h0}; 
  assign mux_cond_65_pad={8'h0,mux_cond_65_shl}; 
  assign mux_cond_66_shl={mux_cond_66,6'h0}; 
  assign mux_cond_66_pad={13'h0,mux_cond_66_shl}; 
  assign mux_cond_67_shl={mux_cond_67,10'h0}; 
  assign mux_cond_67_pad={9'h0,mux_cond_67_shl}; 
  assign mux_cond_68_shl={mux_cond_68,13'h0}; 
  assign mux_cond_68_pad={6'h0,mux_cond_68_shl}; 
  assign sectored_entries_0_0_valid_3_shl={sectored_entries_0_0_valid_3,16'h0}; 
  assign sectored_entries_0_0_valid_3_pad={3'h0,sectored_entries_0_0_valid_3_shl}; 
  assign sectored_entries_0_0_valid_2_shl={sectored_entries_0_0_valid_2,8'h0}; 
  assign sectored_entries_0_0_valid_2_pad={11'h0,sectored_entries_0_0_valid_2_shl}; 
  assign sectored_entries_0_2_valid_0_shl={sectored_entries_0_2_valid_0,8'h0}; 
  assign sectored_entries_0_2_valid_0_pad={11'h0,sectored_entries_0_2_valid_0_shl}; 
  assign sectored_entries_0_3_valid_0_shl={sectored_entries_0_3_valid_0,8'h0}; 
  assign sectored_entries_0_3_valid_0_pad={11'h0,sectored_entries_0_3_valid_0_shl}; 
  assign superpage_entries_2_level_shl=superpage_entries_2_level; 
  assign superpage_entries_2_level_pad={18'h0,superpage_entries_2_level_shl}; 
  assign sectored_entries_0_7_valid_1_shl=sectored_entries_0_7_valid_1; 
  assign sectored_entries_0_7_valid_1_pad={19'h0,sectored_entries_0_7_valid_1_shl}; 
  assign sectored_entries_0_4_valid_0_shl={sectored_entries_0_4_valid_0,8'h0}; 
  assign sectored_entries_0_4_valid_0_pad={11'h0,sectored_entries_0_4_valid_0_shl}; 
  assign sectored_entries_0_1_valid_3_shl={sectored_entries_0_1_valid_3,16'h0}; 
  assign sectored_entries_0_1_valid_3_pad={3'h0,sectored_entries_0_1_valid_3_shl}; 
  assign sectored_entries_0_1_valid_1_shl=sectored_entries_0_1_valid_1; 
  assign sectored_entries_0_1_valid_1_pad={19'h0,sectored_entries_0_1_valid_1_shl}; 
  assign sectored_entries_0_2_valid_3_shl={sectored_entries_0_2_valid_3,16'h0}; 
  assign sectored_entries_0_2_valid_3_pad={3'h0,sectored_entries_0_2_valid_3_shl}; 
  assign sectored_entries_0_2_valid_1_shl=sectored_entries_0_2_valid_1; 
  assign sectored_entries_0_2_valid_1_pad={19'h0,sectored_entries_0_2_valid_1_shl}; 
  assign superpage_entries_1_valid_0_shl={superpage_entries_1_valid_0,11'h0}; 
  assign superpage_entries_1_valid_0_pad={8'h0,superpage_entries_1_valid_0_shl}; 
  assign sectored_entries_0_7_valid_0_shl={sectored_entries_0_7_valid_0,8'h0}; 
  assign sectored_entries_0_7_valid_0_pad={11'h0,sectored_entries_0_7_valid_0_shl}; 
  assign superpage_entries_3_valid_0_shl={superpage_entries_3_valid_0,11'h0}; 
  assign superpage_entries_3_valid_0_pad={8'h0,superpage_entries_3_valid_0_shl}; 
  assign sectored_entries_0_5_valid_3_shl={sectored_entries_0_5_valid_3,16'h0}; 
  assign sectored_entries_0_5_valid_3_pad={3'h0,sectored_entries_0_5_valid_3_shl}; 
  assign sectored_entries_0_5_valid_1_shl=sectored_entries_0_5_valid_1; 
  assign sectored_entries_0_5_valid_1_pad={19'h0,sectored_entries_0_5_valid_1_shl}; 
  assign sectored_entries_0_4_valid_3_shl={sectored_entries_0_4_valid_3,16'h0}; 
  assign sectored_entries_0_4_valid_3_pad={3'h0,sectored_entries_0_4_valid_3_shl}; 
  assign sectored_entries_0_5_valid_2_shl={sectored_entries_0_5_valid_2,8'h0}; 
  assign sectored_entries_0_5_valid_2_pad={11'h0,sectored_entries_0_5_valid_2_shl}; 
  assign sectored_entries_0_1_valid_2_shl={sectored_entries_0_1_valid_2,8'h0}; 
  assign sectored_entries_0_1_valid_2_pad={11'h0,sectored_entries_0_1_valid_2_shl}; 
  assign sectored_entries_0_3_valid_1_shl=sectored_entries_0_3_valid_1; 
  assign sectored_entries_0_3_valid_1_pad={19'h0,sectored_entries_0_3_valid_1_shl}; 
  assign sectored_entries_0_1_valid_0_shl={sectored_entries_0_1_valid_0,8'h0}; 
  assign sectored_entries_0_1_valid_0_pad={11'h0,sectored_entries_0_1_valid_0_shl}; 
  assign sectored_entries_0_4_valid_2_shl={sectored_entries_0_4_valid_2,8'h0}; 
  assign sectored_entries_0_4_valid_2_pad={11'h0,sectored_entries_0_4_valid_2_shl}; 
  assign sectored_entries_0_4_valid_1_shl=sectored_entries_0_4_valid_1; 
  assign sectored_entries_0_4_valid_1_pad={19'h0,sectored_entries_0_4_valid_1_shl}; 
  assign superpage_entries_3_level_shl=superpage_entries_3_level; 
  assign superpage_entries_3_level_pad={18'h0,superpage_entries_3_level_shl}; 
  assign sectored_entries_0_0_valid_1_shl=sectored_entries_0_0_valid_1; 
  assign sectored_entries_0_0_valid_1_pad={19'h0,sectored_entries_0_0_valid_1_shl}; 
  assign sectored_entries_0_3_valid_2_shl={sectored_entries_0_3_valid_2,8'h0}; 
  assign sectored_entries_0_3_valid_2_pad={11'h0,sectored_entries_0_3_valid_2_shl}; 
  assign sectored_entries_0_6_valid_1_shl=sectored_entries_0_6_valid_1; 
  assign sectored_entries_0_6_valid_1_pad={19'h0,sectored_entries_0_6_valid_1_shl}; 
  assign sectored_entries_0_7_valid_3_shl={sectored_entries_0_7_valid_3,16'h0}; 
  assign sectored_entries_0_7_valid_3_pad={3'h0,sectored_entries_0_7_valid_3_shl}; 
  assign sectored_entries_0_3_valid_3_shl={sectored_entries_0_3_valid_3,16'h0}; 
  assign sectored_entries_0_3_valid_3_pad={3'h0,sectored_entries_0_3_valid_3_shl}; 
  assign sectored_entries_0_0_valid_0_shl={sectored_entries_0_0_valid_0,8'h0}; 
  assign sectored_entries_0_0_valid_0_pad={11'h0,sectored_entries_0_0_valid_0_shl}; 
  assign superpage_entries_0_valid_0_shl={superpage_entries_0_valid_0,11'h0}; 
  assign superpage_entries_0_valid_0_pad={8'h0,superpage_entries_0_valid_0_shl}; 
  assign sectored_entries_0_2_valid_2_shl={sectored_entries_0_2_valid_2,8'h0}; 
  assign sectored_entries_0_2_valid_2_pad={11'h0,sectored_entries_0_2_valid_2_shl}; 
  assign sectored_entries_0_6_valid_2_shl={sectored_entries_0_6_valid_2,8'h0}; 
  assign sectored_entries_0_6_valid_2_pad={11'h0,sectored_entries_0_6_valid_2_shl}; 
  assign superpage_entries_2_valid_0_shl={superpage_entries_2_valid_0,11'h0}; 
  assign superpage_entries_2_valid_0_pad={8'h0,superpage_entries_2_valid_0_shl}; 
  assign sectored_entries_0_6_valid_3_shl={sectored_entries_0_6_valid_3,16'h0}; 
  assign sectored_entries_0_6_valid_3_pad={3'h0,sectored_entries_0_6_valid_3_shl}; 
  assign sectored_entries_0_6_valid_0_shl={sectored_entries_0_6_valid_0,8'h0}; 
  assign sectored_entries_0_6_valid_0_pad={11'h0,sectored_entries_0_6_valid_0_shl}; 
  assign sectored_entries_0_7_valid_2_shl={sectored_entries_0_7_valid_2,8'h0}; 
  assign sectored_entries_0_7_valid_2_pad={11'h0,sectored_entries_0_7_valid_2_shl}; 
  assign superpage_entries_0_level_shl=superpage_entries_0_level; 
  assign superpage_entries_0_level_pad={18'h0,superpage_entries_0_level_shl}; 
  assign superpage_entries_1_level_shl=superpage_entries_1_level; 
  assign superpage_entries_1_level_pad={18'h0,superpage_entries_1_level_shl}; 
  assign sectored_entries_0_5_valid_0_shl={sectored_entries_0_5_valid_0,8'h0}; 
  assign sectored_entries_0_5_valid_0_pad={11'h0,sectored_entries_0_5_valid_0_shl}; 
  assign TLB_xor64=r_sectored_repl_addr_pad^r_superpage_repl_addr_pad; 
  assign TLB_xor31=r_sectored_hit_pad^TLB_xor64; 
  assign TLB_xor65=special_entry_valid_0_pad^special_entry_level_pad; 
  assign TLB_xor66=state_pad^r_sectored_hit_addr_pad; 
  assign TLB_xor32=TLB_xor65^TLB_xor66; 
  assign TLB_xor15=TLB_xor31^TLB_xor32; 
  assign TLB_xor68=mux_cond_1_pad^mux_cond_2_pad; 
  assign TLB_xor33=mux_cond_0_pad^TLB_xor68; 
  assign TLB_xor69=mux_cond_3_pad^mux_cond_4_pad; 
  assign TLB_xor70=mux_cond_5_pad^mux_cond_6_pad; 
  assign TLB_xor34=TLB_xor69^TLB_xor70; 
  assign TLB_xor16=TLB_xor33^TLB_xor34; 
  assign TLB_xor7=TLB_xor15^TLB_xor16; 
  assign TLB_xor72=mux_cond_8_pad^mux_cond_9_pad; 
  assign TLB_xor35=mux_cond_7_pad^TLB_xor72; 
  assign TLB_xor73=mux_cond_10_pad^mux_cond_11_pad; 
  assign TLB_xor74=mux_cond_12_pad^mux_cond_13_pad; 
  assign TLB_xor36=TLB_xor73^TLB_xor74; 
  assign TLB_xor17=TLB_xor35^TLB_xor36; 
  assign TLB_xor75=mux_cond_14_pad^mux_cond_15_pad; 
  assign TLB_xor76=mux_cond_16_pad^mux_cond_17_pad; 
  assign TLB_xor37=TLB_xor75^TLB_xor76; 
  assign TLB_xor77=mux_cond_18_pad^mux_cond_19_pad; 
  assign TLB_xor78=mux_cond_20_pad^mux_cond_21_pad; 
  assign TLB_xor38=TLB_xor77^TLB_xor78; 
  assign TLB_xor18=TLB_xor37^TLB_xor38; 
  assign TLB_xor8=TLB_xor17^TLB_xor18; 
  assign TLB_xor3=TLB_xor7^TLB_xor8; 
  assign TLB_xor80=mux_cond_23_pad^mux_cond_24_pad; 
  assign TLB_xor39=mux_cond_22_pad^TLB_xor80; 
  assign TLB_xor81=mux_cond_25_pad^mux_cond_26_pad; 
  assign TLB_xor82=mux_cond_27_pad^mux_cond_28_pad; 
  assign TLB_xor40=TLB_xor81^TLB_xor82; 
  assign TLB_xor19=TLB_xor39^TLB_xor40; 
  assign TLB_xor84=mux_cond_30_pad^mux_cond_31_pad; 
  assign TLB_xor41=mux_cond_29_pad^TLB_xor84; 
  assign TLB_xor85=mux_cond_32_pad^mux_cond_33_pad; 
  assign TLB_xor86=mux_cond_34_pad^mux_cond_35_pad; 
  assign TLB_xor42=TLB_xor85^TLB_xor86; 
  assign TLB_xor20=TLB_xor41^TLB_xor42; 
  assign TLB_xor9=TLB_xor19^TLB_xor20; 
  assign TLB_xor88=mux_cond_37_pad^mux_cond_38_pad; 
  assign TLB_xor43=mux_cond_36_pad^TLB_xor88; 
  assign TLB_xor89=mux_cond_39_pad^mux_cond_40_pad; 
  assign TLB_xor90=mux_cond_41_pad^mux_cond_42_pad; 
  assign TLB_xor44=TLB_xor89^TLB_xor90; 
  assign TLB_xor21=TLB_xor43^TLB_xor44; 
  assign TLB_xor91=mux_cond_43_pad^mux_cond_44_pad; 
  assign TLB_xor92=mux_cond_45_pad^mux_cond_46_pad; 
  assign TLB_xor45=TLB_xor91^TLB_xor92; 
  assign TLB_xor93=mux_cond_47_pad^mux_cond_48_pad; 
  assign TLB_xor94=mux_cond_49_pad^mux_cond_50_pad; 
  assign TLB_xor46=TLB_xor93^TLB_xor94; 
  assign TLB_xor22=TLB_xor45^TLB_xor46; 
  assign TLB_xor10=TLB_xor21^TLB_xor22; 
  assign TLB_xor4=TLB_xor9^TLB_xor10; 
  assign TLB_xor1=TLB_xor3^TLB_xor4; 
  assign TLB_xor96=mux_cond_52_pad^mux_cond_53_pad; 
  assign TLB_xor47=mux_cond_51_pad^TLB_xor96; 
  assign TLB_xor97=mux_cond_54_pad^mux_cond_55_pad; 
  assign TLB_xor98=mux_cond_56_pad^mux_cond_57_pad; 
  assign TLB_xor48=TLB_xor97^TLB_xor98; 
  assign TLB_xor23=TLB_xor47^TLB_xor48; 
  assign TLB_xor100=mux_cond_59_pad^mux_cond_60_pad; 
  assign TLB_xor49=mux_cond_58_pad^TLB_xor100; 
  assign TLB_xor101=mux_cond_61_pad^mux_cond_62_pad; 
  assign TLB_xor102=mux_cond_63_pad^mux_cond_64_pad; 
  assign TLB_xor50=TLB_xor101^TLB_xor102; 
  assign TLB_xor24=TLB_xor49^TLB_xor50; 
  assign TLB_xor11=TLB_xor23^TLB_xor24; 
  assign TLB_xor104=mux_cond_66_pad^mux_cond_67_pad; 
  assign TLB_xor51=mux_cond_65_pad^TLB_xor104; 
  assign TLB_xor105=mux_cond_68_pad^sectored_entries_0_0_valid_3_pad; 
  assign TLB_xor106=sectored_entries_0_0_valid_2_pad^sectored_entries_0_2_valid_0_pad; 
  assign TLB_xor52=TLB_xor105^TLB_xor106; 
  assign TLB_xor25=TLB_xor51^TLB_xor52; 
  assign TLB_xor107=sectored_entries_0_3_valid_0_pad^superpage_entries_2_level_pad; 
  assign TLB_xor108=sectored_entries_0_7_valid_1_pad^sectored_entries_0_4_valid_0_pad; 
  assign TLB_xor53=TLB_xor107^TLB_xor108; 
  assign TLB_xor109=sectored_entries_0_1_valid_3_pad^sectored_entries_0_1_valid_1_pad; 
  assign TLB_xor110=sectored_entries_0_2_valid_3_pad^sectored_entries_0_2_valid_1_pad; 
  assign TLB_xor54=TLB_xor109^TLB_xor110; 
  assign TLB_xor26=TLB_xor53^TLB_xor54; 
  assign TLB_xor12=TLB_xor25^TLB_xor26; 
  assign TLB_xor5=TLB_xor11^TLB_xor12; 
  assign TLB_xor112=sectored_entries_0_7_valid_0_pad^superpage_entries_3_valid_0_pad; 
  assign TLB_xor55=superpage_entries_1_valid_0_pad^TLB_xor112; 
  assign TLB_xor113=sectored_entries_0_5_valid_3_pad^sectored_entries_0_5_valid_1_pad; 
  assign TLB_xor114=sectored_entries_0_4_valid_3_pad^sectored_entries_0_5_valid_2_pad; 
  assign TLB_xor56=TLB_xor113^TLB_xor114; 
  assign TLB_xor27=TLB_xor55^TLB_xor56; 
  assign TLB_xor116=sectored_entries_0_3_valid_1_pad^sectored_entries_0_1_valid_0_pad; 
  assign TLB_xor57=sectored_entries_0_1_valid_2_pad^TLB_xor116; 
  assign TLB_xor117=sectored_entries_0_4_valid_2_pad^sectored_entries_0_4_valid_1_pad; 
  assign TLB_xor118=superpage_entries_3_level_pad^sectored_entries_0_0_valid_1_pad; 
  assign TLB_xor58=TLB_xor117^TLB_xor118; 
  assign TLB_xor28=TLB_xor57^TLB_xor58; 
  assign TLB_xor13=TLB_xor27^TLB_xor28; 
  assign TLB_xor120=sectored_entries_0_6_valid_1_pad^sectored_entries_0_7_valid_3_pad; 
  assign TLB_xor59=sectored_entries_0_3_valid_2_pad^TLB_xor120; 
  assign TLB_xor121=sectored_entries_0_3_valid_3_pad^sectored_entries_0_0_valid_0_pad; 
  assign TLB_xor122=superpage_entries_0_valid_0_pad^sectored_entries_0_2_valid_2_pad; 
  assign TLB_xor60=TLB_xor121^TLB_xor122; 
  assign TLB_xor29=TLB_xor59^TLB_xor60; 
  assign TLB_xor123=sectored_entries_0_6_valid_2_pad^superpage_entries_2_valid_0_pad; 
  assign TLB_xor124=sectored_entries_0_6_valid_3_pad^sectored_entries_0_6_valid_0_pad; 
  assign TLB_xor61=TLB_xor123^TLB_xor124; 
  assign TLB_xor125=sectored_entries_0_7_valid_2_pad^superpage_entries_0_level_pad; 
  assign TLB_xor126=superpage_entries_1_level_pad^sectored_entries_0_5_valid_0_pad; 
  assign TLB_xor62=TLB_xor125^TLB_xor126; 
  assign TLB_xor30=TLB_xor61^TLB_xor62; 
  assign TLB_xor14=TLB_xor29^TLB_xor30; 
  assign TLB_xor6=TLB_xor13^TLB_xor14; 
  assign TLB_xor2=TLB_xor5^TLB_xor6; 
  assign TLB_xor0=TLB_xor1^TLB_xor2; 
  assign mpu_ppn_barrier_sum=TLB_covSum+mpu_ppn_barrier_io_covSum; 
  assign entries_barrier_10_sum=mpu_ppn_barrier_sum+entries_barrier_10_io_covSum; 
  assign entries_barrier_9_sum=entries_barrier_10_sum+entries_barrier_9_io_covSum; 
  assign entries_barrier_7_sum=entries_barrier_9_sum+entries_barrier_7_io_covSum; 
  assign entries_barrier_sum=entries_barrier_7_sum+entries_barrier_io_covSum; 
  assign entries_barrier_6_sum=entries_barrier_sum+entries_barrier_6_io_covSum; 
  assign entries_barrier_12_sum=entries_barrier_6_sum+entries_barrier_12_io_covSum; 
  assign entries_barrier_1_sum=entries_barrier_12_sum+entries_barrier_1_io_covSum; 
  assign entries_barrier_11_sum=entries_barrier_1_sum+entries_barrier_11_io_covSum; 
  assign entries_barrier_8_sum=entries_barrier_11_sum+entries_barrier_8_io_covSum; 
  assign pmp_sum=entries_barrier_8_sum+pmp_io_covSum; 
  assign entries_barrier_2_sum=pmp_sum+entries_barrier_2_io_covSum; 
  assign entries_barrier_4_sum=entries_barrier_2_sum+entries_barrier_4_io_covSum; 
  assign entries_barrier_5_sum=entries_barrier_4_sum+entries_barrier_5_io_covSum; 
  assign entries_barrier_3_sum=entries_barrier_5_sum+entries_barrier_3_io_covSum; 
  assign io_covSum=entries_barrier_3_sum; 
  assign stopEn0=io_sfence_valid&~_T_51; 
  assign entries_barrier_12_metaAssert_wire=entries_barrier_12_metaAssert; 
  assign entries_barrier_metaAssert_wire=entries_barrier_metaAssert; 
  assign entries_barrier_10_metaAssert_wire=entries_barrier_10_metaAssert; 
  assign entries_barrier_5_metaAssert_wire=entries_barrier_5_metaAssert; 
  assign entries_barrier_11_metaAssert_wire=entries_barrier_11_metaAssert; 
  assign entries_barrier_9_metaAssert_wire=entries_barrier_9_metaAssert; 
  assign entries_barrier_8_metaAssert_wire=entries_barrier_8_metaAssert; 
  assign entries_barrier_1_metaAssert_wire=entries_barrier_1_metaAssert; 
  assign mpu_ppn_barrier_metaAssert_wire=mpu_ppn_barrier_metaAssert; 
  assign entries_barrier_4_metaAssert_wire=entries_barrier_4_metaAssert; 
  assign entries_barrier_6_metaAssert_wire=entries_barrier_6_metaAssert; 
  assign entries_barrier_3_metaAssert_wire=entries_barrier_3_metaAssert; 
  assign pmp_metaAssert_wire=pmp_metaAssert; 
  assign entries_barrier_7_metaAssert_wire=entries_barrier_7_metaAssert; 
  assign entries_barrier_2_metaAssert_wire=entries_barrier_2_metaAssert; 
  assign TLB_or7=stopEn0|entries_barrier_6_metaAssert_wire; 
  assign TLB_or8=entries_barrier_10_metaAssert_wire|entries_barrier_7_metaAssert_wire; 
  assign TLB_or3=TLB_or7|TLB_or8; 
  assign TLB_or9=entries_barrier_4_metaAssert_wire|entries_barrier_11_metaAssert_wire; 
  assign TLB_or10=entries_barrier_8_metaAssert_wire|entries_barrier_9_metaAssert_wire; 
  assign TLB_or4=TLB_or9|TLB_or10; 
  assign TLB_or1=TLB_or3|TLB_or4; 
  assign TLB_or11=entries_barrier_metaAssert_wire|entries_barrier_3_metaAssert_wire; 
  assign TLB_or12=pmp_metaAssert_wire|mpu_ppn_barrier_metaAssert_wire; 
  assign TLB_or5=TLB_or11|TLB_or12; 
  assign TLB_or13=entries_barrier_12_metaAssert_wire|entries_barrier_5_metaAssert_wire; 
  assign TLB_or14=entries_barrier_2_metaAssert_wire|entries_barrier_1_metaAssert_wire; 
  assign TLB_or6=TLB_or13|TLB_or14; 
  assign TLB_or2=TLB_or5|TLB_or6; 
  assign TLB_or0=TLB_or1|TLB_or2; 
  assign metaAssert=TLB_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              sectored_entries_0_0_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                sectored_entries_0_0_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_0_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_0_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_0_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_0_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_0[0])
                                 begin 
                                   sectored_entries_0_0_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_0 <=_GEN_53;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=_GEN_53;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=_GEN_53;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_0 <=_GEN_53;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_0 <=_GEN_621;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_0 <=_GEN_473;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_1[0])
                                 begin 
                                   sectored_entries_0_0_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_1 <=_GEN_54;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=_GEN_54;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=_GEN_54;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_1 <=_GEN_54;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_1 <=_GEN_622;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_1 <=_GEN_474;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_2[0])
                                 begin 
                                   sectored_entries_0_0_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_2 <=_GEN_55;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=_GEN_55;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=_GEN_55;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_2 <=_GEN_55;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_2 <=_GEN_623;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_2 <=_GEN_475;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_3[0])
                                 begin 
                                   sectored_entries_0_0_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_3 <=_GEN_56;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=_GEN_56;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=_GEN_56;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_3 <=_GEN_56;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_3 <=_GEN_624;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_3 <=_GEN_476;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                sectored_entries_0_1_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_1_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_1_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_1_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_1_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_0[0])
                                 begin 
                                   sectored_entries_0_1_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_0 <=_GEN_79;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=_GEN_79;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=_GEN_79;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_0 <=_GEN_79;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_0 <=_GEN_649;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_0 <=_GEN_483;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_1[0])
                                 begin 
                                   sectored_entries_0_1_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_1 <=_GEN_80;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=_GEN_80;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=_GEN_80;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_1 <=_GEN_80;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_1 <=_GEN_650;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_1 <=_GEN_484;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_2[0])
                                 begin 
                                   sectored_entries_0_1_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_2 <=_GEN_81;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=_GEN_81;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=_GEN_81;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_2 <=_GEN_81;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_2 <=_GEN_651;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_2 <=_GEN_485;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_3[0])
                                 begin 
                                   sectored_entries_0_1_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_3 <=_GEN_82;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=_GEN_82;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=_GEN_82;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_3 <=_GEN_82;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_3 <=_GEN_652;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_3 <=_GEN_486;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                sectored_entries_0_2_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_2_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_2_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_2_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_2_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_0[0])
                                 begin 
                                   sectored_entries_0_2_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_0 <=_GEN_105;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=_GEN_105;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=_GEN_105;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_0 <=_GEN_105;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_0 <=_GEN_677;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_0 <=_GEN_493;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_1[0])
                                 begin 
                                   sectored_entries_0_2_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_1 <=_GEN_106;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=_GEN_106;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=_GEN_106;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_1 <=_GEN_106;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_1 <=_GEN_678;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_1 <=_GEN_494;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_2[0])
                                 begin 
                                   sectored_entries_0_2_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_2 <=_GEN_107;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=_GEN_107;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=_GEN_107;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_2 <=_GEN_107;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_2 <=_GEN_679;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_2 <=_GEN_495;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_3[0])
                                 begin 
                                   sectored_entries_0_2_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_3 <=_GEN_108;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=_GEN_108;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=_GEN_108;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_3 <=_GEN_108;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_3 <=_GEN_680;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_3 <=_GEN_496;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                sectored_entries_0_3_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_3_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_3_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_3_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_3_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_0[0])
                                 begin 
                                   sectored_entries_0_3_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_0 <=_GEN_131;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=_GEN_131;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=_GEN_131;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_0 <=_GEN_131;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_0 <=_GEN_705;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_0 <=_GEN_503;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_1[0])
                                 begin 
                                   sectored_entries_0_3_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_1 <=_GEN_132;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=_GEN_132;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=_GEN_132;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_1 <=_GEN_132;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_1 <=_GEN_706;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_1 <=_GEN_504;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_2[0])
                                 begin 
                                   sectored_entries_0_3_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_2 <=_GEN_133;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=_GEN_133;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=_GEN_133;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_2 <=_GEN_133;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_2 <=_GEN_707;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_2 <=_GEN_505;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_3[0])
                                 begin 
                                   sectored_entries_0_3_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_3 <=_GEN_134;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=_GEN_134;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=_GEN_134;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_3 <=_GEN_134;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_3 <=_GEN_708;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_3 <=_GEN_506;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                sectored_entries_0_4_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_4_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_4_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_4_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_4_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_0[0])
                                 begin 
                                   sectored_entries_0_4_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_0 <=_GEN_157;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=_GEN_157;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=_GEN_157;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_0 <=_GEN_157;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_0 <=_GEN_733;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_0 <=_GEN_513;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_1[0])
                                 begin 
                                   sectored_entries_0_4_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_1 <=_GEN_158;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=_GEN_158;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=_GEN_158;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_1 <=_GEN_158;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_1 <=_GEN_734;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_1 <=_GEN_514;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_2[0])
                                 begin 
                                   sectored_entries_0_4_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_2 <=_GEN_159;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=_GEN_159;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=_GEN_159;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_2 <=_GEN_159;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_2 <=_GEN_735;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_2 <=_GEN_515;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_3[0])
                                 begin 
                                   sectored_entries_0_4_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_3 <=_GEN_160;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=_GEN_160;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=_GEN_160;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_3 <=_GEN_160;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_3 <=_GEN_736;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_3 <=_GEN_516;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                sectored_entries_0_5_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_5_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_5_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_5_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_5_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_0[0])
                                 begin 
                                   sectored_entries_0_5_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_0 <=_GEN_183;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=_GEN_183;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=_GEN_183;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_0 <=_GEN_183;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_0 <=_GEN_761;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_0 <=_GEN_523;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_1[0])
                                 begin 
                                   sectored_entries_0_5_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_1 <=_GEN_184;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=_GEN_184;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=_GEN_184;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_1 <=_GEN_184;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_1 <=_GEN_762;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_1 <=_GEN_524;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_2[0])
                                 begin 
                                   sectored_entries_0_5_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_2 <=_GEN_185;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=_GEN_185;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=_GEN_185;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_2 <=_GEN_185;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_2 <=_GEN_763;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_2 <=_GEN_525;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_3[0])
                                 begin 
                                   sectored_entries_0_5_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_3 <=_GEN_186;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=_GEN_186;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=_GEN_186;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_3 <=_GEN_186;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_3 <=_GEN_764;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_3 <=_GEN_526;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                sectored_entries_0_6_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_6_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_6_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_6_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_6_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_0[0])
                                 begin 
                                   sectored_entries_0_6_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_0 <=_GEN_209;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=_GEN_209;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=_GEN_209;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_0 <=_GEN_209;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_0 <=_GEN_789;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_0 <=_GEN_533;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_1[0])
                                 begin 
                                   sectored_entries_0_6_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_1 <=_GEN_210;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=_GEN_210;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=_GEN_210;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_1 <=_GEN_210;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_1 <=_GEN_790;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_1 <=_GEN_534;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_2[0])
                                 begin 
                                   sectored_entries_0_6_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_2 <=_GEN_211;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=_GEN_211;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=_GEN_211;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_2 <=_GEN_211;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_2 <=_GEN_791;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_2 <=_GEN_535;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_3[0])
                                 begin 
                                   sectored_entries_0_6_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_3 <=_GEN_212;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=_GEN_212;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=_GEN_212;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_3 <=_GEN_212;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_3 <=_GEN_792;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_3 <=_GEN_536;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                sectored_entries_0_7_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_7_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_7_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_7_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_7_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_0[0])
                                 begin 
                                   sectored_entries_0_7_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_0 <=_GEN_235;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=_GEN_235;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=_GEN_235;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_0 <=_GEN_235;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_0 <=_GEN_817;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_0 <=_GEN_543;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_1[0])
                                 begin 
                                   sectored_entries_0_7_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_1 <=_GEN_236;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=_GEN_236;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=_GEN_236;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_1 <=_GEN_236;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_1 <=_GEN_818;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_1 <=_GEN_544;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_2[0])
                                 begin 
                                   sectored_entries_0_7_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_2 <=_GEN_237;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=_GEN_237;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=_GEN_237;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_2 <=_GEN_237;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_2 <=_GEN_819;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_2 <=_GEN_545;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_3[0])
                                 begin 
                                   sectored_entries_0_7_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_3 <=_GEN_238;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=_GEN_238;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=_GEN_238;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_3 <=_GEN_238;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_3 <=_GEN_820;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_3 <=_GEN_546;
                  end 
         if (metaReset)
            begin 
              superpage_entries_0_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_3)
                              begin 
                                superpage_entries_0_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_0_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_3)
                              begin 
                                superpage_entries_0_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_0_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_3)
                              begin 
                                superpage_entries_0_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_0_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_0_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_0)
                            begin 
                              superpage_entries_0_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_3)
                                              begin 
                                                if (invalidate_refill)
                                                   begin 
                                                     superpage_entries_0_valid_0 <=1'h0;
                                                   end 
                                                 else 
                                                   begin 
                                                     superpage_entries_0_valid_0 <=1'h1;
                                                   end 
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_0_valid_0 <=_GEN_827;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_3)
                                    begin 
                                      if (invalidate_refill)
                                         begin 
                                           superpage_entries_0_valid_0 <=1'h0;
                                         end 
                                       else 
                                         begin 
                                           superpage_entries_0_valid_0 <=1'h1;
                                         end 
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              superpage_entries_1_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_4)
                              begin 
                                superpage_entries_1_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_1_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_4)
                              begin 
                                superpage_entries_1_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_1_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_4)
                              begin 
                                superpage_entries_1_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_1_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_1_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_1)
                            begin 
                              superpage_entries_1_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_4)
                                              begin 
                                                if (invalidate_refill)
                                                   begin 
                                                     superpage_entries_1_valid_0 <=1'h0;
                                                   end 
                                                 else 
                                                   begin 
                                                     superpage_entries_1_valid_0 <=1'h1;
                                                   end 
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_1_valid_0 <=_GEN_831;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_4)
                                    begin 
                                      if (invalidate_refill)
                                         begin 
                                           superpage_entries_1_valid_0 <=1'h0;
                                         end 
                                       else 
                                         begin 
                                           superpage_entries_1_valid_0 <=1'h1;
                                         end 
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              superpage_entries_2_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_5)
                              begin 
                                superpage_entries_2_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_2_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_5)
                              begin 
                                superpage_entries_2_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_2_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_5)
                              begin 
                                superpage_entries_2_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_2_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_2_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_2)
                            begin 
                              superpage_entries_2_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_5)
                                              begin 
                                                superpage_entries_2_valid_0 <=_GEN_32;
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_2_valid_0 <=_GEN_835;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_5)
                                    begin 
                                      superpage_entries_2_valid_0 <=_GEN_32;
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              superpage_entries_3_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_6)
                              begin 
                                superpage_entries_3_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_3_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_6)
                              begin 
                                superpage_entries_3_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_3_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_6)
                              begin 
                                superpage_entries_3_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_3_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_3_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_3)
                            begin 
                              superpage_entries_3_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_6)
                                              begin 
                                                superpage_entries_3_valid_0 <=_GEN_32;
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_3_valid_0 <=_GEN_839;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_6)
                                    begin 
                                      superpage_entries_3_valid_0 <=_GEN_32;
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              special_entry_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (~io_ptw_resp_bits_homogeneous)
                    begin 
                      special_entry_level <=io_ptw_resp_bits_level;
                    end 
               end 
         if (metaReset)
            begin 
              special_entry_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (~io_ptw_resp_bits_homogeneous)
                    begin 
                      special_entry_tag <=r_refill_tag;
                    end 
               end 
         if (metaReset)
            begin 
              special_entry_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (~io_ptw_resp_bits_homogeneous)
                    begin 
                      special_entry_data_0 <=_special_entry_data_0_T;
                    end 
               end 
         if (metaReset)
            begin 
              special_entry_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 special_entry_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_hitsVec_T_106)
                            begin 
                              special_entry_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (~io_ptw_resp_bits_homogeneous)
                                    begin 
                                      special_entry_valid_0 <=_GEN_32;
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         special_entry_valid_0 <=_GEN_843;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (~io_ptw_resp_bits_homogeneous)
                          begin 
                            special_entry_valid_0 <=_GEN_32;
                          end 
                     end 
         if (metaReset)
            begin 
              state <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 state <=2'h0;
               end 
             else 
               if (io_ptw_resp_valid)
                  begin 
                    state <=2'h0;
                  end 
                else 
                  if (_T_45)
                     begin 
                       state <=2'h3;
                     end 
                   else 
                     if (_invalidate_refill_T)
                        begin 
                          if (io_ptw_req_ready)
                             begin 
                               if (io_sfence_valid)
                                  begin 
                                    state <=2'h3;
                                  end 
                                else 
                                  begin 
                                    state <=2'h2;
                                  end 
                             end 
                           else 
                             if (io_sfence_valid)
                                begin 
                                  state <=2'h0;
                                end 
                              else 
                                if (_T_42)
                                   begin 
                                     state <=2'h1;
                                   end 
                        end 
                      else 
                        if (_T_42)
                           begin 
                             state <=2'h1;
                           end 
         if (metaReset)
            begin 
              r_refill_tag <=27'h0;
            end 
          else 
            if (_T_42)
               begin 
                 r_refill_tag <=vpn;
               end 
         if (metaReset)
            begin 
              r_superpage_repl_addr <=2'h0;
            end 
          else 
            if (_T_42)
               begin 
                 if (_r_superpage_repl_addr_T_3)
                    begin 
                      r_superpage_repl_addr <=_r_superpage_repl_addr_T_2;
                    end 
                  else 
                    if (_r_superpage_repl_addr_T_5)
                       begin 
                         r_superpage_repl_addr <=2'h0;
                       end 
                     else 
                       if (_r_superpage_repl_addr_T_6)
                          begin 
                            r_superpage_repl_addr <=2'h1;
                          end 
                        else 
                          if (_r_superpage_repl_addr_T_7)
                             begin 
                               r_superpage_repl_addr <=2'h2;
                             end 
                           else 
                             begin 
                               r_superpage_repl_addr <=2'h3;
                             end 
               end 
         if (metaReset)
            begin 
              r_sectored_repl_addr <=3'h0;
            end 
          else 
            if (_T_42)
               begin 
                 if (_r_sectored_repl_addr_T_7)
                    begin 
                      r_sectored_repl_addr <=_r_sectored_repl_addr_T_6;
                    end 
                  else 
                    if (_r_sectored_repl_addr_T_9)
                       begin 
                         r_sectored_repl_addr <=3'h0;
                       end 
                     else 
                       if (_r_sectored_repl_addr_T_10)
                          begin 
                            r_sectored_repl_addr <=3'h1;
                          end 
                        else 
                          if (_r_sectored_repl_addr_T_11)
                             begin 
                               r_sectored_repl_addr <=3'h2;
                             end 
                           else 
                             if (_r_sectored_repl_addr_T_12)
                                begin 
                                  r_sectored_repl_addr <=3'h3;
                                end 
                              else 
                                if (_r_sectored_repl_addr_T_13)
                                   begin 
                                     r_sectored_repl_addr <=3'h4;
                                   end 
                                 else 
                                   if (_r_sectored_repl_addr_T_14)
                                      begin 
                                        r_sectored_repl_addr <=3'h5;
                                      end 
                                    else 
                                      if (_r_sectored_repl_addr_T_15)
                                         begin 
                                           r_sectored_repl_addr <=3'h6;
                                         end 
                                       else 
                                         begin 
                                           r_sectored_repl_addr <=3'h7;
                                         end 
               end 
         if (metaReset)
            begin 
              r_sectored_hit_addr <=3'h0;
            end 
          else 
            if (_T_42)
               begin 
                 r_sectored_hit_addr <=state_vec_0_touch_way_sized;
               end 
         if (metaReset)
            begin 
              r_sectored_hit <=1'h0;
            end 
          else 
            if (_T_42)
               begin 
                 r_sectored_hit <=_T_30;
               end 
         if (metaReset)
            begin 
              state_vec_0 <=7'h0;
            end 
          else 
            if (reset)
               begin 
                 state_vec_0 <=7'h0;
               end 
             else 
               if (_T_23)
                  begin 
                    if (_T_30)
                       begin 
                         state_vec_0 <=_state_vec_0_T_16;
                       end 
                  end 
         if (metaReset)
            begin 
              state_reg_1 <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 state_reg_1 <=3'h0;
               end 
             else 
               if (_T_23)
                  begin 
                    if (_T_37)
                       begin 
                         state_reg_1 <=_state_reg_T_6;
                       end 
                  end 
         if (io_sfence_valid&~_T_51)
            begin $display("Assertion failed\n    at TLB.scala:385 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n");
            end 
         if (io_sfence_valid&~_T_51)
            begin $display("fatal");
            end 
         TLB_state <=TLB_xor0;
         if (!(TLB_cov_read_data))
            begin 
              TLB_covSum <=TLB_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              TLB_metaAssert <=1'h0;
            end 
          else 
            begin 
              TLB_metaAssert <=TLB_metaAssert|TLB_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (TLB_cov_write_en&TLB_cov_write_mask)
            begin 
              TLB_cov [TLB_cov_write_addr]<=TLB_cov_write_data;
            end 
       end
  
endmodule
 
module MaxPeriodFibonacciLFSR (
  input clock,
  input reset,
  input io_increment,
  output io_out_0,
  output io_out_1,
  output io_out_2,
  output io_out_3,
  output io_out_4,
  output io_out_5,
  output io_out_6,
  output io_out_7,
  output io_out_8,
  output io_out_9,
  output io_out_10,
  output io_out_11,
  output io_out_12,
  output io_out_13,
  output io_out_14,
  output io_out_15,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg state_0 ;  
   reg [31:0] _RAND_0 ;  
   reg state_1 ;  
   reg [31:0] _RAND_1 ;  
   reg state_2 ;  
   reg [31:0] _RAND_2 ;  
   reg state_3 ;  
   reg [31:0] _RAND_3 ;  
   reg state_4 ;  
   reg [31:0] _RAND_4 ;  
   reg state_5 ;  
   reg [31:0] _RAND_5 ;  
   reg state_6 ;  
   reg [31:0] _RAND_6 ;  
   reg state_7 ;  
   reg [31:0] _RAND_7 ;  
   reg state_8 ;  
   reg [31:0] _RAND_8 ;  
   reg state_9 ;  
   reg [31:0] _RAND_9 ;  
   reg state_10 ;  
   reg [31:0] _RAND_10 ;  
   reg state_11 ;  
   reg [31:0] _RAND_11 ;  
   reg state_12 ;  
   reg [31:0] _RAND_12 ;  
   reg state_13 ;  
   reg [31:0] _RAND_13 ;  
   reg state_14 ;  
   reg [31:0] _RAND_14 ;  
   reg state_15 ;  
   reg [31:0] _RAND_15 ;  
   wire _T ;  
   wire _T_1 ;  
   wire _T_2 ;  
   wire _GEN_0 ;  
   wire [29:0] MaxPeriodFibonacciLFSR_covSum ;  
  assign _T=state_15^state_13; 
  assign _T_1=_T^state_12; 
  assign _T_2=_T_1^state_10; 
  assign _GEN_0=io_increment ? _T_2:state_0; 
  assign io_out_0=state_0; 
  assign io_out_1=state_1; 
  assign io_out_2=state_2; 
  assign io_out_3=state_3; 
  assign io_out_4=state_4; 
  assign io_out_5=state_5; 
  assign io_out_6=state_6; 
  assign io_out_7=state_7; 
  assign io_out_8=state_8; 
  assign io_out_9=state_9; 
  assign io_out_10=state_10; 
  assign io_out_11=state_11; 
  assign io_out_12=state_12; 
  assign io_out_13=state_13; 
  assign io_out_14=state_14; 
  assign io_out_15=state_15; 
  assign MaxPeriodFibonacciLFSR_covSum=30'h0; 
  assign io_covSum=MaxPeriodFibonacciLFSR_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              state_0 <=1'h0;
            end 
          else 
            begin 
              state_0 <=reset|_GEN_0;
            end 
         if (metaReset)
            begin 
              state_1 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_1 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_1 <=state_0;
                  end 
         if (metaReset)
            begin 
              state_2 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_2 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_2 <=state_1;
                  end 
         if (metaReset)
            begin 
              state_3 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_3 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_3 <=state_2;
                  end 
         if (metaReset)
            begin 
              state_4 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_4 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_4 <=state_3;
                  end 
         if (metaReset)
            begin 
              state_5 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_5 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_5 <=state_4;
                  end 
         if (metaReset)
            begin 
              state_6 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_6 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_6 <=state_5;
                  end 
         if (metaReset)
            begin 
              state_7 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_7 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_7 <=state_6;
                  end 
         if (metaReset)
            begin 
              state_8 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_8 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_8 <=state_7;
                  end 
         if (metaReset)
            begin 
              state_9 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_9 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_9 <=state_8;
                  end 
         if (metaReset)
            begin 
              state_10 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_10 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_10 <=state_9;
                  end 
         if (metaReset)
            begin 
              state_11 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_11 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_11 <=state_10;
                  end 
         if (metaReset)
            begin 
              state_12 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_12 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_12 <=state_11;
                  end 
         if (metaReset)
            begin 
              state_13 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_13 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_13 <=state_12;
                  end 
         if (metaReset)
            begin 
              state_14 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_14 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_14 <=state_13;
                  end 
         if (metaReset)
            begin 
              state_15 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 state_15 <=1'h0;
               end 
             else 
               if (io_increment)
                  begin 
                    state_15 <=state_14;
                  end 
       end
  
endmodule
 
module DCacheModuleImpl_Anon_1 (
  input io_in_0_valid,
  input [39:0] io_in_0_bits_addr,
  input [5:0] io_in_0_bits_idx,
  input io_in_1_valid,
  input [39:0] io_in_1_bits_addr,
  input [5:0] io_in_1_bits_idx,
  input [21:0] io_in_1_bits_data,
  input io_in_2_valid,
  input [39:0] io_in_2_bits_addr,
  input [5:0] io_in_2_bits_idx,
  input [3:0] io_in_2_bits_way_en,
  input [21:0] io_in_2_bits_data,
  input io_in_3_valid,
  input [39:0] io_in_3_bits_addr,
  input [5:0] io_in_3_bits_idx,
  input [3:0] io_in_3_bits_way_en,
  input [21:0] io_in_3_bits_data,
  output io_in_4_ready,
  input io_in_4_valid,
  input [39:0] io_in_4_bits_addr,
  input [5:0] io_in_4_bits_idx,
  input [3:0] io_in_4_bits_way_en,
  input [21:0] io_in_4_bits_data,
  output io_in_5_ready,
  input io_in_5_valid,
  input [39:0] io_in_5_bits_addr,
  input [5:0] io_in_5_bits_idx,
  output io_in_6_ready,
  input io_in_6_valid,
  input [39:0] io_in_6_bits_addr,
  input [5:0] io_in_6_bits_idx,
  input [3:0] io_in_6_bits_way_en,
  input [21:0] io_in_6_bits_data,
  output io_in_7_ready,
  input io_in_7_valid,
  input [39:0] io_in_7_bits_addr,
  input [5:0] io_in_7_bits_idx,
  input [3:0] io_in_7_bits_way_en,
  input [21:0] io_in_7_bits_data,
  output io_out_valid,
  output io_out_bits_write,
  output [39:0] io_out_bits_addr,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [21:0] io_out_bits_data,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [21:0] _GEN_1 ;  
   wire [3:0] _GEN_2 ;  
   wire [5:0] _GEN_3 ;  
   wire [39:0] _GEN_4 ;  
   wire [21:0] _GEN_13 ;  
   wire [3:0] _GEN_14 ;  
   wire [5:0] _GEN_15 ;  
   wire [39:0] _GEN_16 ;  
   wire [21:0] _GEN_19 ;  
   wire [3:0] _GEN_20 ;  
   wire [5:0] _GEN_21 ;  
   wire [39:0] _GEN_22 ;  
   wire _GEN_23 ;  
   wire [21:0] _GEN_25 ;  
   wire [3:0] _GEN_26 ;  
   wire [5:0] _GEN_27 ;  
   wire [39:0] _GEN_28 ;  
   wire _GEN_29 ;  
   wire [21:0] _GEN_31 ;  
   wire [3:0] _GEN_32 ;  
   wire [5:0] _GEN_33 ;  
   wire [39:0] _GEN_34 ;  
   wire _GEN_35 ;  
   wire _grant_T ;  
   wire _grant_T_1 ;  
   wire _grant_T_2 ;  
   wire _grant_T_3 ;  
   wire _grant_T_5 ;  
   wire grant_7 ;  
   wire [29:0] DCacheModuleImpl_Anon_1_covSum ;  
  assign _GEN_1=io_in_6_valid ? io_in_6_bits_data:io_in_7_bits_data; 
  assign _GEN_2=io_in_6_valid ? io_in_6_bits_way_en:io_in_7_bits_way_en; 
  assign _GEN_3=io_in_6_valid ? io_in_6_bits_idx:io_in_7_bits_idx; 
  assign _GEN_4=io_in_6_valid ? io_in_6_bits_addr:io_in_7_bits_addr; 
  assign _GEN_13=io_in_4_valid ? io_in_4_bits_data:_GEN_1; 
  assign _GEN_14=io_in_4_valid ? io_in_4_bits_way_en:_GEN_2; 
  assign _GEN_15=io_in_4_valid ? io_in_4_bits_idx:_GEN_3; 
  assign _GEN_16=io_in_4_valid ? io_in_4_bits_addr:_GEN_4; 
  assign _GEN_19=io_in_3_valid ? io_in_3_bits_data:_GEN_13; 
  assign _GEN_20=io_in_3_valid ? io_in_3_bits_way_en:_GEN_14; 
  assign _GEN_21=io_in_3_valid ? io_in_3_bits_idx:_GEN_15; 
  assign _GEN_22=io_in_3_valid ? io_in_3_bits_addr:_GEN_16; 
  assign _GEN_23=io_in_3_valid|io_in_4_valid; 
  assign _GEN_25=io_in_2_valid ? io_in_2_bits_data:_GEN_19; 
  assign _GEN_26=io_in_2_valid ? io_in_2_bits_way_en:_GEN_20; 
  assign _GEN_27=io_in_2_valid ? io_in_2_bits_idx:_GEN_21; 
  assign _GEN_28=io_in_2_valid ? io_in_2_bits_addr:_GEN_22; 
  assign _GEN_29=io_in_2_valid|_GEN_23; 
  assign _GEN_31=io_in_1_valid ? io_in_1_bits_data:_GEN_25; 
  assign _GEN_32=io_in_1_valid ? 4'h0:_GEN_26; 
  assign _GEN_33=io_in_1_valid ? io_in_1_bits_idx:_GEN_27; 
  assign _GEN_34=io_in_1_valid ? io_in_1_bits_addr:_GEN_28; 
  assign _GEN_35=io_in_1_valid|_GEN_29; 
  assign _grant_T=io_in_0_valid|io_in_1_valid; 
  assign _grant_T_1=_grant_T|io_in_2_valid; 
  assign _grant_T_2=_grant_T_1|io_in_3_valid; 
  assign _grant_T_3=_grant_T_2|io_in_4_valid; 
  assign _grant_T_5=_grant_T_3|io_in_6_valid; 
  assign grant_7=~_grant_T_5; 
  assign io_in_4_ready=~_grant_T_2; 
  assign io_in_5_ready=~_grant_T_3; 
  assign io_in_6_ready=~_grant_T_3; 
  assign io_in_7_ready=~_grant_T_5; 
  assign io_out_valid=~grant_7|io_in_7_valid; 
  assign io_out_bits_write=io_in_0_valid|_GEN_35; 
  assign io_out_bits_addr=io_in_0_valid ? io_in_0_bits_addr:_GEN_34; 
  assign io_out_bits_idx=io_in_0_valid ? io_in_0_bits_idx:_GEN_33; 
  assign io_out_bits_way_en=io_in_0_valid ? 4'hf:_GEN_32; 
  assign io_out_bits_data=io_in_0_valid ? 22'h0:_GEN_31; 
  assign DCacheModuleImpl_Anon_1_covSum=30'h0; 
  assign io_covSum=DCacheModuleImpl_Anon_1_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module DCacheDataArray (
  input clock,
  input io_req_valid,
  input [11:0] io_req_bits_addr,
  input io_req_bits_write,
  input [63:0] io_req_bits_wdata,
  input [7:0] io_req_bits_eccMask,
  input [3:0] io_req_bits_way_en,
  output [63:0] io_resp_0,
  output [63:0] io_resp_1,
  output [63:0] io_resp_2,
  output [63:0] io_resp_3,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg [7:0] data_arrays_0_0[0:511] ;  
   reg [31:0] _RAND_0 ;  
   wire [7:0] data_arrays_0_0_rdata_data_data ;  
   wire [8:0] data_arrays_0_0_rdata_data_addr ;  
   wire [7:0] data_arrays_0_0_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_0_rdata_MPORT_addr ;  
   wire data_arrays_0_0_rdata_MPORT_mask ;  
   wire data_arrays_0_0_rdata_MPORT_en ;  
   reg data_arrays_0_0_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_1 ;  
   reg [8:0] data_arrays_0_0_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_2 ;  
   reg [7:0] data_arrays_0_1[0:511] ;  
   reg [31:0] _RAND_3 ;  
   wire [7:0] data_arrays_0_1_rdata_data_data ;  
   wire [8:0] data_arrays_0_1_rdata_data_addr ;  
   wire [7:0] data_arrays_0_1_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_1_rdata_MPORT_addr ;  
   wire data_arrays_0_1_rdata_MPORT_mask ;  
   wire data_arrays_0_1_rdata_MPORT_en ;  
   reg data_arrays_0_1_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_4 ;  
   reg [8:0] data_arrays_0_1_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_5 ;  
   reg [7:0] data_arrays_0_2[0:511] ;  
   reg [31:0] _RAND_6 ;  
   wire [7:0] data_arrays_0_2_rdata_data_data ;  
   wire [8:0] data_arrays_0_2_rdata_data_addr ;  
   wire [7:0] data_arrays_0_2_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_2_rdata_MPORT_addr ;  
   wire data_arrays_0_2_rdata_MPORT_mask ;  
   wire data_arrays_0_2_rdata_MPORT_en ;  
   reg data_arrays_0_2_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_7 ;  
   reg [8:0] data_arrays_0_2_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_8 ;  
   reg [7:0] data_arrays_0_3[0:511] ;  
   reg [31:0] _RAND_9 ;  
   wire [7:0] data_arrays_0_3_rdata_data_data ;  
   wire [8:0] data_arrays_0_3_rdata_data_addr ;  
   wire [7:0] data_arrays_0_3_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_3_rdata_MPORT_addr ;  
   wire data_arrays_0_3_rdata_MPORT_mask ;  
   wire data_arrays_0_3_rdata_MPORT_en ;  
   reg data_arrays_0_3_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_10 ;  
   reg [8:0] data_arrays_0_3_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_11 ;  
   reg [7:0] data_arrays_0_4[0:511] ;  
   reg [31:0] _RAND_12 ;  
   wire [7:0] data_arrays_0_4_rdata_data_data ;  
   wire [8:0] data_arrays_0_4_rdata_data_addr ;  
   wire [7:0] data_arrays_0_4_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_4_rdata_MPORT_addr ;  
   wire data_arrays_0_4_rdata_MPORT_mask ;  
   wire data_arrays_0_4_rdata_MPORT_en ;  
   reg data_arrays_0_4_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_13 ;  
   reg [8:0] data_arrays_0_4_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_14 ;  
   reg [7:0] data_arrays_0_5[0:511] ;  
   reg [31:0] _RAND_15 ;  
   wire [7:0] data_arrays_0_5_rdata_data_data ;  
   wire [8:0] data_arrays_0_5_rdata_data_addr ;  
   wire [7:0] data_arrays_0_5_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_5_rdata_MPORT_addr ;  
   wire data_arrays_0_5_rdata_MPORT_mask ;  
   wire data_arrays_0_5_rdata_MPORT_en ;  
   reg data_arrays_0_5_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_16 ;  
   reg [8:0] data_arrays_0_5_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_17 ;  
   reg [7:0] data_arrays_0_6[0:511] ;  
   reg [31:0] _RAND_18 ;  
   wire [7:0] data_arrays_0_6_rdata_data_data ;  
   wire [8:0] data_arrays_0_6_rdata_data_addr ;  
   wire [7:0] data_arrays_0_6_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_6_rdata_MPORT_addr ;  
   wire data_arrays_0_6_rdata_MPORT_mask ;  
   wire data_arrays_0_6_rdata_MPORT_en ;  
   reg data_arrays_0_6_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_19 ;  
   reg [8:0] data_arrays_0_6_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_20 ;  
   reg [7:0] data_arrays_0_7[0:511] ;  
   reg [31:0] _RAND_21 ;  
   wire [7:0] data_arrays_0_7_rdata_data_data ;  
   wire [8:0] data_arrays_0_7_rdata_data_addr ;  
   wire [7:0] data_arrays_0_7_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_7_rdata_MPORT_addr ;  
   wire data_arrays_0_7_rdata_MPORT_mask ;  
   wire data_arrays_0_7_rdata_MPORT_en ;  
   reg data_arrays_0_7_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_22 ;  
   reg [8:0] data_arrays_0_7_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_23 ;  
   reg [7:0] data_arrays_0_8[0:511] ;  
   reg [31:0] _RAND_24 ;  
   wire [7:0] data_arrays_0_8_rdata_data_data ;  
   wire [8:0] data_arrays_0_8_rdata_data_addr ;  
   wire [7:0] data_arrays_0_8_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_8_rdata_MPORT_addr ;  
   wire data_arrays_0_8_rdata_MPORT_mask ;  
   wire data_arrays_0_8_rdata_MPORT_en ;  
   reg data_arrays_0_8_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_25 ;  
   reg [8:0] data_arrays_0_8_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_26 ;  
   reg [7:0] data_arrays_0_9[0:511] ;  
   reg [31:0] _RAND_27 ;  
   wire [7:0] data_arrays_0_9_rdata_data_data ;  
   wire [8:0] data_arrays_0_9_rdata_data_addr ;  
   wire [7:0] data_arrays_0_9_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_9_rdata_MPORT_addr ;  
   wire data_arrays_0_9_rdata_MPORT_mask ;  
   wire data_arrays_0_9_rdata_MPORT_en ;  
   reg data_arrays_0_9_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_28 ;  
   reg [8:0] data_arrays_0_9_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_29 ;  
   reg [7:0] data_arrays_0_10[0:511] ;  
   reg [31:0] _RAND_30 ;  
   wire [7:0] data_arrays_0_10_rdata_data_data ;  
   wire [8:0] data_arrays_0_10_rdata_data_addr ;  
   wire [7:0] data_arrays_0_10_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_10_rdata_MPORT_addr ;  
   wire data_arrays_0_10_rdata_MPORT_mask ;  
   wire data_arrays_0_10_rdata_MPORT_en ;  
   reg data_arrays_0_10_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_31 ;  
   reg [8:0] data_arrays_0_10_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_32 ;  
   reg [7:0] data_arrays_0_11[0:511] ;  
   reg [31:0] _RAND_33 ;  
   wire [7:0] data_arrays_0_11_rdata_data_data ;  
   wire [8:0] data_arrays_0_11_rdata_data_addr ;  
   wire [7:0] data_arrays_0_11_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_11_rdata_MPORT_addr ;  
   wire data_arrays_0_11_rdata_MPORT_mask ;  
   wire data_arrays_0_11_rdata_MPORT_en ;  
   reg data_arrays_0_11_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_34 ;  
   reg [8:0] data_arrays_0_11_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_35 ;  
   reg [7:0] data_arrays_0_12[0:511] ;  
   reg [31:0] _RAND_36 ;  
   wire [7:0] data_arrays_0_12_rdata_data_data ;  
   wire [8:0] data_arrays_0_12_rdata_data_addr ;  
   wire [7:0] data_arrays_0_12_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_12_rdata_MPORT_addr ;  
   wire data_arrays_0_12_rdata_MPORT_mask ;  
   wire data_arrays_0_12_rdata_MPORT_en ;  
   reg data_arrays_0_12_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_37 ;  
   reg [8:0] data_arrays_0_12_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_38 ;  
   reg [7:0] data_arrays_0_13[0:511] ;  
   reg [31:0] _RAND_39 ;  
   wire [7:0] data_arrays_0_13_rdata_data_data ;  
   wire [8:0] data_arrays_0_13_rdata_data_addr ;  
   wire [7:0] data_arrays_0_13_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_13_rdata_MPORT_addr ;  
   wire data_arrays_0_13_rdata_MPORT_mask ;  
   wire data_arrays_0_13_rdata_MPORT_en ;  
   reg data_arrays_0_13_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_40 ;  
   reg [8:0] data_arrays_0_13_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_41 ;  
   reg [7:0] data_arrays_0_14[0:511] ;  
   reg [31:0] _RAND_42 ;  
   wire [7:0] data_arrays_0_14_rdata_data_data ;  
   wire [8:0] data_arrays_0_14_rdata_data_addr ;  
   wire [7:0] data_arrays_0_14_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_14_rdata_MPORT_addr ;  
   wire data_arrays_0_14_rdata_MPORT_mask ;  
   wire data_arrays_0_14_rdata_MPORT_en ;  
   reg data_arrays_0_14_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_43 ;  
   reg [8:0] data_arrays_0_14_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_44 ;  
   reg [7:0] data_arrays_0_15[0:511] ;  
   reg [31:0] _RAND_45 ;  
   wire [7:0] data_arrays_0_15_rdata_data_data ;  
   wire [8:0] data_arrays_0_15_rdata_data_addr ;  
   wire [7:0] data_arrays_0_15_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_15_rdata_MPORT_addr ;  
   wire data_arrays_0_15_rdata_MPORT_mask ;  
   wire data_arrays_0_15_rdata_MPORT_en ;  
   reg data_arrays_0_15_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_46 ;  
   reg [8:0] data_arrays_0_15_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_47 ;  
   reg [7:0] data_arrays_0_16[0:511] ;  
   reg [31:0] _RAND_48 ;  
   wire [7:0] data_arrays_0_16_rdata_data_data ;  
   wire [8:0] data_arrays_0_16_rdata_data_addr ;  
   wire [7:0] data_arrays_0_16_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_16_rdata_MPORT_addr ;  
   wire data_arrays_0_16_rdata_MPORT_mask ;  
   wire data_arrays_0_16_rdata_MPORT_en ;  
   reg data_arrays_0_16_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_49 ;  
   reg [8:0] data_arrays_0_16_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_50 ;  
   reg [7:0] data_arrays_0_17[0:511] ;  
   reg [31:0] _RAND_51 ;  
   wire [7:0] data_arrays_0_17_rdata_data_data ;  
   wire [8:0] data_arrays_0_17_rdata_data_addr ;  
   wire [7:0] data_arrays_0_17_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_17_rdata_MPORT_addr ;  
   wire data_arrays_0_17_rdata_MPORT_mask ;  
   wire data_arrays_0_17_rdata_MPORT_en ;  
   reg data_arrays_0_17_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_52 ;  
   reg [8:0] data_arrays_0_17_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_53 ;  
   reg [7:0] data_arrays_0_18[0:511] ;  
   reg [31:0] _RAND_54 ;  
   wire [7:0] data_arrays_0_18_rdata_data_data ;  
   wire [8:0] data_arrays_0_18_rdata_data_addr ;  
   wire [7:0] data_arrays_0_18_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_18_rdata_MPORT_addr ;  
   wire data_arrays_0_18_rdata_MPORT_mask ;  
   wire data_arrays_0_18_rdata_MPORT_en ;  
   reg data_arrays_0_18_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_55 ;  
   reg [8:0] data_arrays_0_18_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_56 ;  
   reg [7:0] data_arrays_0_19[0:511] ;  
   reg [31:0] _RAND_57 ;  
   wire [7:0] data_arrays_0_19_rdata_data_data ;  
   wire [8:0] data_arrays_0_19_rdata_data_addr ;  
   wire [7:0] data_arrays_0_19_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_19_rdata_MPORT_addr ;  
   wire data_arrays_0_19_rdata_MPORT_mask ;  
   wire data_arrays_0_19_rdata_MPORT_en ;  
   reg data_arrays_0_19_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_58 ;  
   reg [8:0] data_arrays_0_19_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_59 ;  
   reg [7:0] data_arrays_0_20[0:511] ;  
   reg [31:0] _RAND_60 ;  
   wire [7:0] data_arrays_0_20_rdata_data_data ;  
   wire [8:0] data_arrays_0_20_rdata_data_addr ;  
   wire [7:0] data_arrays_0_20_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_20_rdata_MPORT_addr ;  
   wire data_arrays_0_20_rdata_MPORT_mask ;  
   wire data_arrays_0_20_rdata_MPORT_en ;  
   reg data_arrays_0_20_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_61 ;  
   reg [8:0] data_arrays_0_20_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_62 ;  
   reg [7:0] data_arrays_0_21[0:511] ;  
   reg [31:0] _RAND_63 ;  
   wire [7:0] data_arrays_0_21_rdata_data_data ;  
   wire [8:0] data_arrays_0_21_rdata_data_addr ;  
   wire [7:0] data_arrays_0_21_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_21_rdata_MPORT_addr ;  
   wire data_arrays_0_21_rdata_MPORT_mask ;  
   wire data_arrays_0_21_rdata_MPORT_en ;  
   reg data_arrays_0_21_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_64 ;  
   reg [8:0] data_arrays_0_21_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_65 ;  
   reg [7:0] data_arrays_0_22[0:511] ;  
   reg [31:0] _RAND_66 ;  
   wire [7:0] data_arrays_0_22_rdata_data_data ;  
   wire [8:0] data_arrays_0_22_rdata_data_addr ;  
   wire [7:0] data_arrays_0_22_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_22_rdata_MPORT_addr ;  
   wire data_arrays_0_22_rdata_MPORT_mask ;  
   wire data_arrays_0_22_rdata_MPORT_en ;  
   reg data_arrays_0_22_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_67 ;  
   reg [8:0] data_arrays_0_22_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_68 ;  
   reg [7:0] data_arrays_0_23[0:511] ;  
   reg [31:0] _RAND_69 ;  
   wire [7:0] data_arrays_0_23_rdata_data_data ;  
   wire [8:0] data_arrays_0_23_rdata_data_addr ;  
   wire [7:0] data_arrays_0_23_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_23_rdata_MPORT_addr ;  
   wire data_arrays_0_23_rdata_MPORT_mask ;  
   wire data_arrays_0_23_rdata_MPORT_en ;  
   reg data_arrays_0_23_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_70 ;  
   reg [8:0] data_arrays_0_23_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_71 ;  
   reg [7:0] data_arrays_0_24[0:511] ;  
   reg [31:0] _RAND_72 ;  
   wire [7:0] data_arrays_0_24_rdata_data_data ;  
   wire [8:0] data_arrays_0_24_rdata_data_addr ;  
   wire [7:0] data_arrays_0_24_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_24_rdata_MPORT_addr ;  
   wire data_arrays_0_24_rdata_MPORT_mask ;  
   wire data_arrays_0_24_rdata_MPORT_en ;  
   reg data_arrays_0_24_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_73 ;  
   reg [8:0] data_arrays_0_24_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_74 ;  
   reg [7:0] data_arrays_0_25[0:511] ;  
   reg [31:0] _RAND_75 ;  
   wire [7:0] data_arrays_0_25_rdata_data_data ;  
   wire [8:0] data_arrays_0_25_rdata_data_addr ;  
   wire [7:0] data_arrays_0_25_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_25_rdata_MPORT_addr ;  
   wire data_arrays_0_25_rdata_MPORT_mask ;  
   wire data_arrays_0_25_rdata_MPORT_en ;  
   reg data_arrays_0_25_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_76 ;  
   reg [8:0] data_arrays_0_25_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_77 ;  
   reg [7:0] data_arrays_0_26[0:511] ;  
   reg [31:0] _RAND_78 ;  
   wire [7:0] data_arrays_0_26_rdata_data_data ;  
   wire [8:0] data_arrays_0_26_rdata_data_addr ;  
   wire [7:0] data_arrays_0_26_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_26_rdata_MPORT_addr ;  
   wire data_arrays_0_26_rdata_MPORT_mask ;  
   wire data_arrays_0_26_rdata_MPORT_en ;  
   reg data_arrays_0_26_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_79 ;  
   reg [8:0] data_arrays_0_26_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_80 ;  
   reg [7:0] data_arrays_0_27[0:511] ;  
   reg [31:0] _RAND_81 ;  
   wire [7:0] data_arrays_0_27_rdata_data_data ;  
   wire [8:0] data_arrays_0_27_rdata_data_addr ;  
   wire [7:0] data_arrays_0_27_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_27_rdata_MPORT_addr ;  
   wire data_arrays_0_27_rdata_MPORT_mask ;  
   wire data_arrays_0_27_rdata_MPORT_en ;  
   reg data_arrays_0_27_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_82 ;  
   reg [8:0] data_arrays_0_27_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_83 ;  
   reg [7:0] data_arrays_0_28[0:511] ;  
   reg [31:0] _RAND_84 ;  
   wire [7:0] data_arrays_0_28_rdata_data_data ;  
   wire [8:0] data_arrays_0_28_rdata_data_addr ;  
   wire [7:0] data_arrays_0_28_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_28_rdata_MPORT_addr ;  
   wire data_arrays_0_28_rdata_MPORT_mask ;  
   wire data_arrays_0_28_rdata_MPORT_en ;  
   reg data_arrays_0_28_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_85 ;  
   reg [8:0] data_arrays_0_28_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_86 ;  
   reg [7:0] data_arrays_0_29[0:511] ;  
   reg [31:0] _RAND_87 ;  
   wire [7:0] data_arrays_0_29_rdata_data_data ;  
   wire [8:0] data_arrays_0_29_rdata_data_addr ;  
   wire [7:0] data_arrays_0_29_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_29_rdata_MPORT_addr ;  
   wire data_arrays_0_29_rdata_MPORT_mask ;  
   wire data_arrays_0_29_rdata_MPORT_en ;  
   reg data_arrays_0_29_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_88 ;  
   reg [8:0] data_arrays_0_29_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_89 ;  
   reg [7:0] data_arrays_0_30[0:511] ;  
   reg [31:0] _RAND_90 ;  
   wire [7:0] data_arrays_0_30_rdata_data_data ;  
   wire [8:0] data_arrays_0_30_rdata_data_addr ;  
   wire [7:0] data_arrays_0_30_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_30_rdata_MPORT_addr ;  
   wire data_arrays_0_30_rdata_MPORT_mask ;  
   wire data_arrays_0_30_rdata_MPORT_en ;  
   reg data_arrays_0_30_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_91 ;  
   reg [8:0] data_arrays_0_30_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_92 ;  
   reg [7:0] data_arrays_0_31[0:511] ;  
   reg [31:0] _RAND_93 ;  
   wire [7:0] data_arrays_0_31_rdata_data_data ;  
   wire [8:0] data_arrays_0_31_rdata_data_addr ;  
   wire [7:0] data_arrays_0_31_rdata_MPORT_data ;  
   wire [8:0] data_arrays_0_31_rdata_MPORT_addr ;  
   wire data_arrays_0_31_rdata_MPORT_mask ;  
   wire data_arrays_0_31_rdata_MPORT_en ;  
   reg data_arrays_0_31_rdata_data_en_pipe_0 ;  
   reg [31:0] _RAND_94 ;  
   reg [8:0] data_arrays_0_31_rdata_data_addr_pipe_0 ;  
   reg [31:0] _RAND_95 ;  
   wire eccMask_0 ;  
   wire eccMask_1 ;  
   wire eccMask_2 ;  
   wire eccMask_3 ;  
   wire eccMask_4 ;  
   wire eccMask_5 ;  
   wire eccMask_6 ;  
   wire eccMask_7 ;  
   wire [31:0] rdata_lo ;  
   wire [31:0] rdata_hi ;  
   wire [31:0] lo ;  
   wire [31:0] hi ;  
   wire [31:0] lo_1 ;  
   wire [31:0] hi_1 ;  
   wire [31:0] lo_2 ;  
   wire [31:0] hi_2 ;  
   wire [29:0] DCacheDataArray_covSum ;  
  assign data_arrays_0_0_rdata_data_addr=data_arrays_0_0_rdata_data_addr_pipe_0; 
  assign data_arrays_0_0_rdata_data_data=data_arrays_0_0[data_arrays_0_0_rdata_data_addr]; 
  assign data_arrays_0_0_rdata_MPORT_data=io_req_bits_wdata[7:0]; 
  assign data_arrays_0_0_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_0_rdata_MPORT_mask=eccMask_0&io_req_bits_way_en[0]; 
  assign data_arrays_0_0_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_1_rdata_data_addr=data_arrays_0_1_rdata_data_addr_pipe_0; 
  assign data_arrays_0_1_rdata_data_data=data_arrays_0_1[data_arrays_0_1_rdata_data_addr]; 
  assign data_arrays_0_1_rdata_MPORT_data=io_req_bits_wdata[15:8]; 
  assign data_arrays_0_1_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_1_rdata_MPORT_mask=eccMask_1&io_req_bits_way_en[0]; 
  assign data_arrays_0_1_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_2_rdata_data_addr=data_arrays_0_2_rdata_data_addr_pipe_0; 
  assign data_arrays_0_2_rdata_data_data=data_arrays_0_2[data_arrays_0_2_rdata_data_addr]; 
  assign data_arrays_0_2_rdata_MPORT_data=io_req_bits_wdata[23:16]; 
  assign data_arrays_0_2_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_2_rdata_MPORT_mask=eccMask_2&io_req_bits_way_en[0]; 
  assign data_arrays_0_2_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_3_rdata_data_addr=data_arrays_0_3_rdata_data_addr_pipe_0; 
  assign data_arrays_0_3_rdata_data_data=data_arrays_0_3[data_arrays_0_3_rdata_data_addr]; 
  assign data_arrays_0_3_rdata_MPORT_data=io_req_bits_wdata[31:24]; 
  assign data_arrays_0_3_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_3_rdata_MPORT_mask=eccMask_3&io_req_bits_way_en[0]; 
  assign data_arrays_0_3_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_4_rdata_data_addr=data_arrays_0_4_rdata_data_addr_pipe_0; 
  assign data_arrays_0_4_rdata_data_data=data_arrays_0_4[data_arrays_0_4_rdata_data_addr]; 
  assign data_arrays_0_4_rdata_MPORT_data=io_req_bits_wdata[39:32]; 
  assign data_arrays_0_4_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_4_rdata_MPORT_mask=eccMask_4&io_req_bits_way_en[0]; 
  assign data_arrays_0_4_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_5_rdata_data_addr=data_arrays_0_5_rdata_data_addr_pipe_0; 
  assign data_arrays_0_5_rdata_data_data=data_arrays_0_5[data_arrays_0_5_rdata_data_addr]; 
  assign data_arrays_0_5_rdata_MPORT_data=io_req_bits_wdata[47:40]; 
  assign data_arrays_0_5_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_5_rdata_MPORT_mask=eccMask_5&io_req_bits_way_en[0]; 
  assign data_arrays_0_5_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_6_rdata_data_addr=data_arrays_0_6_rdata_data_addr_pipe_0; 
  assign data_arrays_0_6_rdata_data_data=data_arrays_0_6[data_arrays_0_6_rdata_data_addr]; 
  assign data_arrays_0_6_rdata_MPORT_data=io_req_bits_wdata[55:48]; 
  assign data_arrays_0_6_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_6_rdata_MPORT_mask=eccMask_6&io_req_bits_way_en[0]; 
  assign data_arrays_0_6_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_7_rdata_data_addr=data_arrays_0_7_rdata_data_addr_pipe_0; 
  assign data_arrays_0_7_rdata_data_data=data_arrays_0_7[data_arrays_0_7_rdata_data_addr]; 
  assign data_arrays_0_7_rdata_MPORT_data=io_req_bits_wdata[63:56]; 
  assign data_arrays_0_7_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_7_rdata_MPORT_mask=eccMask_7&io_req_bits_way_en[0]; 
  assign data_arrays_0_7_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_8_rdata_data_addr=data_arrays_0_8_rdata_data_addr_pipe_0; 
  assign data_arrays_0_8_rdata_data_data=data_arrays_0_8[data_arrays_0_8_rdata_data_addr]; 
  assign data_arrays_0_8_rdata_MPORT_data=io_req_bits_wdata[7:0]; 
  assign data_arrays_0_8_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_8_rdata_MPORT_mask=eccMask_0&io_req_bits_way_en[1]; 
  assign data_arrays_0_8_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_9_rdata_data_addr=data_arrays_0_9_rdata_data_addr_pipe_0; 
  assign data_arrays_0_9_rdata_data_data=data_arrays_0_9[data_arrays_0_9_rdata_data_addr]; 
  assign data_arrays_0_9_rdata_MPORT_data=io_req_bits_wdata[15:8]; 
  assign data_arrays_0_9_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_9_rdata_MPORT_mask=eccMask_1&io_req_bits_way_en[1]; 
  assign data_arrays_0_9_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_10_rdata_data_addr=data_arrays_0_10_rdata_data_addr_pipe_0; 
  assign data_arrays_0_10_rdata_data_data=data_arrays_0_10[data_arrays_0_10_rdata_data_addr]; 
  assign data_arrays_0_10_rdata_MPORT_data=io_req_bits_wdata[23:16]; 
  assign data_arrays_0_10_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_10_rdata_MPORT_mask=eccMask_2&io_req_bits_way_en[1]; 
  assign data_arrays_0_10_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_11_rdata_data_addr=data_arrays_0_11_rdata_data_addr_pipe_0; 
  assign data_arrays_0_11_rdata_data_data=data_arrays_0_11[data_arrays_0_11_rdata_data_addr]; 
  assign data_arrays_0_11_rdata_MPORT_data=io_req_bits_wdata[31:24]; 
  assign data_arrays_0_11_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_11_rdata_MPORT_mask=eccMask_3&io_req_bits_way_en[1]; 
  assign data_arrays_0_11_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_12_rdata_data_addr=data_arrays_0_12_rdata_data_addr_pipe_0; 
  assign data_arrays_0_12_rdata_data_data=data_arrays_0_12[data_arrays_0_12_rdata_data_addr]; 
  assign data_arrays_0_12_rdata_MPORT_data=io_req_bits_wdata[39:32]; 
  assign data_arrays_0_12_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_12_rdata_MPORT_mask=eccMask_4&io_req_bits_way_en[1]; 
  assign data_arrays_0_12_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_13_rdata_data_addr=data_arrays_0_13_rdata_data_addr_pipe_0; 
  assign data_arrays_0_13_rdata_data_data=data_arrays_0_13[data_arrays_0_13_rdata_data_addr]; 
  assign data_arrays_0_13_rdata_MPORT_data=io_req_bits_wdata[47:40]; 
  assign data_arrays_0_13_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_13_rdata_MPORT_mask=eccMask_5&io_req_bits_way_en[1]; 
  assign data_arrays_0_13_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_14_rdata_data_addr=data_arrays_0_14_rdata_data_addr_pipe_0; 
  assign data_arrays_0_14_rdata_data_data=data_arrays_0_14[data_arrays_0_14_rdata_data_addr]; 
  assign data_arrays_0_14_rdata_MPORT_data=io_req_bits_wdata[55:48]; 
  assign data_arrays_0_14_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_14_rdata_MPORT_mask=eccMask_6&io_req_bits_way_en[1]; 
  assign data_arrays_0_14_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_15_rdata_data_addr=data_arrays_0_15_rdata_data_addr_pipe_0; 
  assign data_arrays_0_15_rdata_data_data=data_arrays_0_15[data_arrays_0_15_rdata_data_addr]; 
  assign data_arrays_0_15_rdata_MPORT_data=io_req_bits_wdata[63:56]; 
  assign data_arrays_0_15_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_15_rdata_MPORT_mask=eccMask_7&io_req_bits_way_en[1]; 
  assign data_arrays_0_15_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_16_rdata_data_addr=data_arrays_0_16_rdata_data_addr_pipe_0; 
  assign data_arrays_0_16_rdata_data_data=data_arrays_0_16[data_arrays_0_16_rdata_data_addr]; 
  assign data_arrays_0_16_rdata_MPORT_data=io_req_bits_wdata[7:0]; 
  assign data_arrays_0_16_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_16_rdata_MPORT_mask=eccMask_0&io_req_bits_way_en[2]; 
  assign data_arrays_0_16_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_17_rdata_data_addr=data_arrays_0_17_rdata_data_addr_pipe_0; 
  assign data_arrays_0_17_rdata_data_data=data_arrays_0_17[data_arrays_0_17_rdata_data_addr]; 
  assign data_arrays_0_17_rdata_MPORT_data=io_req_bits_wdata[15:8]; 
  assign data_arrays_0_17_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_17_rdata_MPORT_mask=eccMask_1&io_req_bits_way_en[2]; 
  assign data_arrays_0_17_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_18_rdata_data_addr=data_arrays_0_18_rdata_data_addr_pipe_0; 
  assign data_arrays_0_18_rdata_data_data=data_arrays_0_18[data_arrays_0_18_rdata_data_addr]; 
  assign data_arrays_0_18_rdata_MPORT_data=io_req_bits_wdata[23:16]; 
  assign data_arrays_0_18_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_18_rdata_MPORT_mask=eccMask_2&io_req_bits_way_en[2]; 
  assign data_arrays_0_18_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_19_rdata_data_addr=data_arrays_0_19_rdata_data_addr_pipe_0; 
  assign data_arrays_0_19_rdata_data_data=data_arrays_0_19[data_arrays_0_19_rdata_data_addr]; 
  assign data_arrays_0_19_rdata_MPORT_data=io_req_bits_wdata[31:24]; 
  assign data_arrays_0_19_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_19_rdata_MPORT_mask=eccMask_3&io_req_bits_way_en[2]; 
  assign data_arrays_0_19_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_20_rdata_data_addr=data_arrays_0_20_rdata_data_addr_pipe_0; 
  assign data_arrays_0_20_rdata_data_data=data_arrays_0_20[data_arrays_0_20_rdata_data_addr]; 
  assign data_arrays_0_20_rdata_MPORT_data=io_req_bits_wdata[39:32]; 
  assign data_arrays_0_20_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_20_rdata_MPORT_mask=eccMask_4&io_req_bits_way_en[2]; 
  assign data_arrays_0_20_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_21_rdata_data_addr=data_arrays_0_21_rdata_data_addr_pipe_0; 
  assign data_arrays_0_21_rdata_data_data=data_arrays_0_21[data_arrays_0_21_rdata_data_addr]; 
  assign data_arrays_0_21_rdata_MPORT_data=io_req_bits_wdata[47:40]; 
  assign data_arrays_0_21_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_21_rdata_MPORT_mask=eccMask_5&io_req_bits_way_en[2]; 
  assign data_arrays_0_21_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_22_rdata_data_addr=data_arrays_0_22_rdata_data_addr_pipe_0; 
  assign data_arrays_0_22_rdata_data_data=data_arrays_0_22[data_arrays_0_22_rdata_data_addr]; 
  assign data_arrays_0_22_rdata_MPORT_data=io_req_bits_wdata[55:48]; 
  assign data_arrays_0_22_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_22_rdata_MPORT_mask=eccMask_6&io_req_bits_way_en[2]; 
  assign data_arrays_0_22_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_23_rdata_data_addr=data_arrays_0_23_rdata_data_addr_pipe_0; 
  assign data_arrays_0_23_rdata_data_data=data_arrays_0_23[data_arrays_0_23_rdata_data_addr]; 
  assign data_arrays_0_23_rdata_MPORT_data=io_req_bits_wdata[63:56]; 
  assign data_arrays_0_23_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_23_rdata_MPORT_mask=eccMask_7&io_req_bits_way_en[2]; 
  assign data_arrays_0_23_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_24_rdata_data_addr=data_arrays_0_24_rdata_data_addr_pipe_0; 
  assign data_arrays_0_24_rdata_data_data=data_arrays_0_24[data_arrays_0_24_rdata_data_addr]; 
  assign data_arrays_0_24_rdata_MPORT_data=io_req_bits_wdata[7:0]; 
  assign data_arrays_0_24_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_24_rdata_MPORT_mask=eccMask_0&io_req_bits_way_en[3]; 
  assign data_arrays_0_24_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_25_rdata_data_addr=data_arrays_0_25_rdata_data_addr_pipe_0; 
  assign data_arrays_0_25_rdata_data_data=data_arrays_0_25[data_arrays_0_25_rdata_data_addr]; 
  assign data_arrays_0_25_rdata_MPORT_data=io_req_bits_wdata[15:8]; 
  assign data_arrays_0_25_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_25_rdata_MPORT_mask=eccMask_1&io_req_bits_way_en[3]; 
  assign data_arrays_0_25_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_26_rdata_data_addr=data_arrays_0_26_rdata_data_addr_pipe_0; 
  assign data_arrays_0_26_rdata_data_data=data_arrays_0_26[data_arrays_0_26_rdata_data_addr]; 
  assign data_arrays_0_26_rdata_MPORT_data=io_req_bits_wdata[23:16]; 
  assign data_arrays_0_26_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_26_rdata_MPORT_mask=eccMask_2&io_req_bits_way_en[3]; 
  assign data_arrays_0_26_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_27_rdata_data_addr=data_arrays_0_27_rdata_data_addr_pipe_0; 
  assign data_arrays_0_27_rdata_data_data=data_arrays_0_27[data_arrays_0_27_rdata_data_addr]; 
  assign data_arrays_0_27_rdata_MPORT_data=io_req_bits_wdata[31:24]; 
  assign data_arrays_0_27_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_27_rdata_MPORT_mask=eccMask_3&io_req_bits_way_en[3]; 
  assign data_arrays_0_27_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_28_rdata_data_addr=data_arrays_0_28_rdata_data_addr_pipe_0; 
  assign data_arrays_0_28_rdata_data_data=data_arrays_0_28[data_arrays_0_28_rdata_data_addr]; 
  assign data_arrays_0_28_rdata_MPORT_data=io_req_bits_wdata[39:32]; 
  assign data_arrays_0_28_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_28_rdata_MPORT_mask=eccMask_4&io_req_bits_way_en[3]; 
  assign data_arrays_0_28_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_29_rdata_data_addr=data_arrays_0_29_rdata_data_addr_pipe_0; 
  assign data_arrays_0_29_rdata_data_data=data_arrays_0_29[data_arrays_0_29_rdata_data_addr]; 
  assign data_arrays_0_29_rdata_MPORT_data=io_req_bits_wdata[47:40]; 
  assign data_arrays_0_29_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_29_rdata_MPORT_mask=eccMask_5&io_req_bits_way_en[3]; 
  assign data_arrays_0_29_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_30_rdata_data_addr=data_arrays_0_30_rdata_data_addr_pipe_0; 
  assign data_arrays_0_30_rdata_data_data=data_arrays_0_30[data_arrays_0_30_rdata_data_addr]; 
  assign data_arrays_0_30_rdata_MPORT_data=io_req_bits_wdata[55:48]; 
  assign data_arrays_0_30_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_30_rdata_MPORT_mask=eccMask_6&io_req_bits_way_en[3]; 
  assign data_arrays_0_30_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_31_rdata_data_addr=data_arrays_0_31_rdata_data_addr_pipe_0; 
  assign data_arrays_0_31_rdata_data_data=data_arrays_0_31[data_arrays_0_31_rdata_data_addr]; 
  assign data_arrays_0_31_rdata_MPORT_data=io_req_bits_wdata[63:56]; 
  assign data_arrays_0_31_rdata_MPORT_addr=io_req_bits_addr[11:3]; 
  assign data_arrays_0_31_rdata_MPORT_mask=eccMask_7&io_req_bits_way_en[3]; 
  assign data_arrays_0_31_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign eccMask_0=io_req_bits_eccMask[0]; 
  assign eccMask_1=io_req_bits_eccMask[1]; 
  assign eccMask_2=io_req_bits_eccMask[2]; 
  assign eccMask_3=io_req_bits_eccMask[3]; 
  assign eccMask_4=io_req_bits_eccMask[4]; 
  assign eccMask_5=io_req_bits_eccMask[5]; 
  assign eccMask_6=io_req_bits_eccMask[6]; 
  assign eccMask_7=io_req_bits_eccMask[7]; 
  assign rdata_lo={data_arrays_0_3_rdata_data_data,data_arrays_0_2_rdata_data_data,data_arrays_0_1_rdata_data_data,data_arrays_0_0_rdata_data_data}; 
  assign rdata_hi={data_arrays_0_7_rdata_data_data,data_arrays_0_6_rdata_data_data,data_arrays_0_5_rdata_data_data,data_arrays_0_4_rdata_data_data}; 
  assign lo={data_arrays_0_11_rdata_data_data,data_arrays_0_10_rdata_data_data,data_arrays_0_9_rdata_data_data,data_arrays_0_8_rdata_data_data}; 
  assign hi={data_arrays_0_15_rdata_data_data,data_arrays_0_14_rdata_data_data,data_arrays_0_13_rdata_data_data,data_arrays_0_12_rdata_data_data}; 
  assign lo_1={data_arrays_0_19_rdata_data_data,data_arrays_0_18_rdata_data_data,data_arrays_0_17_rdata_data_data,data_arrays_0_16_rdata_data_data}; 
  assign hi_1={data_arrays_0_23_rdata_data_data,data_arrays_0_22_rdata_data_data,data_arrays_0_21_rdata_data_data,data_arrays_0_20_rdata_data_data}; 
  assign lo_2={data_arrays_0_27_rdata_data_data,data_arrays_0_26_rdata_data_data,data_arrays_0_25_rdata_data_data,data_arrays_0_24_rdata_data_data}; 
  assign hi_2={data_arrays_0_31_rdata_data_data,data_arrays_0_30_rdata_data_data,data_arrays_0_29_rdata_data_data,data_arrays_0_28_rdata_data_data}; 
  assign io_resp_0={rdata_hi,rdata_lo}; 
  assign io_resp_1={hi,lo}; 
  assign io_resp_2={hi_1,lo_1}; 
  assign io_resp_3={hi_2,lo_2}; 
  assign DCacheDataArray_covSum=30'h0; 
  assign io_covSum=DCacheDataArray_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (data_arrays_0_0_rdata_MPORT_en&data_arrays_0_0_rdata_MPORT_mask)
            begin 
              data_arrays_0_0 [data_arrays_0_0_rdata_MPORT_addr]<=data_arrays_0_0_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_0_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_0_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_0_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_0_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_1_rdata_MPORT_en&data_arrays_0_1_rdata_MPORT_mask)
            begin 
              data_arrays_0_1 [data_arrays_0_1_rdata_MPORT_addr]<=data_arrays_0_1_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_1_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_1_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_1_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_1_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_2_rdata_MPORT_en&data_arrays_0_2_rdata_MPORT_mask)
            begin 
              data_arrays_0_2 [data_arrays_0_2_rdata_MPORT_addr]<=data_arrays_0_2_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_2_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_2_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_2_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_2_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_3_rdata_MPORT_en&data_arrays_0_3_rdata_MPORT_mask)
            begin 
              data_arrays_0_3 [data_arrays_0_3_rdata_MPORT_addr]<=data_arrays_0_3_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_3_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_3_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_3_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_3_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_4_rdata_MPORT_en&data_arrays_0_4_rdata_MPORT_mask)
            begin 
              data_arrays_0_4 [data_arrays_0_4_rdata_MPORT_addr]<=data_arrays_0_4_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_4_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_4_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_4_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_4_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_5_rdata_MPORT_en&data_arrays_0_5_rdata_MPORT_mask)
            begin 
              data_arrays_0_5 [data_arrays_0_5_rdata_MPORT_addr]<=data_arrays_0_5_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_5_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_5_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_5_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_5_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_6_rdata_MPORT_en&data_arrays_0_6_rdata_MPORT_mask)
            begin 
              data_arrays_0_6 [data_arrays_0_6_rdata_MPORT_addr]<=data_arrays_0_6_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_6_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_6_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_6_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_6_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_7_rdata_MPORT_en&data_arrays_0_7_rdata_MPORT_mask)
            begin 
              data_arrays_0_7 [data_arrays_0_7_rdata_MPORT_addr]<=data_arrays_0_7_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_7_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_7_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_7_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_7_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_8_rdata_MPORT_en&data_arrays_0_8_rdata_MPORT_mask)
            begin 
              data_arrays_0_8 [data_arrays_0_8_rdata_MPORT_addr]<=data_arrays_0_8_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_8_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_8_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_8_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_8_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_9_rdata_MPORT_en&data_arrays_0_9_rdata_MPORT_mask)
            begin 
              data_arrays_0_9 [data_arrays_0_9_rdata_MPORT_addr]<=data_arrays_0_9_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_9_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_9_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_9_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_9_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_10_rdata_MPORT_en&data_arrays_0_10_rdata_MPORT_mask)
            begin 
              data_arrays_0_10 [data_arrays_0_10_rdata_MPORT_addr]<=data_arrays_0_10_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_10_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_10_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_10_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_10_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_11_rdata_MPORT_en&data_arrays_0_11_rdata_MPORT_mask)
            begin 
              data_arrays_0_11 [data_arrays_0_11_rdata_MPORT_addr]<=data_arrays_0_11_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_11_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_11_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_11_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_11_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_12_rdata_MPORT_en&data_arrays_0_12_rdata_MPORT_mask)
            begin 
              data_arrays_0_12 [data_arrays_0_12_rdata_MPORT_addr]<=data_arrays_0_12_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_12_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_12_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_12_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_12_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_13_rdata_MPORT_en&data_arrays_0_13_rdata_MPORT_mask)
            begin 
              data_arrays_0_13 [data_arrays_0_13_rdata_MPORT_addr]<=data_arrays_0_13_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_13_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_13_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_13_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_13_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_14_rdata_MPORT_en&data_arrays_0_14_rdata_MPORT_mask)
            begin 
              data_arrays_0_14 [data_arrays_0_14_rdata_MPORT_addr]<=data_arrays_0_14_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_14_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_14_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_14_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_14_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_15_rdata_MPORT_en&data_arrays_0_15_rdata_MPORT_mask)
            begin 
              data_arrays_0_15 [data_arrays_0_15_rdata_MPORT_addr]<=data_arrays_0_15_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_15_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_15_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_15_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_15_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_16_rdata_MPORT_en&data_arrays_0_16_rdata_MPORT_mask)
            begin 
              data_arrays_0_16 [data_arrays_0_16_rdata_MPORT_addr]<=data_arrays_0_16_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_16_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_16_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_16_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_16_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_17_rdata_MPORT_en&data_arrays_0_17_rdata_MPORT_mask)
            begin 
              data_arrays_0_17 [data_arrays_0_17_rdata_MPORT_addr]<=data_arrays_0_17_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_17_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_17_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_17_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_17_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_18_rdata_MPORT_en&data_arrays_0_18_rdata_MPORT_mask)
            begin 
              data_arrays_0_18 [data_arrays_0_18_rdata_MPORT_addr]<=data_arrays_0_18_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_18_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_18_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_18_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_18_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_19_rdata_MPORT_en&data_arrays_0_19_rdata_MPORT_mask)
            begin 
              data_arrays_0_19 [data_arrays_0_19_rdata_MPORT_addr]<=data_arrays_0_19_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_19_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_19_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_19_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_19_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_20_rdata_MPORT_en&data_arrays_0_20_rdata_MPORT_mask)
            begin 
              data_arrays_0_20 [data_arrays_0_20_rdata_MPORT_addr]<=data_arrays_0_20_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_20_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_20_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_20_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_20_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_21_rdata_MPORT_en&data_arrays_0_21_rdata_MPORT_mask)
            begin 
              data_arrays_0_21 [data_arrays_0_21_rdata_MPORT_addr]<=data_arrays_0_21_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_21_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_21_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_21_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_21_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_22_rdata_MPORT_en&data_arrays_0_22_rdata_MPORT_mask)
            begin 
              data_arrays_0_22 [data_arrays_0_22_rdata_MPORT_addr]<=data_arrays_0_22_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_22_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_22_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_22_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_22_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_23_rdata_MPORT_en&data_arrays_0_23_rdata_MPORT_mask)
            begin 
              data_arrays_0_23 [data_arrays_0_23_rdata_MPORT_addr]<=data_arrays_0_23_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_23_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_23_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_23_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_23_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_24_rdata_MPORT_en&data_arrays_0_24_rdata_MPORT_mask)
            begin 
              data_arrays_0_24 [data_arrays_0_24_rdata_MPORT_addr]<=data_arrays_0_24_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_24_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_24_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_24_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_24_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_25_rdata_MPORT_en&data_arrays_0_25_rdata_MPORT_mask)
            begin 
              data_arrays_0_25 [data_arrays_0_25_rdata_MPORT_addr]<=data_arrays_0_25_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_25_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_25_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_25_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_25_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_26_rdata_MPORT_en&data_arrays_0_26_rdata_MPORT_mask)
            begin 
              data_arrays_0_26 [data_arrays_0_26_rdata_MPORT_addr]<=data_arrays_0_26_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_26_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_26_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_26_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_26_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_27_rdata_MPORT_en&data_arrays_0_27_rdata_MPORT_mask)
            begin 
              data_arrays_0_27 [data_arrays_0_27_rdata_MPORT_addr]<=data_arrays_0_27_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_27_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_27_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_27_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_27_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_28_rdata_MPORT_en&data_arrays_0_28_rdata_MPORT_mask)
            begin 
              data_arrays_0_28 [data_arrays_0_28_rdata_MPORT_addr]<=data_arrays_0_28_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_28_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_28_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_28_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_28_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_29_rdata_MPORT_en&data_arrays_0_29_rdata_MPORT_mask)
            begin 
              data_arrays_0_29 [data_arrays_0_29_rdata_MPORT_addr]<=data_arrays_0_29_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_29_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_29_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_29_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_29_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_30_rdata_MPORT_en&data_arrays_0_30_rdata_MPORT_mask)
            begin 
              data_arrays_0_30 [data_arrays_0_30_rdata_MPORT_addr]<=data_arrays_0_30_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_30_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_30_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_30_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_30_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
         if (data_arrays_0_31_rdata_MPORT_en&data_arrays_0_31_rdata_MPORT_mask)
            begin 
              data_arrays_0_31 [data_arrays_0_31_rdata_MPORT_addr]<=data_arrays_0_31_rdata_MPORT_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_31_rdata_data_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_31_rdata_data_en_pipe_0 <=io_req_valid&~io_req_bits_write;
            end 
         if (metaReset)
            begin 
              data_arrays_0_31_rdata_data_addr_pipe_0 <=9'h0;
            end 
          else 
            if (io_req_valid&~io_req_bits_write)
               begin 
                 data_arrays_0_31_rdata_data_addr_pipe_0 <=io_req_bits_addr[11:3];
               end 
       end
  
endmodule
 
module DCacheModuleImpl_Anon_2 (
  input io_in_0_valid,
  input [11:0] io_in_0_bits_addr,
  input io_in_0_bits_write,
  input [63:0] io_in_0_bits_wdata,
  input [7:0] io_in_0_bits_eccMask,
  input [3:0] io_in_0_bits_way_en,
  output io_in_1_ready,
  input io_in_1_valid,
  input [11:0] io_in_1_bits_addr,
  input io_in_1_bits_write,
  input [63:0] io_in_1_bits_wdata,
  input [3:0] io_in_1_bits_way_en,
  output io_in_2_ready,
  input io_in_2_valid,
  input [11:0] io_in_2_bits_addr,
  input [63:0] io_in_2_bits_wdata,
  output io_in_3_ready,
  input io_in_3_valid,
  input [11:0] io_in_3_bits_addr,
  input [63:0] io_in_3_bits_wdata,
  input io_in_3_bits_wordMask,
  output io_out_valid,
  output [11:0] io_out_bits_addr,
  output io_out_bits_write,
  output [63:0] io_out_bits_wdata,
  output [7:0] io_out_bits_eccMask,
  output [3:0] io_out_bits_way_en,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [63:0] _GEN_4 ;  
   wire [11:0] _GEN_6 ;  
   wire [3:0] _GEN_8 ;  
   wire [63:0] _GEN_11 ;  
   wire _GEN_12 ;  
   wire [11:0] _GEN_13 ;  
   wire _grant_T ;  
   wire _grant_T_1 ;  
   wire grant_3 ;  
   wire [29:0] DCacheModuleImpl_Anon_2_covSum ;  
  assign _GEN_4=io_in_2_valid ? io_in_2_bits_wdata:io_in_3_bits_wdata; 
  assign _GEN_6=io_in_2_valid ? io_in_2_bits_addr:io_in_3_bits_addr; 
  assign _GEN_8=io_in_1_valid ? io_in_1_bits_way_en:4'hf; 
  assign _GEN_11=io_in_1_valid ? io_in_1_bits_wdata:_GEN_4; 
  assign _GEN_12=io_in_1_valid&io_in_1_bits_write; 
  assign _GEN_13=io_in_1_valid ? io_in_1_bits_addr:_GEN_6; 
  assign _grant_T=io_in_0_valid|io_in_1_valid; 
  assign _grant_T_1=_grant_T|io_in_2_valid; 
  assign grant_3=~_grant_T_1; 
  assign io_in_1_ready=~io_in_0_valid; 
  assign io_in_2_ready=~_grant_T; 
  assign io_in_3_ready=~_grant_T_1; 
  assign io_out_valid=~grant_3|io_in_3_valid; 
  assign io_out_bits_addr=io_in_0_valid ? io_in_0_bits_addr:_GEN_13; 
  assign io_out_bits_write=io_in_0_valid ? io_in_0_bits_write:_GEN_12; 
  assign io_out_bits_wdata=io_in_0_valid ? io_in_0_bits_wdata:_GEN_11; 
  assign io_out_bits_eccMask=io_in_0_valid ? io_in_0_bits_eccMask:8'hff; 
  assign io_out_bits_way_en=io_in_0_valid ? io_in_0_bits_way_en:_GEN_8; 
  assign DCacheModuleImpl_Anon_2_covSum=30'h0; 
  assign io_covSum=DCacheModuleImpl_Anon_2_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module AMOALU (
  input [7:0] io_mask,
  input [4:0] io_cmd,
  input [63:0] io_lhs,
  input [63:0] io_rhs,
  output [63:0] io_out,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire _max_T ;  
   wire _max_T_1 ;  
   wire max ;  
   wire _min_T ;  
   wire _min_T_1 ;  
   wire min ;  
   wire add ;  
   wire _logic_and_T ;  
   wire _logic_and_T_1 ;  
   wire logic_and ;  
   wire _logic_xor_T ;  
   wire logic_xor ;  
   wire [31:0] _adder_out_mask_T_2 ;  
   wire [63:0] _adder_out_mask_T_3 ;  
   wire [63:0] adder_out_mask ;  
   wire [63:0] _adder_out_T ;  
   wire [63:0] _adder_out_T_1 ;  
   wire [63:0] adder_out ;  
   wire [4:0] _less_signed_T ;  
   wire less_signed ;  
   wire _less_T_3 ;  
   wire _less_T_6 ;  
   wire _less_T_9 ;  
   wire _less_T_12 ;  
   wire _less_T_13 ;  
   wire _less_T_14 ;  
   wire _less_T_17 ;  
   wire _less_T_18 ;  
   wire _less_T_22 ;  
   wire _less_T_28 ;  
   wire _less_T_29 ;  
   wire less ;  
   wire _minmax_T ;  
   wire [63:0] minmax ;  
   wire [63:0] _logic_T ;  
   wire [63:0] _logic_T_1 ;  
   wire [63:0] _logic_T_2 ;  
   wire [63:0] _logic_T_3 ;  
   wire [63:0] logic_ ;  
   wire _out_T ;  
   wire [63:0] _out_T_1 ;  
   wire [63:0] out ;  
   wire [7:0] wmask_lo_lo_lo ;  
   wire [7:0] wmask_lo_lo_hi ;  
   wire [7:0] wmask_lo_hi_lo ;  
   wire [7:0] wmask_lo_hi_hi ;  
   wire [7:0] wmask_hi_lo_lo ;  
   wire [7:0] wmask_hi_lo_hi ;  
   wire [7:0] wmask_hi_hi_lo ;  
   wire [7:0] wmask_hi_hi_hi ;  
   wire [63:0] wmask ;  
   wire [63:0] _io_out_T ;  
   wire [63:0] _io_out_T_2 ;  
   wire [29:0] AMOALU_covSum ;  
  assign _max_T=io_cmd==5'hd; 
  assign _max_T_1=io_cmd==5'hf; 
  assign max=_max_T|_max_T_1; 
  assign _min_T=io_cmd==5'hc; 
  assign _min_T_1=io_cmd==5'he; 
  assign min=_min_T|_min_T_1; 
  assign add=io_cmd==5'h8; 
  assign _logic_and_T=io_cmd==5'ha; 
  assign _logic_and_T_1=io_cmd==5'hb; 
  assign logic_and=_logic_and_T|_logic_and_T_1; 
  assign _logic_xor_T=io_cmd==5'h9; 
  assign logic_xor=_logic_xor_T|_logic_and_T; 
  assign _adder_out_mask_T_2={~io_mask[3],31'h0}; 
  assign _adder_out_mask_T_3={32'b0,_adder_out_mask_T_2}; 
  assign adder_out_mask=~_adder_out_mask_T_3; 
  assign _adder_out_T=io_lhs&adder_out_mask; 
  assign _adder_out_T_1=io_rhs&adder_out_mask; 
  assign adder_out=_adder_out_T+_adder_out_T_1; 
  assign _less_signed_T=io_cmd&5'h2; 
  assign less_signed=_less_signed_T==5'h0; 
  assign _less_T_3=io_lhs[63]==io_rhs[63]; 
  assign _less_T_6=io_lhs[63:32]<io_rhs[63:32]; 
  assign _less_T_9=io_lhs[63:32]==io_rhs[63:32]; 
  assign _less_T_12=io_lhs[31:0]<io_rhs[31:0]; 
  assign _less_T_13=_less_T_9&_less_T_12; 
  assign _less_T_14=_less_T_6|_less_T_13; 
  assign _less_T_17=less_signed ? io_lhs[63]:io_rhs[63]; 
  assign _less_T_18=_less_T_3 ? _less_T_14:_less_T_17; 
  assign _less_T_22=io_lhs[31]==io_rhs[31]; 
  assign _less_T_28=less_signed ? io_lhs[31]:io_rhs[31]; 
  assign _less_T_29=_less_T_22 ? _less_T_12:_less_T_28; 
  assign less=io_mask[4] ? _less_T_18:_less_T_29; 
  assign _minmax_T=less ? min:max; 
  assign minmax=_minmax_T ? io_lhs:io_rhs; 
  assign _logic_T=io_lhs&io_rhs; 
  assign _logic_T_1=logic_and ? _logic_T:64'h0; 
  assign _logic_T_2=io_lhs^io_rhs; 
  assign _logic_T_3=logic_xor ? _logic_T_2:64'h0; 
  assign logic_=_logic_T_1|_logic_T_3; 
  assign _out_T=logic_and|logic_xor; 
  assign _out_T_1=_out_T ? logic_:minmax; 
  assign out=add ? adder_out:_out_T_1; 
  assign wmask_lo_lo_lo=io_mask[0] ? 8'hff:8'h0; 
  assign wmask_lo_lo_hi=io_mask[1] ? 8'hff:8'h0; 
  assign wmask_lo_hi_lo=io_mask[2] ? 8'hff:8'h0; 
  assign wmask_lo_hi_hi=io_mask[3] ? 8'hff:8'h0; 
  assign wmask_hi_lo_lo=io_mask[4] ? 8'hff:8'h0; 
  assign wmask_hi_lo_hi=io_mask[5] ? 8'hff:8'h0; 
  assign wmask_hi_hi_lo=io_mask[6] ? 8'hff:8'h0; 
  assign wmask_hi_hi_hi=io_mask[7] ? 8'hff:8'h0; 
  assign wmask={wmask_hi_hi_hi,wmask_hi_hi_lo,wmask_hi_lo_hi,wmask_hi_lo_lo,wmask_lo_hi_hi,wmask_lo_hi_lo,wmask_lo_lo_hi,wmask_lo_lo_lo}; 
  assign _io_out_T=wmask&out; 
  assign _io_out_T_2=~wmask&io_lhs; 
  assign io_out=_io_out_T|_io_out_T_2; 
  assign AMOALU_covSum=30'h0; 
  assign io_covSum=AMOALU_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module ICache (
  input clock,
  input reset,
  input auto_master_out_a_ready,
  output auto_master_out_a_valid,
  output [31:0] auto_master_out_a_bits_address,
  input auto_master_out_d_valid,
  input [2:0] auto_master_out_d_bits_opcode,
  input [3:0] auto_master_out_d_bits_size,
  input [63:0] auto_master_out_d_bits_data,
  input auto_master_out_d_bits_corrupt,
  output io_req_ready,
  input io_req_valid,
  input [38:0] io_req_bits_addr,
  input [31:0] io_s1_paddr,
  input io_s1_kill,
  input io_s2_kill,
  output io_resp_valid,
  output [31:0] io_resp_bits_data,
  output io_resp_bits_replay,
  output io_resp_bits_ae,
  input io_invalidate,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input repl_way_v0_prng_halt) ; 
   wire repl_way_v0_prng_clock ;  
   wire repl_way_v0_prng_reset ;  
   wire repl_way_v0_prng_io_increment ;  
   wire repl_way_v0_prng_io_out_0 ;  
   wire repl_way_v0_prng_io_out_1 ;  
   wire repl_way_v0_prng_io_out_2 ;  
   wire repl_way_v0_prng_io_out_3 ;  
   wire repl_way_v0_prng_io_out_4 ;  
   wire repl_way_v0_prng_io_out_5 ;  
   wire repl_way_v0_prng_io_out_6 ;  
   wire repl_way_v0_prng_io_out_7 ;  
   wire repl_way_v0_prng_io_out_8 ;  
   wire repl_way_v0_prng_io_out_9 ;  
   wire repl_way_v0_prng_io_out_10 ;  
   wire repl_way_v0_prng_io_out_11 ;  
   wire repl_way_v0_prng_io_out_12 ;  
   wire repl_way_v0_prng_io_out_13 ;  
   wire repl_way_v0_prng_io_out_14 ;  
   wire repl_way_v0_prng_io_out_15 ;  
   wire [29:0] repl_way_v0_prng_io_covSum ;  
   wire repl_way_v0_prng_metaAssert ;  
   wire repl_way_v0_prng_metaReset ;  
   reg [20:0] tag_array_0[0:63] ;  
   reg [31:0] _RAND_0 ;  
   wire [20:0] tag_array_0_tag_rdata_data ;  
   wire [5:0] tag_array_0_tag_rdata_addr ;  
   wire [20:0] tag_array_0_MPORT_data ;  
   wire [5:0] tag_array_0_MPORT_addr ;  
   wire tag_array_0_MPORT_mask ;  
   wire tag_array_0_MPORT_en ;  
   reg tag_array_0_tag_rdata_en_pipe_0 ;  
   reg [31:0] _RAND_1 ;  
   reg [5:0] tag_array_0_tag_rdata_addr_pipe_0 ;  
   reg [31:0] _RAND_2 ;  
   reg [20:0] tag_array_1[0:63] ;  
   reg [31:0] _RAND_3 ;  
   wire [20:0] tag_array_1_tag_rdata_data ;  
   wire [5:0] tag_array_1_tag_rdata_addr ;  
   wire [20:0] tag_array_1_MPORT_data ;  
   wire [5:0] tag_array_1_MPORT_addr ;  
   wire tag_array_1_MPORT_mask ;  
   wire tag_array_1_MPORT_en ;  
   reg tag_array_1_tag_rdata_en_pipe_0 ;  
   reg [31:0] _RAND_4 ;  
   reg [5:0] tag_array_1_tag_rdata_addr_pipe_0 ;  
   reg [31:0] _RAND_5 ;  
   reg [20:0] tag_array_2[0:63] ;  
   reg [31:0] _RAND_6 ;  
   wire [20:0] tag_array_2_tag_rdata_data ;  
   wire [5:0] tag_array_2_tag_rdata_addr ;  
   wire [20:0] tag_array_2_MPORT_data ;  
   wire [5:0] tag_array_2_MPORT_addr ;  
   wire tag_array_2_MPORT_mask ;  
   wire tag_array_2_MPORT_en ;  
   reg tag_array_2_tag_rdata_en_pipe_0 ;  
   reg [31:0] _RAND_7 ;  
   reg [5:0] tag_array_2_tag_rdata_addr_pipe_0 ;  
   reg [31:0] _RAND_8 ;  
   reg [20:0] tag_array_3[0:63] ;  
   reg [31:0] _RAND_9 ;  
   wire [20:0] tag_array_3_tag_rdata_data ;  
   wire [5:0] tag_array_3_tag_rdata_addr ;  
   wire [20:0] tag_array_3_MPORT_data ;  
   wire [5:0] tag_array_3_MPORT_addr ;  
   wire tag_array_3_MPORT_mask ;  
   wire tag_array_3_MPORT_en ;  
   reg tag_array_3_tag_rdata_en_pipe_0 ;  
   reg [31:0] _RAND_10 ;  
   reg [5:0] tag_array_3_tag_rdata_addr_pipe_0 ;  
   reg [31:0] _RAND_11 ;  
   reg [31:0] data_arrays_0_0[0:511] ;  
   reg [31:0] _RAND_12 ;  
   wire [31:0] data_arrays_0_0_dout_data ;  
   wire [8:0] data_arrays_0_0_dout_addr ;  
   wire [31:0] data_arrays_0_0_MPORT_1_data ;  
   wire [8:0] data_arrays_0_0_MPORT_1_addr ;  
   wire data_arrays_0_0_MPORT_1_mask ;  
   wire data_arrays_0_0_MPORT_1_en ;  
   reg data_arrays_0_0_dout_en_pipe_0 ;  
   reg [31:0] _RAND_13 ;  
   reg [8:0] data_arrays_0_0_dout_addr_pipe_0 ;  
   reg [31:0] _RAND_14 ;  
   reg [31:0] data_arrays_0_1[0:511] ;  
   reg [31:0] _RAND_15 ;  
   wire [31:0] data_arrays_0_1_dout_data ;  
   wire [8:0] data_arrays_0_1_dout_addr ;  
   wire [31:0] data_arrays_0_1_MPORT_1_data ;  
   wire [8:0] data_arrays_0_1_MPORT_1_addr ;  
   wire data_arrays_0_1_MPORT_1_mask ;  
   wire data_arrays_0_1_MPORT_1_en ;  
   reg data_arrays_0_1_dout_en_pipe_0 ;  
   reg [31:0] _RAND_16 ;  
   reg [8:0] data_arrays_0_1_dout_addr_pipe_0 ;  
   reg [31:0] _RAND_17 ;  
   reg [31:0] data_arrays_0_2[0:511] ;  
   reg [31:0] _RAND_18 ;  
   wire [31:0] data_arrays_0_2_dout_data ;  
   wire [8:0] data_arrays_0_2_dout_addr ;  
   wire [31:0] data_arrays_0_2_MPORT_1_data ;  
   wire [8:0] data_arrays_0_2_MPORT_1_addr ;  
   wire data_arrays_0_2_MPORT_1_mask ;  
   wire data_arrays_0_2_MPORT_1_en ;  
   reg data_arrays_0_2_dout_en_pipe_0 ;  
   reg [31:0] _RAND_19 ;  
   reg [8:0] data_arrays_0_2_dout_addr_pipe_0 ;  
   reg [31:0] _RAND_20 ;  
   reg [31:0] data_arrays_0_3[0:511] ;  
   reg [31:0] _RAND_21 ;  
   wire [31:0] data_arrays_0_3_dout_data ;  
   wire [8:0] data_arrays_0_3_dout_addr ;  
   wire [31:0] data_arrays_0_3_MPORT_1_data ;  
   wire [8:0] data_arrays_0_3_MPORT_1_addr ;  
   wire data_arrays_0_3_MPORT_1_mask ;  
   wire data_arrays_0_3_MPORT_1_en ;  
   reg data_arrays_0_3_dout_en_pipe_0 ;  
   reg [31:0] _RAND_22 ;  
   reg [8:0] data_arrays_0_3_dout_addr_pipe_0 ;  
   reg [31:0] _RAND_23 ;  
   reg [31:0] data_arrays_1_0[0:511] ;  
   reg [31:0] _RAND_24 ;  
   wire [31:0] data_arrays_1_0_dout_1_data ;  
   wire [8:0] data_arrays_1_0_dout_1_addr ;  
   wire [31:0] data_arrays_1_0_MPORT_2_data ;  
   wire [8:0] data_arrays_1_0_MPORT_2_addr ;  
   wire data_arrays_1_0_MPORT_2_mask ;  
   wire data_arrays_1_0_MPORT_2_en ;  
   reg data_arrays_1_0_dout_1_en_pipe_0 ;  
   reg [31:0] _RAND_25 ;  
   reg [8:0] data_arrays_1_0_dout_1_addr_pipe_0 ;  
   reg [31:0] _RAND_26 ;  
   reg [31:0] data_arrays_1_1[0:511] ;  
   reg [31:0] _RAND_27 ;  
   wire [31:0] data_arrays_1_1_dout_1_data ;  
   wire [8:0] data_arrays_1_1_dout_1_addr ;  
   wire [31:0] data_arrays_1_1_MPORT_2_data ;  
   wire [8:0] data_arrays_1_1_MPORT_2_addr ;  
   wire data_arrays_1_1_MPORT_2_mask ;  
   wire data_arrays_1_1_MPORT_2_en ;  
   reg data_arrays_1_1_dout_1_en_pipe_0 ;  
   reg [31:0] _RAND_28 ;  
   reg [8:0] data_arrays_1_1_dout_1_addr_pipe_0 ;  
   reg [31:0] _RAND_29 ;  
   reg [31:0] data_arrays_1_2[0:511] ;  
   reg [31:0] _RAND_30 ;  
   wire [31:0] data_arrays_1_2_dout_1_data ;  
   wire [8:0] data_arrays_1_2_dout_1_addr ;  
   wire [31:0] data_arrays_1_2_MPORT_2_data ;  
   wire [8:0] data_arrays_1_2_MPORT_2_addr ;  
   wire data_arrays_1_2_MPORT_2_mask ;  
   wire data_arrays_1_2_MPORT_2_en ;  
   reg data_arrays_1_2_dout_1_en_pipe_0 ;  
   reg [31:0] _RAND_31 ;  
   reg [8:0] data_arrays_1_2_dout_1_addr_pipe_0 ;  
   reg [31:0] _RAND_32 ;  
   reg [31:0] data_arrays_1_3[0:511] ;  
   reg [31:0] _RAND_33 ;  
   wire [31:0] data_arrays_1_3_dout_1_data ;  
   wire [8:0] data_arrays_1_3_dout_1_addr ;  
   wire [31:0] data_arrays_1_3_MPORT_2_data ;  
   wire [8:0] data_arrays_1_3_MPORT_2_addr ;  
   wire data_arrays_1_3_MPORT_2_mask ;  
   wire data_arrays_1_3_MPORT_2_en ;  
   reg data_arrays_1_3_dout_1_en_pipe_0 ;  
   reg [31:0] _RAND_34 ;  
   reg [8:0] data_arrays_1_3_dout_1_addr_pipe_0 ;  
   reg [31:0] _RAND_35 ;  
   wire s0_valid ;  
   reg s1_valid ;  
   reg [31:0] _RAND_36 ;  
   reg [255:0] vb_array ;  
   reg [255:0] _RAND_37 ;  
   wire [5:0] s1_vb_lo ;  
   wire [6:0] _s1_vb_T ;  
   wire [255:0] _s1_vb_T_1 ;  
   wire s1_vb ;  
   wire [19:0] tag ;  
   wire [19:0] s1_tag ;  
   wire _tagMatch_T ;  
   wire tagMatch ;  
   wire [6:0] _s1_vb_T_4 ;  
   wire [255:0] _s1_vb_T_5 ;  
   wire s1_vb_1 ;  
   wire [19:0] tag_1 ;  
   wire _tagMatch_T_1 ;  
   wire tagMatch_1 ;  
   wire _s1_hit_T ;  
   wire [7:0] _s1_vb_T_8 ;  
   wire [255:0] _s1_vb_T_9 ;  
   wire s1_vb_2 ;  
   wire [19:0] tag_2 ;  
   wire _tagMatch_T_2 ;  
   wire tagMatch_2 ;  
   wire _s1_hit_T_1 ;  
   wire [7:0] _s1_vb_T_12 ;  
   wire [255:0] _s1_vb_T_13 ;  
   wire s1_vb_3 ;  
   wire [19:0] tag_3 ;  
   wire _tagMatch_T_3 ;  
   wire tagMatch_3 ;  
   wire _s2_valid_T_1 ;  
   reg s2_valid ;  
   reg [31:0] _RAND_38 ;  
   reg s2_hit ;  
   reg [31:0] _RAND_39 ;  
   reg invalidated ;  
   reg [31:0] _RAND_40 ;  
   reg refill_valid ;  
   reg [31:0] _RAND_41 ;  
   wire _s2_miss_T_1 ;  
   wire s2_miss ;  
   reg s2_request_refill_REG ;  
   reg [31:0] _RAND_42 ;  
   wire s2_request_refill ;  
   wire refill_fire ;  
   wire _s1_can_request_refill_T ;  
   wire s1_can_request_refill ;  
   wire _refill_paddr_T ;  
   reg [31:0] refill_paddr ;  
   reg [31:0] _RAND_43 ;  
   wire [19:0] refill_tag ;  
   wire [5:0] refill_idx ;  
   wire refill_one_beat_opdata ;  
   wire refill_one_beat ;  
   wire [26:0] _beats1_decode_T_1 ;  
   wire [8:0] beats1_decode ;  
   wire [8:0] beats1 ;  
   reg [8:0] counter ;  
   reg [31:0] _RAND_44 ;  
   wire [8:0] counter1 ;  
   wire first ;  
   wire _last_T ;  
   wire _last_T_1 ;  
   wire last ;  
   wire d_done ;  
   wire [8:0] refill_cnt ;  
   wire refill_done ;  
   wire [7:0] repl_way_v0_lo ;  
   wire [15:0] _repl_way_v0_T ;  
   wire [1:0] repl_way_v0 ;  
   wire [7:0] _repl_way_T ;  
   reg accruedRefillError ;  
   reg [31:0] _RAND_45 ;  
   wire _refillError_T ;  
   wire _refillError_T_1 ;  
   wire refillError ;  
   wire _vb_array_T_2 ;  
   wire [255:0] _vb_array_T_3 ;  
   wire [255:0] _vb_array_T_4 ;  
   wire [255:0] _vb_array_T_6 ;  
   wire s2_tag_disparity ;  
   wire _T_40 ;  
   wire invalidate ;  
   wire _GEN_30 ;  
   wire tl_error ;  
   wire s1_tl_error_0 ;  
   wire tl_error_1 ;  
   wire s1_tl_error_1 ;  
   wire tl_error_2 ;  
   wire s1_tl_error_2 ;  
   wire tl_error_3 ;  
   wire s1_tl_error_3 ;  
   wire [1:0] _T_15 ;  
   wire [1:0] _T_17 ;  
   wire [2:0] _T_19 ;  
   wire _T_21 ;  
   wire _T_22 ;  
   wire _T_24 ;  
   wire s0_ren ;  
   wire wen ;  
   wire [8:0] _mem_idx_T ;  
   wire [8:0] _mem_idx_T_1 ;  
   wire [31:0] _GEN_54 ;  
   wire [31:0] _GEN_55 ;  
   wire [31:0] _GEN_56 ;  
   wire [31:0] _GEN_57 ;  
   wire s0_ren_1 ;  
   reg s2_tag_hit_0 ;  
   reg [31:0] _RAND_46 ;  
   reg s2_tag_hit_1 ;  
   reg [31:0] _RAND_47 ;  
   reg s2_tag_hit_2 ;  
   reg [31:0] _RAND_48 ;  
   reg s2_tag_hit_3 ;  
   reg [31:0] _RAND_49 ;  
   reg [31:0] s2_dout_0 ;  
   reg [31:0] _RAND_50 ;  
   reg [31:0] s2_dout_1 ;  
   reg [31:0] _RAND_51 ;  
   reg [31:0] s2_dout_2 ;  
   reg [31:0] _RAND_52 ;  
   reg [31:0] s2_dout_3 ;  
   reg [31:0] _RAND_53 ;  
   wire [31:0] _s2_way_mux_T ;  
   wire [31:0] _s2_way_mux_T_1 ;  
   wire [31:0] _s2_way_mux_T_2 ;  
   wire [31:0] _s2_way_mux_T_3 ;  
   wire [31:0] _s2_way_mux_T_4 ;  
   wire [31:0] _s2_way_mux_T_5 ;  
   wire [3:0] _s2_tl_error_T ;  
   wire _s2_tl_error_T_1 ;  
   reg s2_tl_error ;  
   reg [31:0] _RAND_54 ;  
   wire _GEN_101 ;  
   reg [5:0] ICache_state ;  
   reg [31:0] _RAND_55 ;  
   reg ICache_cov[0:63] ;  
   reg [31:0] _RAND_56 ;  
   wire ICache_cov_read_data ;  
   wire [5:0] ICache_cov_read_addr ;  
   wire ICache_cov_write_data ;  
   wire [5:0] ICache_cov_write_addr ;  
   wire ICache_cov_write_mask ;  
   wire ICache_cov_write_en ;  
   reg [29:0] ICache_covSum ;  
   reg [31:0] _RAND_57 ;  
   wire s2_valid_shl ;  
   wire [5:0] s2_valid_pad ;  
   wire [1:0] s1_valid_shl ;  
   wire [5:0] s1_valid_pad ;  
   wire [2:0] refill_valid_shl ;  
   wire [5:0] refill_valid_pad ;  
   wire [3:0] invalidated_shl ;  
   wire [5:0] invalidated_pad ;  
   wire [4:0] s2_hit_shl ;  
   wire [5:0] s2_hit_pad ;  
   wire [5:0] s2_tag_hit_0_shl ;  
   wire [5:0] s2_tag_hit_0_pad ;  
   wire [5:0] s2_tag_hit_1_shl ;  
   wire [5:0] s2_tag_hit_1_pad ;  
   wire [5:0] s2_tag_hit_2_shl ;  
   wire [5:0] s2_tag_hit_2_pad ;  
   wire [5:0] s2_tag_hit_3_shl ;  
   wire [5:0] s2_tag_hit_3_pad ;  
   wire [5:0] ICache_xor3 ;  
   wire [5:0] ICache_xor4 ;  
   wire [5:0] ICache_xor1 ;  
   wire [5:0] ICache_xor5 ;  
   wire [5:0] ICache_xor14 ;  
   wire [5:0] ICache_xor6 ;  
   wire [5:0] ICache_xor2 ;  
   wire [5:0] ICache_xor0 ;  
   wire [29:0] repl_way_v0_prng_sum ;  
   wire stopEn0 ;  
   wire repl_way_v0_prng_metaAssert_wire ;  
   wire ICache_or0 ;  
   reg ICache_metaAssert ;  
   reg [31:0] _RAND_58 ;  
  MaxPeriodFibonacciLFSR repl_way_v0_prng(.clock(repl_way_v0_prng_clock),.reset(repl_way_v0_prng_reset),.io_increment(repl_way_v0_prng_io_increment),.io_out_0(repl_way_v0_prng_io_out_0),.io_out_1(repl_way_v0_prng_io_out_1),.io_out_2(repl_way_v0_prng_io_out_2),.io_out_3(repl_way_v0_prng_io_out_3),.io_out_4(repl_way_v0_prng_io_out_4),.io_out_5(repl_way_v0_prng_io_out_5),.io_out_6(repl_way_v0_prng_io_out_6),.io_out_7(repl_way_v0_prng_io_out_7),.io_out_8(repl_way_v0_prng_io_out_8),.io_out_9(repl_way_v0_prng_io_out_9),.io_out_10(repl_way_v0_prng_io_out_10),.io_out_11(repl_way_v0_prng_io_out_11),.io_out_12(repl_way_v0_prng_io_out_12),.io_out_13(repl_way_v0_prng_io_out_13),.io_out_14(repl_way_v0_prng_io_out_14),.io_out_15(repl_way_v0_prng_io_out_15),.io_covSum(repl_way_v0_prng_io_covSum),.metaAssert(repl_way_v0_prng_metaAssert),.metaReset(repl_way_v0_prng_metaReset)); 
  assign tag_array_0_tag_rdata_addr=tag_array_0_tag_rdata_addr_pipe_0; 
  assign tag_array_0_tag_rdata_data=tag_array_0[tag_array_0_tag_rdata_addr]; 
  assign tag_array_0_MPORT_data={refillError,refill_tag}; 
  assign tag_array_0_MPORT_addr=refill_paddr[11:6]; 
  assign tag_array_0_MPORT_mask=repl_way_v0==2'h0; 
  assign tag_array_0_MPORT_en=refill_one_beat&d_done; 
  assign tag_array_1_tag_rdata_addr=tag_array_1_tag_rdata_addr_pipe_0; 
  assign tag_array_1_tag_rdata_data=tag_array_1[tag_array_1_tag_rdata_addr]; 
  assign tag_array_1_MPORT_data={refillError,refill_tag}; 
  assign tag_array_1_MPORT_addr=refill_paddr[11:6]; 
  assign tag_array_1_MPORT_mask=repl_way_v0==2'h1; 
  assign tag_array_1_MPORT_en=refill_one_beat&d_done; 
  assign tag_array_2_tag_rdata_addr=tag_array_2_tag_rdata_addr_pipe_0; 
  assign tag_array_2_tag_rdata_data=tag_array_2[tag_array_2_tag_rdata_addr]; 
  assign tag_array_2_MPORT_data={refillError,refill_tag}; 
  assign tag_array_2_MPORT_addr=refill_paddr[11:6]; 
  assign tag_array_2_MPORT_mask=repl_way_v0==2'h2; 
  assign tag_array_2_MPORT_en=refill_one_beat&d_done; 
  assign tag_array_3_tag_rdata_addr=tag_array_3_tag_rdata_addr_pipe_0; 
  assign tag_array_3_tag_rdata_data=tag_array_3[tag_array_3_tag_rdata_addr]; 
  assign tag_array_3_MPORT_data={refillError,refill_tag}; 
  assign tag_array_3_MPORT_addr=refill_paddr[11:6]; 
  assign tag_array_3_MPORT_mask=repl_way_v0==2'h3; 
  assign tag_array_3_MPORT_en=refill_one_beat&d_done; 
  assign data_arrays_0_0_dout_addr=data_arrays_0_0_dout_addr_pipe_0; 
  assign data_arrays_0_0_dout_data=data_arrays_0_0[data_arrays_0_0_dout_addr]; 
  assign data_arrays_0_0_MPORT_1_data=auto_master_out_d_bits_data[31:0]; 
  assign data_arrays_0_0_MPORT_1_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_0_0_MPORT_1_mask=repl_way_v0==2'h0; 
  assign data_arrays_0_0_MPORT_1_en=refill_one_beat&~invalidated; 
  assign data_arrays_0_1_dout_addr=data_arrays_0_1_dout_addr_pipe_0; 
  assign data_arrays_0_1_dout_data=data_arrays_0_1[data_arrays_0_1_dout_addr]; 
  assign data_arrays_0_1_MPORT_1_data=auto_master_out_d_bits_data[31:0]; 
  assign data_arrays_0_1_MPORT_1_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_0_1_MPORT_1_mask=repl_way_v0==2'h1; 
  assign data_arrays_0_1_MPORT_1_en=refill_one_beat&~invalidated; 
  assign data_arrays_0_2_dout_addr=data_arrays_0_2_dout_addr_pipe_0; 
  assign data_arrays_0_2_dout_data=data_arrays_0_2[data_arrays_0_2_dout_addr]; 
  assign data_arrays_0_2_MPORT_1_data=auto_master_out_d_bits_data[31:0]; 
  assign data_arrays_0_2_MPORT_1_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_0_2_MPORT_1_mask=repl_way_v0==2'h2; 
  assign data_arrays_0_2_MPORT_1_en=refill_one_beat&~invalidated; 
  assign data_arrays_0_3_dout_addr=data_arrays_0_3_dout_addr_pipe_0; 
  assign data_arrays_0_3_dout_data=data_arrays_0_3[data_arrays_0_3_dout_addr]; 
  assign data_arrays_0_3_MPORT_1_data=auto_master_out_d_bits_data[31:0]; 
  assign data_arrays_0_3_MPORT_1_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_0_3_MPORT_1_mask=repl_way_v0==2'h3; 
  assign data_arrays_0_3_MPORT_1_en=refill_one_beat&~invalidated; 
  assign data_arrays_1_0_dout_1_addr=data_arrays_1_0_dout_1_addr_pipe_0; 
  assign data_arrays_1_0_dout_1_data=data_arrays_1_0[data_arrays_1_0_dout_1_addr]; 
  assign data_arrays_1_0_MPORT_2_data=auto_master_out_d_bits_data[63:32]; 
  assign data_arrays_1_0_MPORT_2_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_1_0_MPORT_2_mask=repl_way_v0==2'h0; 
  assign data_arrays_1_0_MPORT_2_en=refill_one_beat&~invalidated; 
  assign data_arrays_1_1_dout_1_addr=data_arrays_1_1_dout_1_addr_pipe_0; 
  assign data_arrays_1_1_dout_1_data=data_arrays_1_1[data_arrays_1_1_dout_1_addr]; 
  assign data_arrays_1_1_MPORT_2_data=auto_master_out_d_bits_data[63:32]; 
  assign data_arrays_1_1_MPORT_2_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_1_1_MPORT_2_mask=repl_way_v0==2'h1; 
  assign data_arrays_1_1_MPORT_2_en=refill_one_beat&~invalidated; 
  assign data_arrays_1_2_dout_1_addr=data_arrays_1_2_dout_1_addr_pipe_0; 
  assign data_arrays_1_2_dout_1_data=data_arrays_1_2[data_arrays_1_2_dout_1_addr]; 
  assign data_arrays_1_2_MPORT_2_data=auto_master_out_d_bits_data[63:32]; 
  assign data_arrays_1_2_MPORT_2_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_1_2_MPORT_2_mask=repl_way_v0==2'h2; 
  assign data_arrays_1_2_MPORT_2_en=refill_one_beat&~invalidated; 
  assign data_arrays_1_3_dout_1_addr=data_arrays_1_3_dout_1_addr_pipe_0; 
  assign data_arrays_1_3_dout_1_data=data_arrays_1_3[data_arrays_1_3_dout_1_addr]; 
  assign data_arrays_1_3_MPORT_2_data=auto_master_out_d_bits_data[63:32]; 
  assign data_arrays_1_3_MPORT_2_addr=refill_one_beat ? _mem_idx_T_1:io_req_bits_addr[11:3]; 
  assign data_arrays_1_3_MPORT_2_mask=repl_way_v0==2'h3; 
  assign data_arrays_1_3_MPORT_2_en=refill_one_beat&~invalidated; 
  assign s0_valid=io_req_ready&io_req_valid; 
  assign s1_vb_lo=io_s1_paddr[11:6]; 
  assign _s1_vb_T={1'h0,s1_vb_lo}; 
  assign _s1_vb_T_1=vb_array>>_s1_vb_T; 
  assign s1_vb=_s1_vb_T_1[0]; 
  assign tag=tag_array_0_tag_rdata_data[19:0]; 
  assign s1_tag=io_s1_paddr[31:12]; 
  assign _tagMatch_T=tag==s1_tag; 
  assign tagMatch=s1_vb&_tagMatch_T; 
  assign _s1_vb_T_4={1'h1,s1_vb_lo}; 
  assign _s1_vb_T_5=vb_array>>_s1_vb_T_4; 
  assign s1_vb_1=_s1_vb_T_5[0]; 
  assign tag_1=tag_array_1_tag_rdata_data[19:0]; 
  assign _tagMatch_T_1=tag_1==s1_tag; 
  assign tagMatch_1=s1_vb_1&_tagMatch_T_1; 
  assign _s1_hit_T=tagMatch|tagMatch_1; 
  assign _s1_vb_T_8={2'h2,s1_vb_lo}; 
  assign _s1_vb_T_9=vb_array>>_s1_vb_T_8; 
  assign s1_vb_2=_s1_vb_T_9[0]; 
  assign tag_2=tag_array_2_tag_rdata_data[19:0]; 
  assign _tagMatch_T_2=tag_2==s1_tag; 
  assign tagMatch_2=s1_vb_2&_tagMatch_T_2; 
  assign _s1_hit_T_1=_s1_hit_T|tagMatch_2; 
  assign _s1_vb_T_12={2'h3,s1_vb_lo}; 
  assign _s1_vb_T_13=vb_array>>_s1_vb_T_12; 
  assign s1_vb_3=_s1_vb_T_13[0]; 
  assign tag_3=tag_array_3_tag_rdata_data[19:0]; 
  assign _tagMatch_T_3=tag_3==s1_tag; 
  assign tagMatch_3=s1_vb_3&_tagMatch_T_3; 
  assign _s2_valid_T_1=s1_valid&~io_s1_kill; 
  assign _s2_miss_T_1=s2_valid&~s2_hit; 
  assign s2_miss=_s2_miss_T_1&~io_s2_kill; 
  assign s2_request_refill=s2_miss&s2_request_refill_REG; 
  assign refill_fire=auto_master_out_a_ready&s2_request_refill; 
  assign _s1_can_request_refill_T=s2_miss|refill_valid; 
  assign s1_can_request_refill=~_s1_can_request_refill_T; 
  assign _refill_paddr_T=s1_valid&s1_can_request_refill; 
  assign refill_tag=refill_paddr[31:12]; 
  assign refill_idx=refill_paddr[11:6]; 
  assign refill_one_beat_opdata=auto_master_out_d_bits_opcode[0]; 
  assign refill_one_beat=auto_master_out_d_valid&refill_one_beat_opdata; 
  assign _beats1_decode_T_1=27'hfff<<auto_master_out_d_bits_size; 
  assign beats1_decode=~_beats1_decode_T_1[11:3]; 
  assign beats1=refill_one_beat_opdata ? beats1_decode:9'h0; 
  assign counter1=counter-9'h1; 
  assign first=counter==9'h0; 
  assign _last_T=counter==9'h1; 
  assign _last_T_1=beats1==9'h0; 
  assign last=_last_T|_last_T_1; 
  assign d_done=last&auto_master_out_d_valid; 
  assign refill_cnt=beats1&~counter1; 
  assign refill_done=refill_one_beat&d_done; 
  assign repl_way_v0_lo={repl_way_v0_prng_io_out_7,repl_way_v0_prng_io_out_6,repl_way_v0_prng_io_out_5,repl_way_v0_prng_io_out_4,repl_way_v0_prng_io_out_3,repl_way_v0_prng_io_out_2,repl_way_v0_prng_io_out_1,repl_way_v0_prng_io_out_0}; 
  assign _repl_way_v0_T={repl_way_v0_prng_io_out_15,repl_way_v0_prng_io_out_14,repl_way_v0_prng_io_out_13,repl_way_v0_prng_io_out_12,repl_way_v0_prng_io_out_11,repl_way_v0_prng_io_out_10,repl_way_v0_prng_io_out_9,repl_way_v0_prng_io_out_8,repl_way_v0_lo}; 
  assign repl_way_v0=_repl_way_v0_T[1:0]; 
  assign _repl_way_T={repl_way_v0,refill_idx}; 
  assign _refillError_T=refill_cnt>9'h0; 
  assign _refillError_T_1=_refillError_T&accruedRefillError; 
  assign refillError=auto_master_out_d_bits_corrupt|_refillError_T_1; 
  assign _vb_array_T_2=refill_done&~invalidated; 
  assign _vb_array_T_3=256'h1<<_repl_way_T; 
  assign _vb_array_T_4=vb_array|_vb_array_T_3; 
  assign _vb_array_T_6=~vb_array|_vb_array_T_3; 
  assign s2_tag_disparity=|4'h0; 
  assign _T_40=s2_valid&s2_tag_disparity; 
  assign invalidate=_T_40|io_invalidate; 
  assign _GEN_30=invalidate|invalidated; 
  assign tl_error=tag_array_0_tag_rdata_data[20]; 
  assign s1_tl_error_0=tagMatch&tl_error; 
  assign tl_error_1=tag_array_1_tag_rdata_data[20]; 
  assign s1_tl_error_1=tagMatch_1&tl_error_1; 
  assign tl_error_2=tag_array_2_tag_rdata_data[20]; 
  assign s1_tl_error_2=tagMatch_2&tl_error_2; 
  assign tl_error_3=tag_array_3_tag_rdata_data[20]; 
  assign s1_tl_error_3=tagMatch_3&tl_error_3; 
  assign _T_15=tagMatch+tagMatch_1; 
  assign _T_17=tagMatch_2+tagMatch_3; 
  assign _T_19=_T_15+_T_17; 
  assign _T_21=_T_19<=3'h1; 
  assign _T_22=~s1_valid|_T_21; 
  assign _T_24=_T_22|reset; 
  assign s0_ren=s0_valid&~io_req_bits_addr[2]; 
  assign wen=refill_one_beat&~invalidated; 
  assign _mem_idx_T={refill_idx,3'h0}; 
  assign _mem_idx_T_1=_mem_idx_T|refill_cnt; 
  assign _GEN_54=data_arrays_0_0_dout_data; 
  assign _GEN_55=data_arrays_0_1_dout_data; 
  assign _GEN_56=data_arrays_0_2_dout_data; 
  assign _GEN_57=data_arrays_0_3_dout_data; 
  assign s0_ren_1=s0_valid&io_req_bits_addr[2]; 
  assign _s2_way_mux_T=s2_tag_hit_0 ? s2_dout_0:32'h0; 
  assign _s2_way_mux_T_1=s2_tag_hit_1 ? s2_dout_1:32'h0; 
  assign _s2_way_mux_T_2=s2_tag_hit_2 ? s2_dout_2:32'h0; 
  assign _s2_way_mux_T_3=s2_tag_hit_3 ? s2_dout_3:32'h0; 
  assign _s2_way_mux_T_4=_s2_way_mux_T|_s2_way_mux_T_1; 
  assign _s2_way_mux_T_5=_s2_way_mux_T_4|_s2_way_mux_T_2; 
  assign _s2_tl_error_T={s1_tl_error_3,s1_tl_error_2,s1_tl_error_1,s1_tl_error_0}; 
  assign _s2_tl_error_T_1=|_s2_tl_error_T; 
  assign _GEN_101=refill_fire|refill_valid; 
  assign auto_master_out_a_valid=s2_miss&s2_request_refill_REG; 
  assign auto_master_out_a_bits_address={refill_paddr[31:6],6'h0}; 
  assign io_req_ready=~refill_one_beat; 
  assign io_resp_valid=s2_valid&s2_hit; 
  assign io_resp_bits_data=_s2_way_mux_T_5|_s2_way_mux_T_3; 
  assign io_resp_bits_replay=|4'h0; 
  assign io_resp_bits_ae=s2_tl_error; 
  assign repl_way_v0_prng_clock=clock; 
  assign repl_way_v0_prng_reset=reset; 
  assign repl_way_v0_prng_io_increment=auto_master_out_a_ready&s2_request_refill; 
  assign ICache_cov_read_addr=ICache_state; 
  assign ICache_cov_read_data=ICache_cov[ICache_cov_read_addr]; 
  assign ICache_cov_write_data=1'h1; 
  assign ICache_cov_write_addr=ICache_state; 
  assign ICache_cov_write_mask=1'h1; 
  assign ICache_cov_write_en=1'h1; 
  assign s2_valid_shl=s2_valid; 
  assign s2_valid_pad={5'h0,s2_valid_shl}; 
  assign s1_valid_shl={s1_valid,1'h0}; 
  assign s1_valid_pad={4'h0,s1_valid_shl}; 
  assign refill_valid_shl={refill_valid,2'h0}; 
  assign refill_valid_pad={3'h0,refill_valid_shl}; 
  assign invalidated_shl={invalidated,3'h0}; 
  assign invalidated_pad={2'h0,invalidated_shl}; 
  assign s2_hit_shl={s2_hit,4'h0}; 
  assign s2_hit_pad={1'h0,s2_hit_shl}; 
  assign s2_tag_hit_0_shl={s2_tag_hit_0,5'h0}; 
  assign s2_tag_hit_0_pad=s2_tag_hit_0_shl; 
  assign s2_tag_hit_1_shl={s2_tag_hit_1,5'h0}; 
  assign s2_tag_hit_1_pad=s2_tag_hit_1_shl; 
  assign s2_tag_hit_2_shl={s2_tag_hit_2,5'h0}; 
  assign s2_tag_hit_2_pad=s2_tag_hit_2_shl; 
  assign s2_tag_hit_3_shl={s2_tag_hit_3,5'h0}; 
  assign s2_tag_hit_3_pad=s2_tag_hit_3_shl; 
  assign ICache_xor3=s2_valid_pad^s1_valid_pad; 
  assign ICache_xor4=refill_valid_pad^invalidated_pad; 
  assign ICache_xor1=ICache_xor3^ICache_xor4; 
  assign ICache_xor5=s2_hit_pad^s2_tag_hit_0_pad; 
  assign ICache_xor14=s2_tag_hit_2_pad^s2_tag_hit_3_pad; 
  assign ICache_xor6=s2_tag_hit_1_pad^ICache_xor14; 
  assign ICache_xor2=ICache_xor5^ICache_xor6; 
  assign ICache_xor0=ICache_xor1^ICache_xor2; 
  assign repl_way_v0_prng_sum=ICache_covSum+repl_way_v0_prng_io_covSum; 
  assign io_covSum=repl_way_v0_prng_sum; 
  assign stopEn0=~_T_24; 
  assign repl_way_v0_prng_metaAssert_wire=repl_way_v0_prng_metaAssert; 
  assign ICache_or0=stopEn0|repl_way_v0_prng_metaAssert_wire; 
  assign metaAssert=ICache_metaAssert; 
  assign repl_way_v0_prng_metaReset=metaReset|repl_way_v0_prng_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (tag_array_0_MPORT_en&tag_array_0_MPORT_mask)
            begin 
              tag_array_0 [tag_array_0_MPORT_addr]<=tag_array_0_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_0_tag_rdata_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_0_tag_rdata_en_pipe_0 <=~refill_done&s0_valid;
            end 
         if (metaReset)
            begin 
              tag_array_0_tag_rdata_addr_pipe_0 <=6'h0;
            end 
          else 
            if (~refill_done&s0_valid)
               begin 
                 tag_array_0_tag_rdata_addr_pipe_0 <=io_req_bits_addr[11:6];
               end 
         if (tag_array_1_MPORT_en&tag_array_1_MPORT_mask)
            begin 
              tag_array_1 [tag_array_1_MPORT_addr]<=tag_array_1_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_1_tag_rdata_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_1_tag_rdata_en_pipe_0 <=~refill_done&s0_valid;
            end 
         if (metaReset)
            begin 
              tag_array_1_tag_rdata_addr_pipe_0 <=6'h0;
            end 
          else 
            if (~refill_done&s0_valid)
               begin 
                 tag_array_1_tag_rdata_addr_pipe_0 <=io_req_bits_addr[11:6];
               end 
         if (tag_array_2_MPORT_en&tag_array_2_MPORT_mask)
            begin 
              tag_array_2 [tag_array_2_MPORT_addr]<=tag_array_2_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_2_tag_rdata_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_2_tag_rdata_en_pipe_0 <=~refill_done&s0_valid;
            end 
         if (metaReset)
            begin 
              tag_array_2_tag_rdata_addr_pipe_0 <=6'h0;
            end 
          else 
            if (~refill_done&s0_valid)
               begin 
                 tag_array_2_tag_rdata_addr_pipe_0 <=io_req_bits_addr[11:6];
               end 
         if (tag_array_3_MPORT_en&tag_array_3_MPORT_mask)
            begin 
              tag_array_3 [tag_array_3_MPORT_addr]<=tag_array_3_MPORT_data;
            end 
         if (metaReset)
            begin 
              tag_array_3_tag_rdata_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              tag_array_3_tag_rdata_en_pipe_0 <=~refill_done&s0_valid;
            end 
         if (metaReset)
            begin 
              tag_array_3_tag_rdata_addr_pipe_0 <=6'h0;
            end 
          else 
            if (~refill_done&s0_valid)
               begin 
                 tag_array_3_tag_rdata_addr_pipe_0 <=io_req_bits_addr[11:6];
               end 
         if (data_arrays_0_0_MPORT_1_en&data_arrays_0_0_MPORT_1_mask)
            begin 
              data_arrays_0_0 [data_arrays_0_0_MPORT_1_addr]<=data_arrays_0_0_MPORT_1_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_0_dout_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_0_dout_en_pipe_0 <=~wen&s0_ren;
            end 
         if (metaReset)
            begin 
              data_arrays_0_0_dout_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_0_0_dout_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_0_0_dout_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (data_arrays_0_1_MPORT_1_en&data_arrays_0_1_MPORT_1_mask)
            begin 
              data_arrays_0_1 [data_arrays_0_1_MPORT_1_addr]<=data_arrays_0_1_MPORT_1_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_1_dout_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_1_dout_en_pipe_0 <=~wen&s0_ren;
            end 
         if (metaReset)
            begin 
              data_arrays_0_1_dout_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_0_1_dout_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_0_1_dout_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (data_arrays_0_2_MPORT_1_en&data_arrays_0_2_MPORT_1_mask)
            begin 
              data_arrays_0_2 [data_arrays_0_2_MPORT_1_addr]<=data_arrays_0_2_MPORT_1_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_2_dout_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_2_dout_en_pipe_0 <=~wen&s0_ren;
            end 
         if (metaReset)
            begin 
              data_arrays_0_2_dout_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_0_2_dout_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_0_2_dout_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (data_arrays_0_3_MPORT_1_en&data_arrays_0_3_MPORT_1_mask)
            begin 
              data_arrays_0_3 [data_arrays_0_3_MPORT_1_addr]<=data_arrays_0_3_MPORT_1_data;
            end 
         if (metaReset)
            begin 
              data_arrays_0_3_dout_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_0_3_dout_en_pipe_0 <=~wen&s0_ren;
            end 
         if (metaReset)
            begin 
              data_arrays_0_3_dout_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_0_3_dout_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_0_3_dout_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (data_arrays_1_0_MPORT_2_en&data_arrays_1_0_MPORT_2_mask)
            begin 
              data_arrays_1_0 [data_arrays_1_0_MPORT_2_addr]<=data_arrays_1_0_MPORT_2_data;
            end 
         if (metaReset)
            begin 
              data_arrays_1_0_dout_1_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_1_0_dout_1_en_pipe_0 <=~wen&s0_ren_1;
            end 
         if (metaReset)
            begin 
              data_arrays_1_0_dout_1_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren_1)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_1_0_dout_1_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_1_0_dout_1_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (data_arrays_1_1_MPORT_2_en&data_arrays_1_1_MPORT_2_mask)
            begin 
              data_arrays_1_1 [data_arrays_1_1_MPORT_2_addr]<=data_arrays_1_1_MPORT_2_data;
            end 
         if (metaReset)
            begin 
              data_arrays_1_1_dout_1_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_1_1_dout_1_en_pipe_0 <=~wen&s0_ren_1;
            end 
         if (metaReset)
            begin 
              data_arrays_1_1_dout_1_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren_1)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_1_1_dout_1_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_1_1_dout_1_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (data_arrays_1_2_MPORT_2_en&data_arrays_1_2_MPORT_2_mask)
            begin 
              data_arrays_1_2 [data_arrays_1_2_MPORT_2_addr]<=data_arrays_1_2_MPORT_2_data;
            end 
         if (metaReset)
            begin 
              data_arrays_1_2_dout_1_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_1_2_dout_1_en_pipe_0 <=~wen&s0_ren_1;
            end 
         if (metaReset)
            begin 
              data_arrays_1_2_dout_1_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren_1)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_1_2_dout_1_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_1_2_dout_1_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (data_arrays_1_3_MPORT_2_en&data_arrays_1_3_MPORT_2_mask)
            begin 
              data_arrays_1_3 [data_arrays_1_3_MPORT_2_addr]<=data_arrays_1_3_MPORT_2_data;
            end 
         if (metaReset)
            begin 
              data_arrays_1_3_dout_1_en_pipe_0 <=1'h0;
            end 
          else 
            begin 
              data_arrays_1_3_dout_1_en_pipe_0 <=~wen&s0_ren_1;
            end 
         if (metaReset)
            begin 
              data_arrays_1_3_dout_1_addr_pipe_0 <=9'h0;
            end 
          else 
            if (~wen&s0_ren_1)
               begin 
                 if (refill_one_beat)
                    begin 
                      data_arrays_1_3_dout_1_addr_pipe_0 <=_mem_idx_T_1;
                    end 
                  else 
                    begin 
                      data_arrays_1_3_dout_1_addr_pipe_0 <=io_req_bits_addr[11:3];
                    end 
               end 
         if (metaReset)
            begin 
              s1_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s1_valid <=1'h0;
               end 
             else 
               begin 
                 s1_valid <=s0_valid;
               end 
         if (metaReset)
            begin 
              vb_array <=256'h0;
            end 
          else 
            if (reset)
               begin 
                 vb_array <=256'h0;
               end 
             else 
               if (invalidate)
                  begin 
                    vb_array <=256'h0;
                  end 
                else 
                  if (refill_one_beat)
                     begin 
                       if (_vb_array_T_2)
                          begin 
                            vb_array <=_vb_array_T_4;
                          end 
                        else 
                          begin 
                            vb_array <=~_vb_array_T_6;
                          end 
                     end 
         if (metaReset)
            begin 
              s2_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 s2_valid <=1'h0;
               end 
             else 
               begin 
                 s2_valid <=_s2_valid_T_1;
               end 
         if (metaReset)
            begin 
              s2_hit <=1'h0;
            end 
          else 
            begin 
              s2_hit <=_s1_hit_T_1|tagMatch_3;
            end 
         if (metaReset)
            begin 
              invalidated <=1'h0;
            end 
          else 
            if (~refill_valid)
               begin 
                 invalidated <=1'h0;
               end 
             else 
               begin 
                 invalidated <=_GEN_30;
               end 
         if (metaReset)
            begin 
              refill_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 refill_valid <=1'h0;
               end 
             else 
               if (refill_done)
                  begin 
                    refill_valid <=1'h0;
                  end 
                else 
                  begin 
                    refill_valid <=_GEN_101;
                  end 
         if (metaReset)
            begin 
              s2_request_refill_REG <=1'h0;
            end 
          else 
            begin 
              s2_request_refill_REG <=~_s1_can_request_refill_T;
            end 
         if (metaReset)
            begin 
              refill_paddr <=32'h0;
            end 
          else 
            if (_refill_paddr_T)
               begin 
                 refill_paddr <=io_s1_paddr;
               end 
         if (metaReset)
            begin 
              counter <=9'h0;
            end 
          else 
            if (reset)
               begin 
                 counter <=9'h0;
               end 
             else 
               if (auto_master_out_d_valid)
                  begin 
                    if (first)
                       begin 
                         if (refill_one_beat_opdata)
                            begin 
                              counter <=beats1_decode;
                            end 
                          else 
                            begin 
                              counter <=9'h0;
                            end 
                       end 
                     else 
                       begin 
                         counter <=counter1;
                       end 
                  end 
         if (metaReset)
            begin 
              accruedRefillError <=1'h0;
            end 
          else 
            if (refill_one_beat)
               begin 
                 accruedRefillError <=refillError;
               end 
         if (metaReset)
            begin 
              s2_tag_hit_0 <=1'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 s2_tag_hit_0 <=tagMatch;
               end 
         if (metaReset)
            begin 
              s2_tag_hit_1 <=1'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 s2_tag_hit_1 <=tagMatch_1;
               end 
         if (metaReset)
            begin 
              s2_tag_hit_2 <=1'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 s2_tag_hit_2 <=tagMatch_2;
               end 
         if (metaReset)
            begin 
              s2_tag_hit_3 <=1'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 s2_tag_hit_3 <=tagMatch_3;
               end 
         if (metaReset)
            begin 
              s2_dout_0 <=32'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 if (io_s1_paddr[2])
                    begin 
                      s2_dout_0 <=data_arrays_1_0_dout_1_data;
                    end 
                  else 
                    begin 
                      s2_dout_0 <=_GEN_54;
                    end 
               end 
         if (metaReset)
            begin 
              s2_dout_1 <=32'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 if (io_s1_paddr[2])
                    begin 
                      s2_dout_1 <=data_arrays_1_1_dout_1_data;
                    end 
                  else 
                    begin 
                      s2_dout_1 <=_GEN_55;
                    end 
               end 
         if (metaReset)
            begin 
              s2_dout_2 <=32'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 if (io_s1_paddr[2])
                    begin 
                      s2_dout_2 <=data_arrays_1_2_dout_1_data;
                    end 
                  else 
                    begin 
                      s2_dout_2 <=_GEN_56;
                    end 
               end 
         if (metaReset)
            begin 
              s2_dout_3 <=32'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 if (io_s1_paddr[2])
                    begin 
                      s2_dout_3 <=data_arrays_1_3_dout_1_data;
                    end 
                  else 
                    begin 
                      s2_dout_3 <=_GEN_57;
                    end 
               end 
         if (metaReset)
            begin 
              s2_tl_error <=1'h0;
            end 
          else 
            if (s1_valid)
               begin 
                 s2_tl_error <=_s2_tl_error_T_1;
               end 
         if (~_T_24)
            begin $display("Assertion failed\n    at ICache.scala:267 assert(!(s1_valid || s1_slaveValid) || PopCount(s1_tag_hit zip s1_tag_disparity map { case (h, d) => h && !d }) <= 1)\n");
            end 
         if (~_T_24)
            begin $display("fatal");
            end 
         ICache_state <=ICache_xor0;
         if (!(ICache_cov_read_data))
            begin 
              ICache_covSum <=ICache_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              ICache_metaAssert <=1'h0;
            end 
          else 
            begin 
              ICache_metaAssert <=ICache_metaAssert|ICache_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (ICache_cov_write_en&ICache_cov_write_mask)
            begin 
              ICache_cov [ICache_cov_write_addr]<=ICache_cov_write_data;
            end 
       end
  
endmodule
 
module ShiftQueue (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input io_enq_bits_btb_taken,
  input io_enq_bits_btb_bridx,
  input [4:0] io_enq_bits_btb_entry,
  input [7:0] io_enq_bits_btb_bht_history,
  input [39:0] io_enq_bits_pc,
  input [31:0] io_enq_bits_data,
  input [1:0] io_enq_bits_mask,
  input io_enq_bits_xcpt_pf_inst,
  input io_enq_bits_xcpt_ae_inst,
  input io_enq_bits_replay,
  input io_deq_ready,
  output io_deq_valid,
  output io_deq_bits_btb_taken,
  output io_deq_bits_btb_bridx,
  output [4:0] io_deq_bits_btb_entry,
  output [7:0] io_deq_bits_btb_bht_history,
  output [39:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_data,
  output io_deq_bits_xcpt_pf_inst,
  output io_deq_bits_xcpt_ae_inst,
  output io_deq_bits_replay,
  output [4:0] io_mask,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg valid_0 ;  
   reg [31:0] _RAND_0 ;  
   reg valid_1 ;  
   reg [31:0] _RAND_1 ;  
   reg valid_2 ;  
   reg [31:0] _RAND_2 ;  
   reg valid_3 ;  
   reg [31:0] _RAND_3 ;  
   reg valid_4 ;  
   reg [31:0] _RAND_4 ;  
   reg elts_0_btb_taken ;  
   reg [31:0] _RAND_5 ;  
   reg elts_0_btb_bridx ;  
   reg [31:0] _RAND_6 ;  
   reg [4:0] elts_0_btb_entry ;  
   reg [31:0] _RAND_7 ;  
   reg [7:0] elts_0_btb_bht_history ;  
   reg [31:0] _RAND_8 ;  
   reg [39:0] elts_0_pc ;  
   reg [63:0] _RAND_9 ;  
   reg [31:0] elts_0_data ;  
   reg [31:0] _RAND_10 ;  
   reg elts_0_xcpt_pf_inst ;  
   reg [31:0] _RAND_11 ;  
   reg elts_0_xcpt_ae_inst ;  
   reg [31:0] _RAND_12 ;  
   reg elts_0_replay ;  
   reg [31:0] _RAND_13 ;  
   reg elts_1_btb_taken ;  
   reg [31:0] _RAND_14 ;  
   reg elts_1_btb_bridx ;  
   reg [31:0] _RAND_15 ;  
   reg [4:0] elts_1_btb_entry ;  
   reg [31:0] _RAND_16 ;  
   reg [7:0] elts_1_btb_bht_history ;  
   reg [31:0] _RAND_17 ;  
   reg [39:0] elts_1_pc ;  
   reg [63:0] _RAND_18 ;  
   reg [31:0] elts_1_data ;  
   reg [31:0] _RAND_19 ;  
   reg elts_1_xcpt_pf_inst ;  
   reg [31:0] _RAND_20 ;  
   reg elts_1_xcpt_ae_inst ;  
   reg [31:0] _RAND_21 ;  
   reg elts_1_replay ;  
   reg [31:0] _RAND_22 ;  
   reg elts_2_btb_taken ;  
   reg [31:0] _RAND_23 ;  
   reg elts_2_btb_bridx ;  
   reg [31:0] _RAND_24 ;  
   reg [4:0] elts_2_btb_entry ;  
   reg [31:0] _RAND_25 ;  
   reg [7:0] elts_2_btb_bht_history ;  
   reg [31:0] _RAND_26 ;  
   reg [39:0] elts_2_pc ;  
   reg [63:0] _RAND_27 ;  
   reg [31:0] elts_2_data ;  
   reg [31:0] _RAND_28 ;  
   reg elts_2_xcpt_pf_inst ;  
   reg [31:0] _RAND_29 ;  
   reg elts_2_xcpt_ae_inst ;  
   reg [31:0] _RAND_30 ;  
   reg elts_2_replay ;  
   reg [31:0] _RAND_31 ;  
   reg elts_3_btb_taken ;  
   reg [31:0] _RAND_32 ;  
   reg elts_3_btb_bridx ;  
   reg [31:0] _RAND_33 ;  
   reg [4:0] elts_3_btb_entry ;  
   reg [31:0] _RAND_34 ;  
   reg [7:0] elts_3_btb_bht_history ;  
   reg [31:0] _RAND_35 ;  
   reg [39:0] elts_3_pc ;  
   reg [63:0] _RAND_36 ;  
   reg [31:0] elts_3_data ;  
   reg [31:0] _RAND_37 ;  
   reg elts_3_xcpt_pf_inst ;  
   reg [31:0] _RAND_38 ;  
   reg elts_3_xcpt_ae_inst ;  
   reg [31:0] _RAND_39 ;  
   reg elts_3_replay ;  
   reg [31:0] _RAND_40 ;  
   reg elts_4_btb_taken ;  
   reg [31:0] _RAND_41 ;  
   reg elts_4_btb_bridx ;  
   reg [31:0] _RAND_42 ;  
   reg [4:0] elts_4_btb_entry ;  
   reg [31:0] _RAND_43 ;  
   reg [7:0] elts_4_btb_bht_history ;  
   reg [31:0] _RAND_44 ;  
   reg [39:0] elts_4_pc ;  
   reg [63:0] _RAND_45 ;  
   reg [31:0] elts_4_data ;  
   reg [31:0] _RAND_46 ;  
   reg elts_4_xcpt_pf_inst ;  
   reg [31:0] _RAND_47 ;  
   reg elts_4_xcpt_ae_inst ;  
   reg [31:0] _RAND_48 ;  
   reg elts_4_replay ;  
   reg [31:0] _RAND_49 ;  
   wire _wen_T ;  
   wire _wen_T_2 ;  
   wire _wen_T_3 ;  
   wire _wen_T_7 ;  
   wire wen ;  
   wire _valid_0_T_6 ;  
   wire _wen_T_10 ;  
   wire _wen_T_11 ;  
   wire _wen_T_15 ;  
   wire wen_1 ;  
   wire _valid_1_T_6 ;  
   wire _wen_T_18 ;  
   wire _wen_T_19 ;  
   wire _wen_T_23 ;  
   wire wen_2 ;  
   wire _valid_2_T_6 ;  
   wire _wen_T_26 ;  
   wire _wen_T_27 ;  
   wire _wen_T_31 ;  
   wire wen_3 ;  
   wire _valid_3_T_6 ;  
   wire _wen_T_34 ;  
   wire _wen_T_39 ;  
   wire wen_4 ;  
   wire _valid_4_T_6 ;  
   wire [1:0] io_mask_lo ;  
   wire [2:0] io_mask_hi ;  
   reg ShiftQueue_state ;  
   reg [31:0] _RAND_50 ;  
   reg ShiftQueue_cov[0:1] ;  
   reg [31:0] _RAND_51 ;  
   wire ShiftQueue_cov_read_data ;  
   wire ShiftQueue_cov_read_addr ;  
   wire ShiftQueue_cov_write_data ;  
   wire ShiftQueue_cov_write_addr ;  
   wire ShiftQueue_cov_write_mask ;  
   wire ShiftQueue_cov_write_en ;  
   reg [29:0] ShiftQueue_covSum ;  
   reg [31:0] _RAND_52 ;  
   wire valid_1_shl ;  
   wire valid_1_pad ;  
   wire valid_0_shl ;  
   wire valid_0_pad ;  
   wire valid_2_shl ;  
   wire valid_2_pad ;  
   wire valid_4_shl ;  
   wire valid_4_pad ;  
   wire valid_3_shl ;  
   wire valid_3_pad ;  
   wire ShiftQueue_xor1 ;  
   wire ShiftQueue_xor6 ;  
   wire ShiftQueue_xor2 ;  
   wire ShiftQueue_xor0 ;  
  assign _wen_T=io_enq_ready&io_enq_valid; 
  assign _wen_T_2=_wen_T&valid_0; 
  assign _wen_T_3=valid_1|_wen_T_2; 
  assign _wen_T_7=_wen_T&~valid_0; 
  assign wen=io_deq_ready ? _wen_T_3:_wen_T_7; 
  assign _valid_0_T_6=_wen_T|valid_0; 
  assign _wen_T_10=_wen_T&valid_1; 
  assign _wen_T_11=valid_2|_wen_T_10; 
  assign _wen_T_15=_wen_T_2&~valid_1; 
  assign wen_1=io_deq_ready ? _wen_T_11:_wen_T_15; 
  assign _valid_1_T_6=_wen_T_2|valid_1; 
  assign _wen_T_18=_wen_T&valid_2; 
  assign _wen_T_19=valid_3|_wen_T_18; 
  assign _wen_T_23=_wen_T_10&~valid_2; 
  assign wen_2=io_deq_ready ? _wen_T_19:_wen_T_23; 
  assign _valid_2_T_6=_wen_T_10|valid_2; 
  assign _wen_T_26=_wen_T&valid_3; 
  assign _wen_T_27=valid_4|_wen_T_26; 
  assign _wen_T_31=_wen_T_18&~valid_3; 
  assign wen_3=io_deq_ready ? _wen_T_27:_wen_T_31; 
  assign _valid_3_T_6=_wen_T_18|valid_3; 
  assign _wen_T_34=_wen_T&valid_4; 
  assign _wen_T_39=_wen_T_26&~valid_4; 
  assign wen_4=io_deq_ready ? _wen_T_34:_wen_T_39; 
  assign _valid_4_T_6=_wen_T_26|valid_4; 
  assign io_mask_lo={valid_1,valid_0}; 
  assign io_mask_hi={valid_4,valid_3,valid_2}; 
  assign io_enq_ready=~valid_4; 
  assign io_deq_valid=io_enq_valid|valid_0; 
  assign io_deq_bits_btb_taken=valid_0 ? elts_0_btb_taken:io_enq_bits_btb_taken; 
  assign io_deq_bits_btb_bridx=valid_0 ? elts_0_btb_bridx:io_enq_bits_btb_bridx; 
  assign io_deq_bits_btb_entry=valid_0 ? elts_0_btb_entry:io_enq_bits_btb_entry; 
  assign io_deq_bits_btb_bht_history=valid_0 ? elts_0_btb_bht_history:io_enq_bits_btb_bht_history; 
  assign io_deq_bits_pc=valid_0 ? elts_0_pc:io_enq_bits_pc; 
  assign io_deq_bits_data=valid_0 ? elts_0_data:io_enq_bits_data; 
  assign io_deq_bits_xcpt_pf_inst=valid_0 ? elts_0_xcpt_pf_inst:io_enq_bits_xcpt_pf_inst; 
  assign io_deq_bits_xcpt_ae_inst=valid_0 ? elts_0_xcpt_ae_inst:io_enq_bits_xcpt_ae_inst; 
  assign io_deq_bits_replay=valid_0 ? elts_0_replay:io_enq_bits_replay; 
  assign io_mask={io_mask_hi,io_mask_lo}; 
  assign ShiftQueue_cov_read_addr=ShiftQueue_state; 
  assign ShiftQueue_cov_read_data=ShiftQueue_cov[ShiftQueue_cov_read_addr]; 
  assign ShiftQueue_cov_write_data=1'h1; 
  assign ShiftQueue_cov_write_addr=ShiftQueue_state; 
  assign ShiftQueue_cov_write_mask=1'h1; 
  assign ShiftQueue_cov_write_en=1'h1; 
  assign valid_1_shl=valid_1; 
  assign valid_1_pad=valid_1_shl; 
  assign valid_0_shl=valid_0; 
  assign valid_0_pad=valid_0_shl; 
  assign valid_2_shl=valid_2; 
  assign valid_2_pad=valid_2_shl; 
  assign valid_4_shl=valid_4; 
  assign valid_4_pad=valid_4_shl; 
  assign valid_3_shl=valid_3; 
  assign valid_3_pad=valid_3_shl; 
  assign ShiftQueue_xor1=valid_1_pad^valid_0_pad; 
  assign ShiftQueue_xor6=valid_4_pad^valid_3_pad; 
  assign ShiftQueue_xor2=valid_2_pad^ShiftQueue_xor6; 
  assign ShiftQueue_xor0=ShiftQueue_xor1^ShiftQueue_xor2; 
  assign io_covSum=ShiftQueue_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              valid_0 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 valid_0 <=1'h0;
               end 
             else 
               if (io_deq_ready)
                  begin 
                    valid_0 <=_wen_T_3;
                  end 
                else 
                  begin 
                    valid_0 <=_valid_0_T_6;
                  end 
         if (metaReset)
            begin 
              valid_1 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 valid_1 <=1'h0;
               end 
             else 
               if (io_deq_ready)
                  begin 
                    valid_1 <=_wen_T_11;
                  end 
                else 
                  begin 
                    valid_1 <=_valid_1_T_6;
                  end 
         if (metaReset)
            begin 
              valid_2 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 valid_2 <=1'h0;
               end 
             else 
               if (io_deq_ready)
                  begin 
                    valid_2 <=_wen_T_19;
                  end 
                else 
                  begin 
                    valid_2 <=_valid_2_T_6;
                  end 
         if (metaReset)
            begin 
              valid_3 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 valid_3 <=1'h0;
               end 
             else 
               if (io_deq_ready)
                  begin 
                    valid_3 <=_wen_T_27;
                  end 
                else 
                  begin 
                    valid_3 <=_valid_3_T_6;
                  end 
         if (metaReset)
            begin 
              valid_4 <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 valid_4 <=1'h0;
               end 
             else 
               if (io_deq_ready)
                  begin 
                    valid_4 <=_wen_T_34;
                  end 
                else 
                  begin 
                    valid_4 <=_valid_4_T_6;
                  end 
         if (metaReset)
            begin 
              elts_0_btb_taken <=1'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_btb_taken <=elts_1_btb_taken;
                    end 
                  else 
                    begin 
                      elts_0_btb_taken <=io_enq_bits_btb_taken;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_btb_bridx <=1'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_btb_bridx <=elts_1_btb_bridx;
                    end 
                  else 
                    begin 
                      elts_0_btb_bridx <=io_enq_bits_btb_bridx;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_btb_entry <=5'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_btb_entry <=elts_1_btb_entry;
                    end 
                  else 
                    begin 
                      elts_0_btb_entry <=io_enq_bits_btb_entry;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_btb_bht_history <=8'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_btb_bht_history <=elts_1_btb_bht_history;
                    end 
                  else 
                    begin 
                      elts_0_btb_bht_history <=io_enq_bits_btb_bht_history;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_pc <=40'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_pc <=elts_1_pc;
                    end 
                  else 
                    begin 
                      elts_0_pc <=io_enq_bits_pc;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_data <=32'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_data <=elts_1_data;
                    end 
                  else 
                    begin 
                      elts_0_data <=io_enq_bits_data;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_xcpt_pf_inst <=1'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_xcpt_pf_inst <=elts_1_xcpt_pf_inst;
                    end 
                  else 
                    begin 
                      elts_0_xcpt_pf_inst <=io_enq_bits_xcpt_pf_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_xcpt_ae_inst <=1'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_xcpt_ae_inst <=elts_1_xcpt_ae_inst;
                    end 
                  else 
                    begin 
                      elts_0_xcpt_ae_inst <=io_enq_bits_xcpt_ae_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_0_replay <=1'h0;
            end 
          else 
            if (wen)
               begin 
                 if (valid_1)
                    begin 
                      elts_0_replay <=elts_1_replay;
                    end 
                  else 
                    begin 
                      elts_0_replay <=io_enq_bits_replay;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_btb_taken <=1'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_btb_taken <=elts_2_btb_taken;
                    end 
                  else 
                    begin 
                      elts_1_btb_taken <=io_enq_bits_btb_taken;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_btb_bridx <=1'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_btb_bridx <=elts_2_btb_bridx;
                    end 
                  else 
                    begin 
                      elts_1_btb_bridx <=io_enq_bits_btb_bridx;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_btb_entry <=5'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_btb_entry <=elts_2_btb_entry;
                    end 
                  else 
                    begin 
                      elts_1_btb_entry <=io_enq_bits_btb_entry;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_btb_bht_history <=8'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_btb_bht_history <=elts_2_btb_bht_history;
                    end 
                  else 
                    begin 
                      elts_1_btb_bht_history <=io_enq_bits_btb_bht_history;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_pc <=40'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_pc <=elts_2_pc;
                    end 
                  else 
                    begin 
                      elts_1_pc <=io_enq_bits_pc;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_data <=32'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_data <=elts_2_data;
                    end 
                  else 
                    begin 
                      elts_1_data <=io_enq_bits_data;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_xcpt_pf_inst <=1'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_xcpt_pf_inst <=elts_2_xcpt_pf_inst;
                    end 
                  else 
                    begin 
                      elts_1_xcpt_pf_inst <=io_enq_bits_xcpt_pf_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_xcpt_ae_inst <=1'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_xcpt_ae_inst <=elts_2_xcpt_ae_inst;
                    end 
                  else 
                    begin 
                      elts_1_xcpt_ae_inst <=io_enq_bits_xcpt_ae_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_1_replay <=1'h0;
            end 
          else 
            if (wen_1)
               begin 
                 if (valid_2)
                    begin 
                      elts_1_replay <=elts_2_replay;
                    end 
                  else 
                    begin 
                      elts_1_replay <=io_enq_bits_replay;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_btb_taken <=1'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_btb_taken <=elts_3_btb_taken;
                    end 
                  else 
                    begin 
                      elts_2_btb_taken <=io_enq_bits_btb_taken;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_btb_bridx <=1'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_btb_bridx <=elts_3_btb_bridx;
                    end 
                  else 
                    begin 
                      elts_2_btb_bridx <=io_enq_bits_btb_bridx;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_btb_entry <=5'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_btb_entry <=elts_3_btb_entry;
                    end 
                  else 
                    begin 
                      elts_2_btb_entry <=io_enq_bits_btb_entry;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_btb_bht_history <=8'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_btb_bht_history <=elts_3_btb_bht_history;
                    end 
                  else 
                    begin 
                      elts_2_btb_bht_history <=io_enq_bits_btb_bht_history;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_pc <=40'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_pc <=elts_3_pc;
                    end 
                  else 
                    begin 
                      elts_2_pc <=io_enq_bits_pc;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_data <=32'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_data <=elts_3_data;
                    end 
                  else 
                    begin 
                      elts_2_data <=io_enq_bits_data;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_xcpt_pf_inst <=1'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_xcpt_pf_inst <=elts_3_xcpt_pf_inst;
                    end 
                  else 
                    begin 
                      elts_2_xcpt_pf_inst <=io_enq_bits_xcpt_pf_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_xcpt_ae_inst <=1'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_xcpt_ae_inst <=elts_3_xcpt_ae_inst;
                    end 
                  else 
                    begin 
                      elts_2_xcpt_ae_inst <=io_enq_bits_xcpt_ae_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_2_replay <=1'h0;
            end 
          else 
            if (wen_2)
               begin 
                 if (valid_3)
                    begin 
                      elts_2_replay <=elts_3_replay;
                    end 
                  else 
                    begin 
                      elts_2_replay <=io_enq_bits_replay;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_btb_taken <=1'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_btb_taken <=elts_4_btb_taken;
                    end 
                  else 
                    begin 
                      elts_3_btb_taken <=io_enq_bits_btb_taken;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_btb_bridx <=1'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_btb_bridx <=elts_4_btb_bridx;
                    end 
                  else 
                    begin 
                      elts_3_btb_bridx <=io_enq_bits_btb_bridx;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_btb_entry <=5'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_btb_entry <=elts_4_btb_entry;
                    end 
                  else 
                    begin 
                      elts_3_btb_entry <=io_enq_bits_btb_entry;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_btb_bht_history <=8'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_btb_bht_history <=elts_4_btb_bht_history;
                    end 
                  else 
                    begin 
                      elts_3_btb_bht_history <=io_enq_bits_btb_bht_history;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_pc <=40'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_pc <=elts_4_pc;
                    end 
                  else 
                    begin 
                      elts_3_pc <=io_enq_bits_pc;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_data <=32'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_data <=elts_4_data;
                    end 
                  else 
                    begin 
                      elts_3_data <=io_enq_bits_data;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_xcpt_pf_inst <=1'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_xcpt_pf_inst <=elts_4_xcpt_pf_inst;
                    end 
                  else 
                    begin 
                      elts_3_xcpt_pf_inst <=io_enq_bits_xcpt_pf_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_xcpt_ae_inst <=1'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_xcpt_ae_inst <=elts_4_xcpt_ae_inst;
                    end 
                  else 
                    begin 
                      elts_3_xcpt_ae_inst <=io_enq_bits_xcpt_ae_inst;
                    end 
               end 
         if (metaReset)
            begin 
              elts_3_replay <=1'h0;
            end 
          else 
            if (wen_3)
               begin 
                 if (valid_4)
                    begin 
                      elts_3_replay <=elts_4_replay;
                    end 
                  else 
                    begin 
                      elts_3_replay <=io_enq_bits_replay;
                    end 
               end 
         if (metaReset)
            begin 
              elts_4_btb_taken <=1'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_btb_taken <=io_enq_bits_btb_taken;
               end 
         if (metaReset)
            begin 
              elts_4_btb_bridx <=1'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_btb_bridx <=io_enq_bits_btb_bridx;
               end 
         if (metaReset)
            begin 
              elts_4_btb_entry <=5'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_btb_entry <=io_enq_bits_btb_entry;
               end 
         if (metaReset)
            begin 
              elts_4_btb_bht_history <=8'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_btb_bht_history <=io_enq_bits_btb_bht_history;
               end 
         if (metaReset)
            begin 
              elts_4_pc <=40'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_pc <=io_enq_bits_pc;
               end 
         if (metaReset)
            begin 
              elts_4_data <=32'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_data <=io_enq_bits_data;
               end 
         if (metaReset)
            begin 
              elts_4_xcpt_pf_inst <=1'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_xcpt_pf_inst <=io_enq_bits_xcpt_pf_inst;
               end 
         if (metaReset)
            begin 
              elts_4_xcpt_ae_inst <=1'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_xcpt_ae_inst <=io_enq_bits_xcpt_ae_inst;
               end 
         if (metaReset)
            begin 
              elts_4_replay <=1'h0;
            end 
          else 
            if (wen_4)
               begin 
                 elts_4_replay <=io_enq_bits_replay;
               end 
         ShiftQueue_state <=ShiftQueue_xor0;
         if (!(ShiftQueue_cov_read_data))
            begin 
              ShiftQueue_covSum <=ShiftQueue_covSum+1'h1;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (ShiftQueue_cov_write_en&ShiftQueue_cov_write_mask)
            begin 
              ShiftQueue_cov [ShiftQueue_cov_write_addr]<=ShiftQueue_cov_write_data;
            end 
       end
  
endmodule
 
module TLB_1 (
  input clock,
  input reset,
  output io_req_ready,
  input io_req_valid,
  input [39:0] io_req_bits_vaddr,
  output io_resp_miss,
  output [31:0] io_resp_paddr,
  output io_resp_pf_inst,
  output io_resp_ae_inst,
  output io_resp_cacheable,
  input io_sfence_valid,
  input io_sfence_bits_rs1,
  input io_sfence_bits_rs2,
  input [38:0] io_sfence_bits_addr,
  input io_ptw_req_ready,
  output io_ptw_req_valid,
  output io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  input io_ptw_resp_valid,
  input io_ptw_resp_bits_ae,
  input [53:0] io_ptw_resp_bits_pte_ppn,
  input io_ptw_resp_bits_pte_d,
  input io_ptw_resp_bits_pte_a,
  input io_ptw_resp_bits_pte_g,
  input io_ptw_resp_bits_pte_u,
  input io_ptw_resp_bits_pte_x,
  input io_ptw_resp_bits_pte_w,
  input io_ptw_resp_bits_pte_r,
  input io_ptw_resp_bits_pte_v,
  input [1:0] io_ptw_resp_bits_level,
  input io_ptw_resp_bits_homogeneous,
  input [3:0] io_ptw_ptbr_mode,
  input io_ptw_status_debug,
  input [1:0] io_ptw_status_prv,
  input io_ptw_pmp_0_cfg_l,
  input [1:0] io_ptw_pmp_0_cfg_a,
  input io_ptw_pmp_0_cfg_x,
  input io_ptw_pmp_0_cfg_w,
  input io_ptw_pmp_0_cfg_r,
  input [29:0] io_ptw_pmp_0_addr,
  input [31:0] io_ptw_pmp_0_mask,
  input io_ptw_pmp_1_cfg_l,
  input [1:0] io_ptw_pmp_1_cfg_a,
  input io_ptw_pmp_1_cfg_x,
  input io_ptw_pmp_1_cfg_w,
  input io_ptw_pmp_1_cfg_r,
  input [29:0] io_ptw_pmp_1_addr,
  input [31:0] io_ptw_pmp_1_mask,
  input io_ptw_pmp_2_cfg_l,
  input [1:0] io_ptw_pmp_2_cfg_a,
  input io_ptw_pmp_2_cfg_x,
  input io_ptw_pmp_2_cfg_w,
  input io_ptw_pmp_2_cfg_r,
  input [29:0] io_ptw_pmp_2_addr,
  input [31:0] io_ptw_pmp_2_mask,
  input io_ptw_pmp_3_cfg_l,
  input [1:0] io_ptw_pmp_3_cfg_a,
  input io_ptw_pmp_3_cfg_x,
  input io_ptw_pmp_3_cfg_w,
  input io_ptw_pmp_3_cfg_r,
  input [29:0] io_ptw_pmp_3_addr,
  input [31:0] io_ptw_pmp_3_mask,
  input io_ptw_pmp_4_cfg_l,
  input [1:0] io_ptw_pmp_4_cfg_a,
  input io_ptw_pmp_4_cfg_x,
  input io_ptw_pmp_4_cfg_w,
  input io_ptw_pmp_4_cfg_r,
  input [29:0] io_ptw_pmp_4_addr,
  input [31:0] io_ptw_pmp_4_mask,
  input io_ptw_pmp_5_cfg_l,
  input [1:0] io_ptw_pmp_5_cfg_a,
  input io_ptw_pmp_5_cfg_x,
  input io_ptw_pmp_5_cfg_w,
  input io_ptw_pmp_5_cfg_r,
  input [29:0] io_ptw_pmp_5_addr,
  input [31:0] io_ptw_pmp_5_mask,
  input io_ptw_pmp_6_cfg_l,
  input [1:0] io_ptw_pmp_6_cfg_a,
  input io_ptw_pmp_6_cfg_x,
  input io_ptw_pmp_6_cfg_w,
  input io_ptw_pmp_6_cfg_r,
  input [29:0] io_ptw_pmp_6_addr,
  input [31:0] io_ptw_pmp_6_mask,
  input io_ptw_pmp_7_cfg_l,
  input [1:0] io_ptw_pmp_7_cfg_a,
  input io_ptw_pmp_7_cfg_x,
  input io_ptw_pmp_7_cfg_w,
  input io_ptw_pmp_7_cfg_r,
  input [29:0] io_ptw_pmp_7_addr,
  input [31:0] io_ptw_pmp_7_mask,
  input io_kill,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [19:0] mpu_ppn_barrier_io_x_ppn ;  
   wire mpu_ppn_barrier_io_x_u ;  
   wire mpu_ppn_barrier_io_x_ae ;  
   wire mpu_ppn_barrier_io_x_sw ;  
   wire mpu_ppn_barrier_io_x_sx ;  
   wire mpu_ppn_barrier_io_x_sr ;  
   wire mpu_ppn_barrier_io_x_pw ;  
   wire mpu_ppn_barrier_io_x_px ;  
   wire mpu_ppn_barrier_io_x_pr ;  
   wire mpu_ppn_barrier_io_x_ppp ;  
   wire mpu_ppn_barrier_io_x_pal ;  
   wire mpu_ppn_barrier_io_x_paa ;  
   wire mpu_ppn_barrier_io_x_eff ;  
   wire mpu_ppn_barrier_io_x_c ;  
   wire [19:0] mpu_ppn_barrier_io_y_ppn ;  
   wire mpu_ppn_barrier_io_y_u ;  
   wire mpu_ppn_barrier_io_y_ae ;  
   wire mpu_ppn_barrier_io_y_sw ;  
   wire mpu_ppn_barrier_io_y_sx ;  
   wire mpu_ppn_barrier_io_y_sr ;  
   wire mpu_ppn_barrier_io_y_pw ;  
   wire mpu_ppn_barrier_io_y_px ;  
   wire mpu_ppn_barrier_io_y_pr ;  
   wire mpu_ppn_barrier_io_y_ppp ;  
   wire mpu_ppn_barrier_io_y_pal ;  
   wire mpu_ppn_barrier_io_y_paa ;  
   wire mpu_ppn_barrier_io_y_eff ;  
   wire mpu_ppn_barrier_io_y_c ;  
   wire [29:0] mpu_ppn_barrier_io_covSum ;  
   wire mpu_ppn_barrier_metaAssert ;  
   wire [1:0] pmp_io_prv ;  
   wire pmp_io_pmp_0_cfg_l ;  
   wire [1:0] pmp_io_pmp_0_cfg_a ;  
   wire pmp_io_pmp_0_cfg_x ;  
   wire pmp_io_pmp_0_cfg_w ;  
   wire pmp_io_pmp_0_cfg_r ;  
   wire [29:0] pmp_io_pmp_0_addr ;  
   wire [31:0] pmp_io_pmp_0_mask ;  
   wire pmp_io_pmp_1_cfg_l ;  
   wire [1:0] pmp_io_pmp_1_cfg_a ;  
   wire pmp_io_pmp_1_cfg_x ;  
   wire pmp_io_pmp_1_cfg_w ;  
   wire pmp_io_pmp_1_cfg_r ;  
   wire [29:0] pmp_io_pmp_1_addr ;  
   wire [31:0] pmp_io_pmp_1_mask ;  
   wire pmp_io_pmp_2_cfg_l ;  
   wire [1:0] pmp_io_pmp_2_cfg_a ;  
   wire pmp_io_pmp_2_cfg_x ;  
   wire pmp_io_pmp_2_cfg_w ;  
   wire pmp_io_pmp_2_cfg_r ;  
   wire [29:0] pmp_io_pmp_2_addr ;  
   wire [31:0] pmp_io_pmp_2_mask ;  
   wire pmp_io_pmp_3_cfg_l ;  
   wire [1:0] pmp_io_pmp_3_cfg_a ;  
   wire pmp_io_pmp_3_cfg_x ;  
   wire pmp_io_pmp_3_cfg_w ;  
   wire pmp_io_pmp_3_cfg_r ;  
   wire [29:0] pmp_io_pmp_3_addr ;  
   wire [31:0] pmp_io_pmp_3_mask ;  
   wire pmp_io_pmp_4_cfg_l ;  
   wire [1:0] pmp_io_pmp_4_cfg_a ;  
   wire pmp_io_pmp_4_cfg_x ;  
   wire pmp_io_pmp_4_cfg_w ;  
   wire pmp_io_pmp_4_cfg_r ;  
   wire [29:0] pmp_io_pmp_4_addr ;  
   wire [31:0] pmp_io_pmp_4_mask ;  
   wire pmp_io_pmp_5_cfg_l ;  
   wire [1:0] pmp_io_pmp_5_cfg_a ;  
   wire pmp_io_pmp_5_cfg_x ;  
   wire pmp_io_pmp_5_cfg_w ;  
   wire pmp_io_pmp_5_cfg_r ;  
   wire [29:0] pmp_io_pmp_5_addr ;  
   wire [31:0] pmp_io_pmp_5_mask ;  
   wire pmp_io_pmp_6_cfg_l ;  
   wire [1:0] pmp_io_pmp_6_cfg_a ;  
   wire pmp_io_pmp_6_cfg_x ;  
   wire pmp_io_pmp_6_cfg_w ;  
   wire pmp_io_pmp_6_cfg_r ;  
   wire [29:0] pmp_io_pmp_6_addr ;  
   wire [31:0] pmp_io_pmp_6_mask ;  
   wire pmp_io_pmp_7_cfg_l ;  
   wire [1:0] pmp_io_pmp_7_cfg_a ;  
   wire pmp_io_pmp_7_cfg_x ;  
   wire pmp_io_pmp_7_cfg_w ;  
   wire pmp_io_pmp_7_cfg_r ;  
   wire [29:0] pmp_io_pmp_7_addr ;  
   wire [31:0] pmp_io_pmp_7_mask ;  
   wire [31:0] pmp_io_addr ;  
   wire pmp_io_r ;  
   wire pmp_io_w ;  
   wire pmp_io_x ;  
   wire [29:0] pmp_io_covSum ;  
   wire pmp_metaAssert ;  
   wire [19:0] entries_barrier_io_x_ppn ;  
   wire entries_barrier_io_x_u ;  
   wire entries_barrier_io_x_ae ;  
   wire entries_barrier_io_x_sw ;  
   wire entries_barrier_io_x_sx ;  
   wire entries_barrier_io_x_sr ;  
   wire entries_barrier_io_x_pw ;  
   wire entries_barrier_io_x_px ;  
   wire entries_barrier_io_x_pr ;  
   wire entries_barrier_io_x_ppp ;  
   wire entries_barrier_io_x_pal ;  
   wire entries_barrier_io_x_paa ;  
   wire entries_barrier_io_x_eff ;  
   wire entries_barrier_io_x_c ;  
   wire [19:0] entries_barrier_io_y_ppn ;  
   wire entries_barrier_io_y_u ;  
   wire entries_barrier_io_y_ae ;  
   wire entries_barrier_io_y_sw ;  
   wire entries_barrier_io_y_sx ;  
   wire entries_barrier_io_y_sr ;  
   wire entries_barrier_io_y_pw ;  
   wire entries_barrier_io_y_px ;  
   wire entries_barrier_io_y_pr ;  
   wire entries_barrier_io_y_ppp ;  
   wire entries_barrier_io_y_pal ;  
   wire entries_barrier_io_y_paa ;  
   wire entries_barrier_io_y_eff ;  
   wire entries_barrier_io_y_c ;  
   wire [29:0] entries_barrier_io_covSum ;  
   wire entries_barrier_metaAssert ;  
   wire [19:0] entries_barrier_1_io_x_ppn ;  
   wire entries_barrier_1_io_x_u ;  
   wire entries_barrier_1_io_x_ae ;  
   wire entries_barrier_1_io_x_sw ;  
   wire entries_barrier_1_io_x_sx ;  
   wire entries_barrier_1_io_x_sr ;  
   wire entries_barrier_1_io_x_pw ;  
   wire entries_barrier_1_io_x_px ;  
   wire entries_barrier_1_io_x_pr ;  
   wire entries_barrier_1_io_x_ppp ;  
   wire entries_barrier_1_io_x_pal ;  
   wire entries_barrier_1_io_x_paa ;  
   wire entries_barrier_1_io_x_eff ;  
   wire entries_barrier_1_io_x_c ;  
   wire [19:0] entries_barrier_1_io_y_ppn ;  
   wire entries_barrier_1_io_y_u ;  
   wire entries_barrier_1_io_y_ae ;  
   wire entries_barrier_1_io_y_sw ;  
   wire entries_barrier_1_io_y_sx ;  
   wire entries_barrier_1_io_y_sr ;  
   wire entries_barrier_1_io_y_pw ;  
   wire entries_barrier_1_io_y_px ;  
   wire entries_barrier_1_io_y_pr ;  
   wire entries_barrier_1_io_y_ppp ;  
   wire entries_barrier_1_io_y_pal ;  
   wire entries_barrier_1_io_y_paa ;  
   wire entries_barrier_1_io_y_eff ;  
   wire entries_barrier_1_io_y_c ;  
   wire [29:0] entries_barrier_1_io_covSum ;  
   wire entries_barrier_1_metaAssert ;  
   wire [19:0] entries_barrier_2_io_x_ppn ;  
   wire entries_barrier_2_io_x_u ;  
   wire entries_barrier_2_io_x_ae ;  
   wire entries_barrier_2_io_x_sw ;  
   wire entries_barrier_2_io_x_sx ;  
   wire entries_barrier_2_io_x_sr ;  
   wire entries_barrier_2_io_x_pw ;  
   wire entries_barrier_2_io_x_px ;  
   wire entries_barrier_2_io_x_pr ;  
   wire entries_barrier_2_io_x_ppp ;  
   wire entries_barrier_2_io_x_pal ;  
   wire entries_barrier_2_io_x_paa ;  
   wire entries_barrier_2_io_x_eff ;  
   wire entries_barrier_2_io_x_c ;  
   wire [19:0] entries_barrier_2_io_y_ppn ;  
   wire entries_barrier_2_io_y_u ;  
   wire entries_barrier_2_io_y_ae ;  
   wire entries_barrier_2_io_y_sw ;  
   wire entries_barrier_2_io_y_sx ;  
   wire entries_barrier_2_io_y_sr ;  
   wire entries_barrier_2_io_y_pw ;  
   wire entries_barrier_2_io_y_px ;  
   wire entries_barrier_2_io_y_pr ;  
   wire entries_barrier_2_io_y_ppp ;  
   wire entries_barrier_2_io_y_pal ;  
   wire entries_barrier_2_io_y_paa ;  
   wire entries_barrier_2_io_y_eff ;  
   wire entries_barrier_2_io_y_c ;  
   wire [29:0] entries_barrier_2_io_covSum ;  
   wire entries_barrier_2_metaAssert ;  
   wire [19:0] entries_barrier_3_io_x_ppn ;  
   wire entries_barrier_3_io_x_u ;  
   wire entries_barrier_3_io_x_ae ;  
   wire entries_barrier_3_io_x_sw ;  
   wire entries_barrier_3_io_x_sx ;  
   wire entries_barrier_3_io_x_sr ;  
   wire entries_barrier_3_io_x_pw ;  
   wire entries_barrier_3_io_x_px ;  
   wire entries_barrier_3_io_x_pr ;  
   wire entries_barrier_3_io_x_ppp ;  
   wire entries_barrier_3_io_x_pal ;  
   wire entries_barrier_3_io_x_paa ;  
   wire entries_barrier_3_io_x_eff ;  
   wire entries_barrier_3_io_x_c ;  
   wire [19:0] entries_barrier_3_io_y_ppn ;  
   wire entries_barrier_3_io_y_u ;  
   wire entries_barrier_3_io_y_ae ;  
   wire entries_barrier_3_io_y_sw ;  
   wire entries_barrier_3_io_y_sx ;  
   wire entries_barrier_3_io_y_sr ;  
   wire entries_barrier_3_io_y_pw ;  
   wire entries_barrier_3_io_y_px ;  
   wire entries_barrier_3_io_y_pr ;  
   wire entries_barrier_3_io_y_ppp ;  
   wire entries_barrier_3_io_y_pal ;  
   wire entries_barrier_3_io_y_paa ;  
   wire entries_barrier_3_io_y_eff ;  
   wire entries_barrier_3_io_y_c ;  
   wire [29:0] entries_barrier_3_io_covSum ;  
   wire entries_barrier_3_metaAssert ;  
   wire [19:0] entries_barrier_4_io_x_ppn ;  
   wire entries_barrier_4_io_x_u ;  
   wire entries_barrier_4_io_x_ae ;  
   wire entries_barrier_4_io_x_sw ;  
   wire entries_barrier_4_io_x_sx ;  
   wire entries_barrier_4_io_x_sr ;  
   wire entries_barrier_4_io_x_pw ;  
   wire entries_barrier_4_io_x_px ;  
   wire entries_barrier_4_io_x_pr ;  
   wire entries_barrier_4_io_x_ppp ;  
   wire entries_barrier_4_io_x_pal ;  
   wire entries_barrier_4_io_x_paa ;  
   wire entries_barrier_4_io_x_eff ;  
   wire entries_barrier_4_io_x_c ;  
   wire [19:0] entries_barrier_4_io_y_ppn ;  
   wire entries_barrier_4_io_y_u ;  
   wire entries_barrier_4_io_y_ae ;  
   wire entries_barrier_4_io_y_sw ;  
   wire entries_barrier_4_io_y_sx ;  
   wire entries_barrier_4_io_y_sr ;  
   wire entries_barrier_4_io_y_pw ;  
   wire entries_barrier_4_io_y_px ;  
   wire entries_barrier_4_io_y_pr ;  
   wire entries_barrier_4_io_y_ppp ;  
   wire entries_barrier_4_io_y_pal ;  
   wire entries_barrier_4_io_y_paa ;  
   wire entries_barrier_4_io_y_eff ;  
   wire entries_barrier_4_io_y_c ;  
   wire [29:0] entries_barrier_4_io_covSum ;  
   wire entries_barrier_4_metaAssert ;  
   wire [19:0] entries_barrier_5_io_x_ppn ;  
   wire entries_barrier_5_io_x_u ;  
   wire entries_barrier_5_io_x_ae ;  
   wire entries_barrier_5_io_x_sw ;  
   wire entries_barrier_5_io_x_sx ;  
   wire entries_barrier_5_io_x_sr ;  
   wire entries_barrier_5_io_x_pw ;  
   wire entries_barrier_5_io_x_px ;  
   wire entries_barrier_5_io_x_pr ;  
   wire entries_barrier_5_io_x_ppp ;  
   wire entries_barrier_5_io_x_pal ;  
   wire entries_barrier_5_io_x_paa ;  
   wire entries_barrier_5_io_x_eff ;  
   wire entries_barrier_5_io_x_c ;  
   wire [19:0] entries_barrier_5_io_y_ppn ;  
   wire entries_barrier_5_io_y_u ;  
   wire entries_barrier_5_io_y_ae ;  
   wire entries_barrier_5_io_y_sw ;  
   wire entries_barrier_5_io_y_sx ;  
   wire entries_barrier_5_io_y_sr ;  
   wire entries_barrier_5_io_y_pw ;  
   wire entries_barrier_5_io_y_px ;  
   wire entries_barrier_5_io_y_pr ;  
   wire entries_barrier_5_io_y_ppp ;  
   wire entries_barrier_5_io_y_pal ;  
   wire entries_barrier_5_io_y_paa ;  
   wire entries_barrier_5_io_y_eff ;  
   wire entries_barrier_5_io_y_c ;  
   wire [29:0] entries_barrier_5_io_covSum ;  
   wire entries_barrier_5_metaAssert ;  
   wire [19:0] entries_barrier_6_io_x_ppn ;  
   wire entries_barrier_6_io_x_u ;  
   wire entries_barrier_6_io_x_ae ;  
   wire entries_barrier_6_io_x_sw ;  
   wire entries_barrier_6_io_x_sx ;  
   wire entries_barrier_6_io_x_sr ;  
   wire entries_barrier_6_io_x_pw ;  
   wire entries_barrier_6_io_x_px ;  
   wire entries_barrier_6_io_x_pr ;  
   wire entries_barrier_6_io_x_ppp ;  
   wire entries_barrier_6_io_x_pal ;  
   wire entries_barrier_6_io_x_paa ;  
   wire entries_barrier_6_io_x_eff ;  
   wire entries_barrier_6_io_x_c ;  
   wire [19:0] entries_barrier_6_io_y_ppn ;  
   wire entries_barrier_6_io_y_u ;  
   wire entries_barrier_6_io_y_ae ;  
   wire entries_barrier_6_io_y_sw ;  
   wire entries_barrier_6_io_y_sx ;  
   wire entries_barrier_6_io_y_sr ;  
   wire entries_barrier_6_io_y_pw ;  
   wire entries_barrier_6_io_y_px ;  
   wire entries_barrier_6_io_y_pr ;  
   wire entries_barrier_6_io_y_ppp ;  
   wire entries_barrier_6_io_y_pal ;  
   wire entries_barrier_6_io_y_paa ;  
   wire entries_barrier_6_io_y_eff ;  
   wire entries_barrier_6_io_y_c ;  
   wire [29:0] entries_barrier_6_io_covSum ;  
   wire entries_barrier_6_metaAssert ;  
   wire [19:0] entries_barrier_7_io_x_ppn ;  
   wire entries_barrier_7_io_x_u ;  
   wire entries_barrier_7_io_x_ae ;  
   wire entries_barrier_7_io_x_sw ;  
   wire entries_barrier_7_io_x_sx ;  
   wire entries_barrier_7_io_x_sr ;  
   wire entries_barrier_7_io_x_pw ;  
   wire entries_barrier_7_io_x_px ;  
   wire entries_barrier_7_io_x_pr ;  
   wire entries_barrier_7_io_x_ppp ;  
   wire entries_barrier_7_io_x_pal ;  
   wire entries_barrier_7_io_x_paa ;  
   wire entries_barrier_7_io_x_eff ;  
   wire entries_barrier_7_io_x_c ;  
   wire [19:0] entries_barrier_7_io_y_ppn ;  
   wire entries_barrier_7_io_y_u ;  
   wire entries_barrier_7_io_y_ae ;  
   wire entries_barrier_7_io_y_sw ;  
   wire entries_barrier_7_io_y_sx ;  
   wire entries_barrier_7_io_y_sr ;  
   wire entries_barrier_7_io_y_pw ;  
   wire entries_barrier_7_io_y_px ;  
   wire entries_barrier_7_io_y_pr ;  
   wire entries_barrier_7_io_y_ppp ;  
   wire entries_barrier_7_io_y_pal ;  
   wire entries_barrier_7_io_y_paa ;  
   wire entries_barrier_7_io_y_eff ;  
   wire entries_barrier_7_io_y_c ;  
   wire [29:0] entries_barrier_7_io_covSum ;  
   wire entries_barrier_7_metaAssert ;  
   wire [19:0] entries_barrier_8_io_x_ppn ;  
   wire entries_barrier_8_io_x_u ;  
   wire entries_barrier_8_io_x_ae ;  
   wire entries_barrier_8_io_x_sw ;  
   wire entries_barrier_8_io_x_sx ;  
   wire entries_barrier_8_io_x_sr ;  
   wire entries_barrier_8_io_x_pw ;  
   wire entries_barrier_8_io_x_px ;  
   wire entries_barrier_8_io_x_pr ;  
   wire entries_barrier_8_io_x_ppp ;  
   wire entries_barrier_8_io_x_pal ;  
   wire entries_barrier_8_io_x_paa ;  
   wire entries_barrier_8_io_x_eff ;  
   wire entries_barrier_8_io_x_c ;  
   wire [19:0] entries_barrier_8_io_y_ppn ;  
   wire entries_barrier_8_io_y_u ;  
   wire entries_barrier_8_io_y_ae ;  
   wire entries_barrier_8_io_y_sw ;  
   wire entries_barrier_8_io_y_sx ;  
   wire entries_barrier_8_io_y_sr ;  
   wire entries_barrier_8_io_y_pw ;  
   wire entries_barrier_8_io_y_px ;  
   wire entries_barrier_8_io_y_pr ;  
   wire entries_barrier_8_io_y_ppp ;  
   wire entries_barrier_8_io_y_pal ;  
   wire entries_barrier_8_io_y_paa ;  
   wire entries_barrier_8_io_y_eff ;  
   wire entries_barrier_8_io_y_c ;  
   wire [29:0] entries_barrier_8_io_covSum ;  
   wire entries_barrier_8_metaAssert ;  
   wire [19:0] entries_barrier_9_io_x_ppn ;  
   wire entries_barrier_9_io_x_u ;  
   wire entries_barrier_9_io_x_ae ;  
   wire entries_barrier_9_io_x_sw ;  
   wire entries_barrier_9_io_x_sx ;  
   wire entries_barrier_9_io_x_sr ;  
   wire entries_barrier_9_io_x_pw ;  
   wire entries_barrier_9_io_x_px ;  
   wire entries_barrier_9_io_x_pr ;  
   wire entries_barrier_9_io_x_ppp ;  
   wire entries_barrier_9_io_x_pal ;  
   wire entries_barrier_9_io_x_paa ;  
   wire entries_barrier_9_io_x_eff ;  
   wire entries_barrier_9_io_x_c ;  
   wire [19:0] entries_barrier_9_io_y_ppn ;  
   wire entries_barrier_9_io_y_u ;  
   wire entries_barrier_9_io_y_ae ;  
   wire entries_barrier_9_io_y_sw ;  
   wire entries_barrier_9_io_y_sx ;  
   wire entries_barrier_9_io_y_sr ;  
   wire entries_barrier_9_io_y_pw ;  
   wire entries_barrier_9_io_y_px ;  
   wire entries_barrier_9_io_y_pr ;  
   wire entries_barrier_9_io_y_ppp ;  
   wire entries_barrier_9_io_y_pal ;  
   wire entries_barrier_9_io_y_paa ;  
   wire entries_barrier_9_io_y_eff ;  
   wire entries_barrier_9_io_y_c ;  
   wire [29:0] entries_barrier_9_io_covSum ;  
   wire entries_barrier_9_metaAssert ;  
   wire [19:0] entries_barrier_10_io_x_ppn ;  
   wire entries_barrier_10_io_x_u ;  
   wire entries_barrier_10_io_x_ae ;  
   wire entries_barrier_10_io_x_sw ;  
   wire entries_barrier_10_io_x_sx ;  
   wire entries_barrier_10_io_x_sr ;  
   wire entries_barrier_10_io_x_pw ;  
   wire entries_barrier_10_io_x_px ;  
   wire entries_barrier_10_io_x_pr ;  
   wire entries_barrier_10_io_x_ppp ;  
   wire entries_barrier_10_io_x_pal ;  
   wire entries_barrier_10_io_x_paa ;  
   wire entries_barrier_10_io_x_eff ;  
   wire entries_barrier_10_io_x_c ;  
   wire [19:0] entries_barrier_10_io_y_ppn ;  
   wire entries_barrier_10_io_y_u ;  
   wire entries_barrier_10_io_y_ae ;  
   wire entries_barrier_10_io_y_sw ;  
   wire entries_barrier_10_io_y_sx ;  
   wire entries_barrier_10_io_y_sr ;  
   wire entries_barrier_10_io_y_pw ;  
   wire entries_barrier_10_io_y_px ;  
   wire entries_barrier_10_io_y_pr ;  
   wire entries_barrier_10_io_y_ppp ;  
   wire entries_barrier_10_io_y_pal ;  
   wire entries_barrier_10_io_y_paa ;  
   wire entries_barrier_10_io_y_eff ;  
   wire entries_barrier_10_io_y_c ;  
   wire [29:0] entries_barrier_10_io_covSum ;  
   wire entries_barrier_10_metaAssert ;  
   wire [19:0] entries_barrier_11_io_x_ppn ;  
   wire entries_barrier_11_io_x_u ;  
   wire entries_barrier_11_io_x_ae ;  
   wire entries_barrier_11_io_x_sw ;  
   wire entries_barrier_11_io_x_sx ;  
   wire entries_barrier_11_io_x_sr ;  
   wire entries_barrier_11_io_x_pw ;  
   wire entries_barrier_11_io_x_px ;  
   wire entries_barrier_11_io_x_pr ;  
   wire entries_barrier_11_io_x_ppp ;  
   wire entries_barrier_11_io_x_pal ;  
   wire entries_barrier_11_io_x_paa ;  
   wire entries_barrier_11_io_x_eff ;  
   wire entries_barrier_11_io_x_c ;  
   wire [19:0] entries_barrier_11_io_y_ppn ;  
   wire entries_barrier_11_io_y_u ;  
   wire entries_barrier_11_io_y_ae ;  
   wire entries_barrier_11_io_y_sw ;  
   wire entries_barrier_11_io_y_sx ;  
   wire entries_barrier_11_io_y_sr ;  
   wire entries_barrier_11_io_y_pw ;  
   wire entries_barrier_11_io_y_px ;  
   wire entries_barrier_11_io_y_pr ;  
   wire entries_barrier_11_io_y_ppp ;  
   wire entries_barrier_11_io_y_pal ;  
   wire entries_barrier_11_io_y_paa ;  
   wire entries_barrier_11_io_y_eff ;  
   wire entries_barrier_11_io_y_c ;  
   wire [29:0] entries_barrier_11_io_covSum ;  
   wire entries_barrier_11_metaAssert ;  
   wire [19:0] entries_barrier_12_io_x_ppn ;  
   wire entries_barrier_12_io_x_u ;  
   wire entries_barrier_12_io_x_ae ;  
   wire entries_barrier_12_io_x_sw ;  
   wire entries_barrier_12_io_x_sx ;  
   wire entries_barrier_12_io_x_sr ;  
   wire entries_barrier_12_io_x_pw ;  
   wire entries_barrier_12_io_x_px ;  
   wire entries_barrier_12_io_x_pr ;  
   wire entries_barrier_12_io_x_ppp ;  
   wire entries_barrier_12_io_x_pal ;  
   wire entries_barrier_12_io_x_paa ;  
   wire entries_barrier_12_io_x_eff ;  
   wire entries_barrier_12_io_x_c ;  
   wire [19:0] entries_barrier_12_io_y_ppn ;  
   wire entries_barrier_12_io_y_u ;  
   wire entries_barrier_12_io_y_ae ;  
   wire entries_barrier_12_io_y_sw ;  
   wire entries_barrier_12_io_y_sx ;  
   wire entries_barrier_12_io_y_sr ;  
   wire entries_barrier_12_io_y_pw ;  
   wire entries_barrier_12_io_y_px ;  
   wire entries_barrier_12_io_y_pr ;  
   wire entries_barrier_12_io_y_ppp ;  
   wire entries_barrier_12_io_y_pal ;  
   wire entries_barrier_12_io_y_paa ;  
   wire entries_barrier_12_io_y_eff ;  
   wire entries_barrier_12_io_y_c ;  
   wire [29:0] entries_barrier_12_io_covSum ;  
   wire entries_barrier_12_metaAssert ;  
   wire [26:0] vpn ;  
   reg [26:0] sectored_entries_0_0_tag ;  
   reg [31:0] _RAND_0 ;  
   reg [34:0] sectored_entries_0_0_data_0 ;  
   reg [63:0] _RAND_1 ;  
   reg [34:0] sectored_entries_0_0_data_1 ;  
   reg [63:0] _RAND_2 ;  
   reg [34:0] sectored_entries_0_0_data_2 ;  
   reg [63:0] _RAND_3 ;  
   reg [34:0] sectored_entries_0_0_data_3 ;  
   reg [63:0] _RAND_4 ;  
   reg sectored_entries_0_0_valid_0 ;  
   reg [31:0] _RAND_5 ;  
   reg sectored_entries_0_0_valid_1 ;  
   reg [31:0] _RAND_6 ;  
   reg sectored_entries_0_0_valid_2 ;  
   reg [31:0] _RAND_7 ;  
   reg sectored_entries_0_0_valid_3 ;  
   reg [31:0] _RAND_8 ;  
   reg [26:0] sectored_entries_0_1_tag ;  
   reg [31:0] _RAND_9 ;  
   reg [34:0] sectored_entries_0_1_data_0 ;  
   reg [63:0] _RAND_10 ;  
   reg [34:0] sectored_entries_0_1_data_1 ;  
   reg [63:0] _RAND_11 ;  
   reg [34:0] sectored_entries_0_1_data_2 ;  
   reg [63:0] _RAND_12 ;  
   reg [34:0] sectored_entries_0_1_data_3 ;  
   reg [63:0] _RAND_13 ;  
   reg sectored_entries_0_1_valid_0 ;  
   reg [31:0] _RAND_14 ;  
   reg sectored_entries_0_1_valid_1 ;  
   reg [31:0] _RAND_15 ;  
   reg sectored_entries_0_1_valid_2 ;  
   reg [31:0] _RAND_16 ;  
   reg sectored_entries_0_1_valid_3 ;  
   reg [31:0] _RAND_17 ;  
   reg [26:0] sectored_entries_0_2_tag ;  
   reg [31:0] _RAND_18 ;  
   reg [34:0] sectored_entries_0_2_data_0 ;  
   reg [63:0] _RAND_19 ;  
   reg [34:0] sectored_entries_0_2_data_1 ;  
   reg [63:0] _RAND_20 ;  
   reg [34:0] sectored_entries_0_2_data_2 ;  
   reg [63:0] _RAND_21 ;  
   reg [34:0] sectored_entries_0_2_data_3 ;  
   reg [63:0] _RAND_22 ;  
   reg sectored_entries_0_2_valid_0 ;  
   reg [31:0] _RAND_23 ;  
   reg sectored_entries_0_2_valid_1 ;  
   reg [31:0] _RAND_24 ;  
   reg sectored_entries_0_2_valid_2 ;  
   reg [31:0] _RAND_25 ;  
   reg sectored_entries_0_2_valid_3 ;  
   reg [31:0] _RAND_26 ;  
   reg [26:0] sectored_entries_0_3_tag ;  
   reg [31:0] _RAND_27 ;  
   reg [34:0] sectored_entries_0_3_data_0 ;  
   reg [63:0] _RAND_28 ;  
   reg [34:0] sectored_entries_0_3_data_1 ;  
   reg [63:0] _RAND_29 ;  
   reg [34:0] sectored_entries_0_3_data_2 ;  
   reg [63:0] _RAND_30 ;  
   reg [34:0] sectored_entries_0_3_data_3 ;  
   reg [63:0] _RAND_31 ;  
   reg sectored_entries_0_3_valid_0 ;  
   reg [31:0] _RAND_32 ;  
   reg sectored_entries_0_3_valid_1 ;  
   reg [31:0] _RAND_33 ;  
   reg sectored_entries_0_3_valid_2 ;  
   reg [31:0] _RAND_34 ;  
   reg sectored_entries_0_3_valid_3 ;  
   reg [31:0] _RAND_35 ;  
   reg [26:0] sectored_entries_0_4_tag ;  
   reg [31:0] _RAND_36 ;  
   reg [34:0] sectored_entries_0_4_data_0 ;  
   reg [63:0] _RAND_37 ;  
   reg [34:0] sectored_entries_0_4_data_1 ;  
   reg [63:0] _RAND_38 ;  
   reg [34:0] sectored_entries_0_4_data_2 ;  
   reg [63:0] _RAND_39 ;  
   reg [34:0] sectored_entries_0_4_data_3 ;  
   reg [63:0] _RAND_40 ;  
   reg sectored_entries_0_4_valid_0 ;  
   reg [31:0] _RAND_41 ;  
   reg sectored_entries_0_4_valid_1 ;  
   reg [31:0] _RAND_42 ;  
   reg sectored_entries_0_4_valid_2 ;  
   reg [31:0] _RAND_43 ;  
   reg sectored_entries_0_4_valid_3 ;  
   reg [31:0] _RAND_44 ;  
   reg [26:0] sectored_entries_0_5_tag ;  
   reg [31:0] _RAND_45 ;  
   reg [34:0] sectored_entries_0_5_data_0 ;  
   reg [63:0] _RAND_46 ;  
   reg [34:0] sectored_entries_0_5_data_1 ;  
   reg [63:0] _RAND_47 ;  
   reg [34:0] sectored_entries_0_5_data_2 ;  
   reg [63:0] _RAND_48 ;  
   reg [34:0] sectored_entries_0_5_data_3 ;  
   reg [63:0] _RAND_49 ;  
   reg sectored_entries_0_5_valid_0 ;  
   reg [31:0] _RAND_50 ;  
   reg sectored_entries_0_5_valid_1 ;  
   reg [31:0] _RAND_51 ;  
   reg sectored_entries_0_5_valid_2 ;  
   reg [31:0] _RAND_52 ;  
   reg sectored_entries_0_5_valid_3 ;  
   reg [31:0] _RAND_53 ;  
   reg [26:0] sectored_entries_0_6_tag ;  
   reg [31:0] _RAND_54 ;  
   reg [34:0] sectored_entries_0_6_data_0 ;  
   reg [63:0] _RAND_55 ;  
   reg [34:0] sectored_entries_0_6_data_1 ;  
   reg [63:0] _RAND_56 ;  
   reg [34:0] sectored_entries_0_6_data_2 ;  
   reg [63:0] _RAND_57 ;  
   reg [34:0] sectored_entries_0_6_data_3 ;  
   reg [63:0] _RAND_58 ;  
   reg sectored_entries_0_6_valid_0 ;  
   reg [31:0] _RAND_59 ;  
   reg sectored_entries_0_6_valid_1 ;  
   reg [31:0] _RAND_60 ;  
   reg sectored_entries_0_6_valid_2 ;  
   reg [31:0] _RAND_61 ;  
   reg sectored_entries_0_6_valid_3 ;  
   reg [31:0] _RAND_62 ;  
   reg [26:0] sectored_entries_0_7_tag ;  
   reg [31:0] _RAND_63 ;  
   reg [34:0] sectored_entries_0_7_data_0 ;  
   reg [63:0] _RAND_64 ;  
   reg [34:0] sectored_entries_0_7_data_1 ;  
   reg [63:0] _RAND_65 ;  
   reg [34:0] sectored_entries_0_7_data_2 ;  
   reg [63:0] _RAND_66 ;  
   reg [34:0] sectored_entries_0_7_data_3 ;  
   reg [63:0] _RAND_67 ;  
   reg sectored_entries_0_7_valid_0 ;  
   reg [31:0] _RAND_68 ;  
   reg sectored_entries_0_7_valid_1 ;  
   reg [31:0] _RAND_69 ;  
   reg sectored_entries_0_7_valid_2 ;  
   reg [31:0] _RAND_70 ;  
   reg sectored_entries_0_7_valid_3 ;  
   reg [31:0] _RAND_71 ;  
   reg [1:0] superpage_entries_0_level ;  
   reg [31:0] _RAND_72 ;  
   reg [26:0] superpage_entries_0_tag ;  
   reg [31:0] _RAND_73 ;  
   reg [34:0] superpage_entries_0_data_0 ;  
   reg [63:0] _RAND_74 ;  
   reg superpage_entries_0_valid_0 ;  
   reg [31:0] _RAND_75 ;  
   reg [1:0] superpage_entries_1_level ;  
   reg [31:0] _RAND_76 ;  
   reg [26:0] superpage_entries_1_tag ;  
   reg [31:0] _RAND_77 ;  
   reg [34:0] superpage_entries_1_data_0 ;  
   reg [63:0] _RAND_78 ;  
   reg superpage_entries_1_valid_0 ;  
   reg [31:0] _RAND_79 ;  
   reg [1:0] superpage_entries_2_level ;  
   reg [31:0] _RAND_80 ;  
   reg [26:0] superpage_entries_2_tag ;  
   reg [31:0] _RAND_81 ;  
   reg [34:0] superpage_entries_2_data_0 ;  
   reg [63:0] _RAND_82 ;  
   reg superpage_entries_2_valid_0 ;  
   reg [31:0] _RAND_83 ;  
   reg [1:0] superpage_entries_3_level ;  
   reg [31:0] _RAND_84 ;  
   reg [26:0] superpage_entries_3_tag ;  
   reg [31:0] _RAND_85 ;  
   reg [34:0] superpage_entries_3_data_0 ;  
   reg [63:0] _RAND_86 ;  
   reg superpage_entries_3_valid_0 ;  
   reg [31:0] _RAND_87 ;  
   reg [1:0] special_entry_level ;  
   reg [31:0] _RAND_88 ;  
   reg [26:0] special_entry_tag ;  
   reg [31:0] _RAND_89 ;  
   reg [34:0] special_entry_data_0 ;  
   reg [63:0] _RAND_90 ;  
   reg special_entry_valid_0 ;  
   reg [31:0] _RAND_91 ;  
   reg [1:0] state ;  
   reg [31:0] _RAND_92 ;  
   reg [26:0] r_refill_tag ;  
   reg [31:0] _RAND_93 ;  
   reg [1:0] r_superpage_repl_addr ;  
   reg [31:0] _RAND_94 ;  
   reg [2:0] r_sectored_repl_addr ;  
   reg [31:0] _RAND_95 ;  
   reg [2:0] r_sectored_hit_addr ;  
   reg [31:0] _RAND_96 ;  
   reg r_sectored_hit ;  
   reg [31:0] _RAND_97 ;  
   wire priv_s ;  
   wire priv_uses_vm ;  
   wire vm_enabled ;  
   wire [19:0] refill_ppn ;  
   wire _invalidate_refill_T ;  
   wire _invalidate_refill_T_1 ;  
   wire _invalidate_refill_T_2 ;  
   wire invalidate_refill ;  
   wire [1:0] mpu_ppn_hi ;  
   wire mpu_ppn_ignore ;  
   wire [26:0] _mpu_ppn_T_17 ;  
   wire [26:0] _GEN_919 ;  
   wire [26:0] _mpu_ppn_T_18 ;  
   wire [8:0] mpu_ppn_lo ;  
   wire mpu_ppn_ignore_1 ;  
   wire [26:0] _mpu_ppn_T_19 ;  
   wire [26:0] _mpu_ppn_T_20 ;  
   wire [8:0] mpu_ppn_lo_1 ;  
   wire [19:0] _mpu_ppn_T_21 ;  
   wire [27:0] _mpu_ppn_T_23 ;  
   wire [27:0] mpu_ppn ;  
   wire [11:0] mpu_physaddr_lo ;  
   wire [39:0] mpu_physaddr ;  
   wire [2:0] _mpu_priv_T_2 ;  
   wire [2:0] mpu_priv ;  
   wire [39:0] _legal_address_T ;  
   wire [40:0] _legal_address_T_1 ;  
   wire [40:0] _legal_address_T_3 ;  
   wire _legal_address_T_4 ;  
   wire [39:0] _legal_address_T_5 ;  
   wire [40:0] _legal_address_T_6 ;  
   wire [40:0] _legal_address_T_8 ;  
   wire _legal_address_T_9 ;  
   wire [39:0] _legal_address_T_10 ;  
   wire [40:0] _legal_address_T_11 ;  
   wire [40:0] _legal_address_T_13 ;  
   wire _legal_address_T_14 ;  
   wire [40:0] _legal_address_T_16 ;  
   wire [40:0] _legal_address_T_18 ;  
   wire _legal_address_T_19 ;  
   wire [39:0] _legal_address_T_20 ;  
   wire [40:0] _legal_address_T_21 ;  
   wire [40:0] _legal_address_T_23 ;  
   wire _legal_address_T_24 ;  
   wire [39:0] _legal_address_T_25 ;  
   wire [40:0] _legal_address_T_26 ;  
   wire [40:0] _legal_address_T_28 ;  
   wire _legal_address_T_29 ;  
   wire [39:0] _legal_address_T_30 ;  
   wire [40:0] _legal_address_T_31 ;  
   wire [40:0] _legal_address_T_33 ;  
   wire _legal_address_T_34 ;  
   wire _legal_address_T_35 ;  
   wire _legal_address_T_36 ;  
   wire _legal_address_T_37 ;  
   wire _legal_address_T_38 ;  
   wire _legal_address_T_39 ;  
   wire legal_address ;  
   wire [40:0] _cacheable_T_8 ;  
   wire _cacheable_T_9 ;  
   wire cacheable ;  
   wire [39:0] _homogeneous_T_54 ;  
   wire [40:0] _homogeneous_T_55 ;  
   wire [40:0] _homogeneous_T_57 ;  
   wire _homogeneous_T_58 ;  
   wire [40:0] _homogeneous_T_71 ;  
   wire _homogeneous_T_72 ;  
   wire _homogeneous_T_79 ;  
   wire _deny_access_to_debug_T ;  
   wire deny_access_to_debug ;  
   wire _prot_r_T_7 ;  
   wire prot_r ;  
   wire [39:0] _prot_w_T_10 ;  
   wire [40:0] _prot_w_T_11 ;  
   wire [40:0] _prot_w_T_13 ;  
   wire _prot_w_T_14 ;  
   wire [40:0] _prot_w_T_18 ;  
   wire _prot_w_T_19 ;  
   wire _prot_w_T_21 ;  
   wire _prot_w_T_22 ;  
   wire _prot_w_T_31 ;  
   wire _prot_w_T_33 ;  
   wire prot_w ;  
   wire prot_al ;  
   wire [40:0] _prot_x_T_3 ;  
   wire _prot_x_T_4 ;  
   wire _prot_x_T_15 ;  
   wire _prot_x_T_16 ;  
   wire _prot_x_T_31 ;  
   wire _prot_x_T_33 ;  
   wire prot_x ;  
   wire [40:0] _prot_eff_T_20 ;  
   wire _prot_eff_T_21 ;  
   wire [40:0] _prot_eff_T_25 ;  
   wire _prot_eff_T_26 ;  
   wire _prot_eff_T_37 ;  
   wire _prot_eff_T_38 ;  
   wire _prot_eff_T_39 ;  
   wire prot_eff ;  
   wire _sector_hits_T ;  
   wire _sector_hits_T_1 ;  
   wire _sector_hits_T_2 ;  
   wire [26:0] _sector_hits_T_3 ;  
   wire _sector_hits_T_5 ;  
   wire sector_hits_0 ;  
   wire _sector_hits_T_6 ;  
   wire _sector_hits_T_7 ;  
   wire _sector_hits_T_8 ;  
   wire [26:0] _sector_hits_T_9 ;  
   wire _sector_hits_T_11 ;  
   wire sector_hits_1 ;  
   wire _sector_hits_T_12 ;  
   wire _sector_hits_T_13 ;  
   wire _sector_hits_T_14 ;  
   wire [26:0] _sector_hits_T_15 ;  
   wire _sector_hits_T_17 ;  
   wire sector_hits_2 ;  
   wire _sector_hits_T_18 ;  
   wire _sector_hits_T_19 ;  
   wire _sector_hits_T_20 ;  
   wire [26:0] _sector_hits_T_21 ;  
   wire _sector_hits_T_23 ;  
   wire sector_hits_3 ;  
   wire _sector_hits_T_24 ;  
   wire _sector_hits_T_25 ;  
   wire _sector_hits_T_26 ;  
   wire [26:0] _sector_hits_T_27 ;  
   wire _sector_hits_T_29 ;  
   wire sector_hits_4 ;  
   wire _sector_hits_T_30 ;  
   wire _sector_hits_T_31 ;  
   wire _sector_hits_T_32 ;  
   wire [26:0] _sector_hits_T_33 ;  
   wire _sector_hits_T_35 ;  
   wire sector_hits_5 ;  
   wire _sector_hits_T_36 ;  
   wire _sector_hits_T_37 ;  
   wire _sector_hits_T_38 ;  
   wire [26:0] _sector_hits_T_39 ;  
   wire _sector_hits_T_41 ;  
   wire sector_hits_6 ;  
   wire _sector_hits_T_42 ;  
   wire _sector_hits_T_43 ;  
   wire _sector_hits_T_44 ;  
   wire [26:0] _sector_hits_T_45 ;  
   wire _sector_hits_T_47 ;  
   wire sector_hits_7 ;  
   wire _superpage_hits_T_2 ;  
   wire _superpage_hits_T_4 ;  
   wire superpage_hits_ignore_1 ;  
   wire _superpage_hits_T_7 ;  
   wire _superpage_hits_T_8 ;  
   wire superpage_hits_0 ;  
   wire _superpage_hits_T_16 ;  
   wire _superpage_hits_T_18 ;  
   wire superpage_hits_ignore_4 ;  
   wire _superpage_hits_T_21 ;  
   wire _superpage_hits_T_22 ;  
   wire superpage_hits_1 ;  
   wire _superpage_hits_T_30 ;  
   wire _superpage_hits_T_32 ;  
   wire superpage_hits_ignore_7 ;  
   wire _superpage_hits_T_35 ;  
   wire _superpage_hits_T_36 ;  
   wire superpage_hits_2 ;  
   wire _superpage_hits_T_44 ;  
   wire _superpage_hits_T_46 ;  
   wire superpage_hits_ignore_10 ;  
   wire _superpage_hits_T_49 ;  
   wire _superpage_hits_T_50 ;  
   wire superpage_hits_3 ;  
   wire [1:0] hitsVec_idx ;  
   wire _GEN_1 ;  
   wire _GEN_2 ;  
   wire _GEN_3 ;  
   wire _hitsVec_T_3 ;  
   wire hitsVec_0 ;  
   wire _GEN_5 ;  
   wire _GEN_6 ;  
   wire _GEN_7 ;  
   wire _hitsVec_T_7 ;  
   wire hitsVec_1 ;  
   wire _GEN_9 ;  
   wire _GEN_10 ;  
   wire _GEN_11 ;  
   wire _hitsVec_T_11 ;  
   wire hitsVec_2 ;  
   wire _GEN_13 ;  
   wire _GEN_14 ;  
   wire _GEN_15 ;  
   wire _hitsVec_T_15 ;  
   wire hitsVec_3 ;  
   wire _GEN_17 ;  
   wire _GEN_18 ;  
   wire _GEN_19 ;  
   wire _hitsVec_T_19 ;  
   wire hitsVec_4 ;  
   wire _GEN_21 ;  
   wire _GEN_22 ;  
   wire _GEN_23 ;  
   wire _hitsVec_T_23 ;  
   wire hitsVec_5 ;  
   wire _GEN_25 ;  
   wire _GEN_26 ;  
   wire _GEN_27 ;  
   wire _hitsVec_T_27 ;  
   wire hitsVec_6 ;  
   wire _GEN_29 ;  
   wire _GEN_30 ;  
   wire _GEN_31 ;  
   wire _hitsVec_T_31 ;  
   wire hitsVec_7 ;  
   wire hitsVec_8 ;  
   wire hitsVec_9 ;  
   wire hitsVec_10 ;  
   wire hitsVec_11 ;  
   wire _hitsVec_T_94 ;  
   wire _hitsVec_T_96 ;  
   wire _hitsVec_T_99 ;  
   wire _hitsVec_T_100 ;  
   wire _hitsVec_T_101 ;  
   wire _hitsVec_T_104 ;  
   wire _hitsVec_T_105 ;  
   wire _hitsVec_T_106 ;  
   wire hitsVec_12 ;  
   wire [5:0] real_hits_lo ;  
   wire [12:0] real_hits ;  
   wire hits_hi ;  
   wire [13:0] hits ;  
   wire newEntry_g ;  
   wire _newEntry_sr_T_1 ;  
   wire _newEntry_sr_T_2 ;  
   wire _newEntry_sr_T_3 ;  
   wire _newEntry_sr_T_4 ;  
   wire newEntry_sr ;  
   wire _newEntry_sw_T_5 ;  
   wire newEntry_sw ;  
   wire newEntry_sx ;  
   wire [7:0] special_entry_data_0_lo ;  
   wire [34:0] _special_entry_data_0_T ;  
   wire _GEN_32 ;  
   wire _T_2 ;  
   wire _T_3 ;  
   wire _GEN_35 ;  
   wire _T_4 ;  
   wire _GEN_39 ;  
   wire _T_5 ;  
   wire _GEN_43 ;  
   wire _T_6 ;  
   wire _GEN_47 ;  
   wire [2:0] waddr ;  
   wire _T_7 ;  
   wire _GEN_49 ;  
   wire _GEN_50 ;  
   wire _GEN_51 ;  
   wire _GEN_52 ;  
   wire [1:0] idx ;  
   wire _GEN_921 ;  
   wire _GEN_53 ;  
   wire _GEN_922 ;  
   wire _GEN_54 ;  
   wire _GEN_923 ;  
   wire _GEN_55 ;  
   wire _GEN_924 ;  
   wire _GEN_56 ;  
   wire _GEN_61 ;  
   wire _GEN_62 ;  
   wire _GEN_63 ;  
   wire _GEN_64 ;  
   wire _GEN_65 ;  
   wire _GEN_66 ;  
   wire _GEN_67 ;  
   wire _GEN_68 ;  
   wire _T_9 ;  
   wire _GEN_75 ;  
   wire _GEN_76 ;  
   wire _GEN_77 ;  
   wire _GEN_78 ;  
   wire _GEN_79 ;  
   wire _GEN_80 ;  
   wire _GEN_81 ;  
   wire _GEN_82 ;  
   wire _GEN_87 ;  
   wire _GEN_88 ;  
   wire _GEN_89 ;  
   wire _GEN_90 ;  
   wire _GEN_91 ;  
   wire _GEN_92 ;  
   wire _GEN_93 ;  
   wire _GEN_94 ;  
   wire _T_11 ;  
   wire _GEN_101 ;  
   wire _GEN_102 ;  
   wire _GEN_103 ;  
   wire _GEN_104 ;  
   wire _GEN_105 ;  
   wire _GEN_106 ;  
   wire _GEN_107 ;  
   wire _GEN_108 ;  
   wire _GEN_113 ;  
   wire _GEN_114 ;  
   wire _GEN_115 ;  
   wire _GEN_116 ;  
   wire _GEN_117 ;  
   wire _GEN_118 ;  
   wire _GEN_119 ;  
   wire _GEN_120 ;  
   wire _T_13 ;  
   wire _GEN_127 ;  
   wire _GEN_128 ;  
   wire _GEN_129 ;  
   wire _GEN_130 ;  
   wire _GEN_131 ;  
   wire _GEN_132 ;  
   wire _GEN_133 ;  
   wire _GEN_134 ;  
   wire _GEN_139 ;  
   wire _GEN_140 ;  
   wire _GEN_141 ;  
   wire _GEN_142 ;  
   wire _GEN_143 ;  
   wire _GEN_144 ;  
   wire _GEN_145 ;  
   wire _GEN_146 ;  
   wire _T_15 ;  
   wire _GEN_153 ;  
   wire _GEN_154 ;  
   wire _GEN_155 ;  
   wire _GEN_156 ;  
   wire _GEN_157 ;  
   wire _GEN_158 ;  
   wire _GEN_159 ;  
   wire _GEN_160 ;  
   wire _GEN_165 ;  
   wire _GEN_166 ;  
   wire _GEN_167 ;  
   wire _GEN_168 ;  
   wire _GEN_169 ;  
   wire _GEN_170 ;  
   wire _GEN_171 ;  
   wire _GEN_172 ;  
   wire _T_17 ;  
   wire _GEN_179 ;  
   wire _GEN_180 ;  
   wire _GEN_181 ;  
   wire _GEN_182 ;  
   wire _GEN_183 ;  
   wire _GEN_184 ;  
   wire _GEN_185 ;  
   wire _GEN_186 ;  
   wire _GEN_191 ;  
   wire _GEN_192 ;  
   wire _GEN_193 ;  
   wire _GEN_194 ;  
   wire _GEN_195 ;  
   wire _GEN_196 ;  
   wire _GEN_197 ;  
   wire _GEN_198 ;  
   wire _T_19 ;  
   wire _GEN_205 ;  
   wire _GEN_206 ;  
   wire _GEN_207 ;  
   wire _GEN_208 ;  
   wire _GEN_209 ;  
   wire _GEN_210 ;  
   wire _GEN_211 ;  
   wire _GEN_212 ;  
   wire _GEN_217 ;  
   wire _GEN_218 ;  
   wire _GEN_219 ;  
   wire _GEN_220 ;  
   wire _GEN_221 ;  
   wire _GEN_222 ;  
   wire _GEN_223 ;  
   wire _GEN_224 ;  
   wire _T_21 ;  
   wire _GEN_231 ;  
   wire _GEN_232 ;  
   wire _GEN_233 ;  
   wire _GEN_234 ;  
   wire _GEN_235 ;  
   wire _GEN_236 ;  
   wire _GEN_237 ;  
   wire _GEN_238 ;  
   wire _GEN_243 ;  
   wire _GEN_244 ;  
   wire _GEN_245 ;  
   wire _GEN_246 ;  
   wire _GEN_247 ;  
   wire _GEN_248 ;  
   wire _GEN_249 ;  
   wire _GEN_250 ;  
   wire _GEN_259 ;  
   wire _GEN_263 ;  
   wire _GEN_267 ;  
   wire _GEN_271 ;  
   wire _GEN_273 ;  
   wire _GEN_274 ;  
   wire _GEN_275 ;  
   wire _GEN_276 ;  
   wire _GEN_283 ;  
   wire _GEN_284 ;  
   wire _GEN_285 ;  
   wire _GEN_286 ;  
   wire _GEN_293 ;  
   wire _GEN_294 ;  
   wire _GEN_295 ;  
   wire _GEN_296 ;  
   wire _GEN_303 ;  
   wire _GEN_304 ;  
   wire _GEN_305 ;  
   wire _GEN_306 ;  
   wire _GEN_313 ;  
   wire _GEN_314 ;  
   wire _GEN_315 ;  
   wire _GEN_316 ;  
   wire _GEN_323 ;  
   wire _GEN_324 ;  
   wire _GEN_325 ;  
   wire _GEN_326 ;  
   wire _GEN_333 ;  
   wire _GEN_334 ;  
   wire _GEN_335 ;  
   wire _GEN_336 ;  
   wire _GEN_343 ;  
   wire _GEN_344 ;  
   wire _GEN_345 ;  
   wire _GEN_346 ;  
   wire _GEN_355 ;  
   wire _GEN_359 ;  
   wire _GEN_363 ;  
   wire _GEN_367 ;  
   wire _GEN_371 ;  
   wire _GEN_373 ;  
   wire _GEN_374 ;  
   wire _GEN_375 ;  
   wire _GEN_376 ;  
   wire _GEN_383 ;  
   wire _GEN_384 ;  
   wire _GEN_385 ;  
   wire _GEN_386 ;  
   wire _GEN_393 ;  
   wire _GEN_394 ;  
   wire _GEN_395 ;  
   wire _GEN_396 ;  
   wire _GEN_403 ;  
   wire _GEN_404 ;  
   wire _GEN_405 ;  
   wire _GEN_406 ;  
   wire _GEN_413 ;  
   wire _GEN_414 ;  
   wire _GEN_415 ;  
   wire _GEN_416 ;  
   wire _GEN_423 ;  
   wire _GEN_424 ;  
   wire _GEN_425 ;  
   wire _GEN_426 ;  
   wire _GEN_433 ;  
   wire _GEN_434 ;  
   wire _GEN_435 ;  
   wire _GEN_436 ;  
   wire _GEN_443 ;  
   wire _GEN_444 ;  
   wire _GEN_445 ;  
   wire _GEN_446 ;  
   wire _GEN_455 ;  
   wire _GEN_459 ;  
   wire _GEN_463 ;  
   wire _GEN_467 ;  
   wire _GEN_471 ;  
   wire _GEN_473 ;  
   wire _GEN_474 ;  
   wire _GEN_475 ;  
   wire _GEN_476 ;  
   wire _GEN_483 ;  
   wire _GEN_484 ;  
   wire _GEN_485 ;  
   wire _GEN_486 ;  
   wire _GEN_493 ;  
   wire _GEN_494 ;  
   wire _GEN_495 ;  
   wire _GEN_496 ;  
   wire _GEN_503 ;  
   wire _GEN_504 ;  
   wire _GEN_505 ;  
   wire _GEN_506 ;  
   wire _GEN_513 ;  
   wire _GEN_514 ;  
   wire _GEN_515 ;  
   wire _GEN_516 ;  
   wire _GEN_523 ;  
   wire _GEN_524 ;  
   wire _GEN_525 ;  
   wire _GEN_526 ;  
   wire _GEN_533 ;  
   wire _GEN_534 ;  
   wire _GEN_535 ;  
   wire _GEN_536 ;  
   wire _GEN_543 ;  
   wire _GEN_544 ;  
   wire _GEN_545 ;  
   wire _GEN_546 ;  
   wire [34:0] _GEN_554 ;  
   wire [34:0] _GEN_555 ;  
   wire [34:0] _GEN_556 ;  
   wire [34:0] _GEN_558 ;  
   wire [34:0] _GEN_559 ;  
   wire [34:0] _GEN_560 ;  
   wire [34:0] _GEN_562 ;  
   wire [34:0] _GEN_563 ;  
   wire [34:0] _GEN_564 ;  
   wire [34:0] _GEN_566 ;  
   wire [34:0] _GEN_567 ;  
   wire [34:0] _GEN_568 ;  
   wire [34:0] _GEN_570 ;  
   wire [34:0] _GEN_571 ;  
   wire [34:0] _GEN_572 ;  
   wire [34:0] _GEN_574 ;  
   wire [34:0] _GEN_575 ;  
   wire [34:0] _GEN_576 ;  
   wire [34:0] _GEN_578 ;  
   wire [34:0] _GEN_579 ;  
   wire [34:0] _GEN_580 ;  
   wire [34:0] _GEN_582 ;  
   wire [34:0] _GEN_583 ;  
   wire [34:0] _GEN_584 ;  
   wire [1:0] ppn_hi ;  
   wire [26:0] _ppn_T_1 ;  
   wire [26:0] _GEN_953 ;  
   wire [26:0] _ppn_T_2 ;  
   wire [8:0] ppn_lo ;  
   wire [26:0] _ppn_T_4 ;  
   wire [8:0] ppn_lo_1 ;  
   wire [19:0] _ppn_T_5 ;  
   wire [1:0] ppn_hi_2 ;  
   wire [26:0] _ppn_T_6 ;  
   wire [26:0] _GEN_955 ;  
   wire [26:0] _ppn_T_7 ;  
   wire [8:0] ppn_lo_2 ;  
   wire [26:0] _ppn_T_9 ;  
   wire [8:0] ppn_lo_3 ;  
   wire [19:0] _ppn_T_10 ;  
   wire [1:0] ppn_hi_4 ;  
   wire [26:0] _ppn_T_11 ;  
   wire [26:0] _GEN_957 ;  
   wire [26:0] _ppn_T_12 ;  
   wire [8:0] ppn_lo_4 ;  
   wire [26:0] _ppn_T_14 ;  
   wire [8:0] ppn_lo_5 ;  
   wire [19:0] _ppn_T_15 ;  
   wire [1:0] ppn_hi_6 ;  
   wire [26:0] _ppn_T_16 ;  
   wire [26:0] _GEN_959 ;  
   wire [26:0] _ppn_T_17 ;  
   wire [8:0] ppn_lo_6 ;  
   wire [26:0] _ppn_T_19 ;  
   wire [8:0] ppn_lo_7 ;  
   wire [19:0] _ppn_T_20 ;  
   wire [1:0] ppn_hi_8 ;  
   wire [26:0] _GEN_961 ;  
   wire [26:0] _ppn_T_22 ;  
   wire [8:0] ppn_lo_8 ;  
   wire [26:0] _ppn_T_24 ;  
   wire [8:0] ppn_lo_9 ;  
   wire [19:0] _ppn_T_25 ;  
   wire [19:0] _ppn_T_27 ;  
   wire [19:0] _ppn_T_28 ;  
   wire [19:0] _ppn_T_29 ;  
   wire [19:0] _ppn_T_30 ;  
   wire [19:0] _ppn_T_31 ;  
   wire [19:0] _ppn_T_32 ;  
   wire [19:0] _ppn_T_33 ;  
   wire [19:0] _ppn_T_34 ;  
   wire [19:0] _ppn_T_35 ;  
   wire [19:0] _ppn_T_36 ;  
   wire [19:0] _ppn_T_37 ;  
   wire [19:0] _ppn_T_38 ;  
   wire [19:0] _ppn_T_39 ;  
   wire [19:0] _ppn_T_40 ;  
   wire [19:0] _ppn_T_41 ;  
   wire [19:0] _ppn_T_42 ;  
   wire [19:0] _ppn_T_43 ;  
   wire [19:0] _ppn_T_44 ;  
   wire [19:0] _ppn_T_45 ;  
   wire [19:0] _ppn_T_46 ;  
   wire [19:0] _ppn_T_47 ;  
   wire [19:0] _ppn_T_48 ;  
   wire [19:0] _ppn_T_49 ;  
   wire [19:0] _ppn_T_50 ;  
   wire [19:0] _ppn_T_51 ;  
   wire [19:0] _ppn_T_52 ;  
   wire [19:0] ppn ;  
   wire [5:0] ptw_ae_array_lo ;  
   wire [13:0] ptw_ae_array ;  
   wire [5:0] priv_rw_ok_lo ;  
   wire [12:0] _priv_rw_ok_T_2 ;  
   wire [12:0] priv_x_ok ;  
   wire [5:0] r_array_lo_1 ;  
   wire [12:0] _r_array_T_1 ;  
   wire [12:0] x_array_lo_1 ;  
   wire [13:0] x_array ;  
   wire [1:0] px_array_hi ;  
   wire [5:0] px_array_lo ;  
   wire [13:0] _px_array_T_1 ;  
   wire [13:0] px_array ;  
   wire [1:0] c_array_hi ;  
   wire [5:0] c_array_lo ;  
   wire [13:0] c_array ;  
   wire [39:0] bad_va_maskedVAddr ;  
   wire _bad_va_T_1 ;  
   wire _bad_va_T_2 ;  
   wire _bad_va_T_3 ;  
   wire bad_va ;  
   wire [13:0] _pf_inst_array_T ;  
   wire [13:0] pf_inst_array ;  
   wire tlb_hit ;  
   wire _tlb_miss_T_1 ;  
   wire tlb_miss ;  
   reg [6:0] state_vec_0 ;  
   reg [31:0] _RAND_98 ;  
   reg [2:0] state_reg_1 ;  
   reg [31:0] _RAND_99 ;  
   wire _T_23 ;  
   wire _T_24 ;  
   wire _T_25 ;  
   wire _T_26 ;  
   wire _T_27 ;  
   wire _T_28 ;  
   wire _T_29 ;  
   wire _T_30 ;  
   wire [7:0] _T_31 ;  
   wire [3:0] hi_1 ;  
   wire [3:0] lo_1 ;  
   wire hi_2 ;  
   wire [3:0] _T_32 ;  
   wire [1:0] hi_3 ;  
   wire [1:0] lo_2 ;  
   wire hi_4 ;  
   wire [1:0] _T_33 ;  
   wire lo_3 ;  
   wire [2:0] state_vec_0_touch_way_sized ;  
   wire state_vec_0_hi_hi ;  
   wire [2:0] state_vec_0_left_subtree_state ;  
   wire [2:0] state_vec_0_right_subtree_state ;  
   wire state_vec_0_hi_hi_1 ;  
   wire state_vec_0_left_subtree_state_1 ;  
   wire state_vec_0_right_subtree_state_1 ;  
   wire state_vec_0_hi_lo ;  
   wire state_vec_0_lo ;  
   wire [2:0] _state_vec_0_T_7 ;  
   wire [2:0] state_vec_0_hi_lo_1 ;  
   wire state_vec_0_left_subtree_state_2 ;  
   wire state_vec_0_right_subtree_state_2 ;  
   wire state_vec_0_hi_lo_2 ;  
   wire state_vec_0_lo_1 ;  
   wire [2:0] _state_vec_0_T_15 ;  
   wire [2:0] state_vec_0_lo_2 ;  
   wire [6:0] _state_vec_0_T_16 ;  
   wire _T_35 ;  
   wire _T_36 ;  
   wire _T_37 ;  
   wire [3:0] _T_38 ;  
   wire [1:0] hi_6 ;  
   wire [1:0] lo_6 ;  
   wire hi_7 ;  
   wire [1:0] _T_39 ;  
   wire lo_7 ;  
   wire [1:0] state_reg_touch_way_sized ;  
   wire state_reg_hi_hi ;  
   wire state_reg_left_subtree_state ;  
   wire state_reg_right_subtree_state ;  
   wire state_reg_hi_lo ;  
   wire state_reg_lo ;  
   wire [2:0] _state_reg_T_6 ;  
   wire multipleHits_leftOne ;  
   wire multipleHits_leftOne_1 ;  
   wire multipleHits_rightOne ;  
   wire multipleHits_rightOne_1 ;  
   wire multipleHits_rightTwo ;  
   wire multipleHits_leftOne_2 ;  
   wire _multipleHits_T_9 ;  
   wire multipleHits_leftTwo ;  
   wire multipleHits_leftOne_3 ;  
   wire multipleHits_leftOne_4 ;  
   wire multipleHits_rightOne_2 ;  
   wire multipleHits_rightOne_3 ;  
   wire multipleHits_rightTwo_1 ;  
   wire multipleHits_rightOne_4 ;  
   wire _multipleHits_T_18 ;  
   wire multipleHits_rightTwo_2 ;  
   wire multipleHits_leftOne_5 ;  
   wire _multipleHits_T_19 ;  
   wire _multipleHits_T_20 ;  
   wire multipleHits_leftTwo_1 ;  
   wire multipleHits_leftOne_6 ;  
   wire multipleHits_leftOne_7 ;  
   wire multipleHits_rightOne_5 ;  
   wire multipleHits_rightOne_6 ;  
   wire multipleHits_rightTwo_3 ;  
   wire multipleHits_leftOne_8 ;  
   wire _multipleHits_T_30 ;  
   wire multipleHits_leftTwo_2 ;  
   wire multipleHits_leftOne_9 ;  
   wire multipleHits_rightOne_7 ;  
   wire multipleHits_leftOne_10 ;  
   wire multipleHits_leftTwo_3 ;  
   wire multipleHits_leftOne_11 ;  
   wire multipleHits_rightOne_8 ;  
   wire multipleHits_rightOne_9 ;  
   wire multipleHits_rightTwo_4 ;  
   wire multipleHits_rightOne_10 ;  
   wire _multipleHits_T_42 ;  
   wire _multipleHits_T_43 ;  
   wire multipleHits_rightTwo_5 ;  
   wire multipleHits_rightOne_11 ;  
   wire _multipleHits_T_44 ;  
   wire _multipleHits_T_45 ;  
   wire multipleHits_rightTwo_6 ;  
   wire _multipleHits_T_47 ;  
   wire _multipleHits_T_48 ;  
   wire multipleHits ;  
   wire [13:0] _io_resp_pf_inst_T ;  
   wire _io_resp_pf_inst_T_1 ;  
   wire [13:0] _io_resp_ae_inst_T_1 ;  
   wire [13:0] _io_resp_cacheable_T ;  
   wire _io_resp_miss_T ;  
   wire _T_41 ;  
   wire _T_42 ;  
   wire r_superpage_repl_addr_hi ;  
   wire r_superpage_repl_addr_lo ;  
   wire [1:0] _r_superpage_repl_addr_T_2 ;  
   wire [3:0] r_superpage_repl_addr_valids ;  
   wire _r_superpage_repl_addr_T_3 ;  
   wire _r_superpage_repl_addr_T_5 ;  
   wire _r_superpage_repl_addr_T_6 ;  
   wire _r_superpage_repl_addr_T_7 ;  
   wire r_sectored_repl_addr_hi ;  
   wire r_sectored_repl_addr_hi_1 ;  
   wire r_sectored_repl_addr_lo ;  
   wire [1:0] _r_sectored_repl_addr_T_2 ;  
   wire r_sectored_repl_addr_hi_2 ;  
   wire r_sectored_repl_addr_lo_1 ;  
   wire [1:0] _r_sectored_repl_addr_T_5 ;  
   wire [1:0] r_sectored_repl_addr_lo_2 ;  
   wire [2:0] _r_sectored_repl_addr_T_6 ;  
   wire [7:0] r_sectored_repl_addr_valids ;  
   wire _r_sectored_repl_addr_T_7 ;  
   wire _r_sectored_repl_addr_T_9 ;  
   wire _r_sectored_repl_addr_T_10 ;  
   wire _r_sectored_repl_addr_T_11 ;  
   wire _r_sectored_repl_addr_T_12 ;  
   wire _r_sectored_repl_addr_T_13 ;  
   wire _r_sectored_repl_addr_T_14 ;  
   wire _r_sectored_repl_addr_T_15 ;  
   wire _T_44 ;  
   wire _T_45 ;  
   wire _T_48 ;  
   wire _T_49 ;  
   wire _T_51 ;  
   wire _T_59 ;  
   wire _GEN_617 ;  
   wire _GEN_618 ;  
   wire _GEN_619 ;  
   wire _GEN_620 ;  
   wire _GEN_621 ;  
   wire _GEN_622 ;  
   wire _GEN_623 ;  
   wire _GEN_624 ;  
   wire _T_198 ;  
   wire _GEN_645 ;  
   wire _GEN_646 ;  
   wire _GEN_647 ;  
   wire _GEN_648 ;  
   wire _GEN_649 ;  
   wire _GEN_650 ;  
   wire _GEN_651 ;  
   wire _GEN_652 ;  
   wire _T_337 ;  
   wire _GEN_673 ;  
   wire _GEN_674 ;  
   wire _GEN_675 ;  
   wire _GEN_676 ;  
   wire _GEN_677 ;  
   wire _GEN_678 ;  
   wire _GEN_679 ;  
   wire _GEN_680 ;  
   wire _T_476 ;  
   wire _GEN_701 ;  
   wire _GEN_702 ;  
   wire _GEN_703 ;  
   wire _GEN_704 ;  
   wire _GEN_705 ;  
   wire _GEN_706 ;  
   wire _GEN_707 ;  
   wire _GEN_708 ;  
   wire _T_615 ;  
   wire _GEN_729 ;  
   wire _GEN_730 ;  
   wire _GEN_731 ;  
   wire _GEN_732 ;  
   wire _GEN_733 ;  
   wire _GEN_734 ;  
   wire _GEN_735 ;  
   wire _GEN_736 ;  
   wire _T_754 ;  
   wire _GEN_757 ;  
   wire _GEN_758 ;  
   wire _GEN_759 ;  
   wire _GEN_760 ;  
   wire _GEN_761 ;  
   wire _GEN_762 ;  
   wire _GEN_763 ;  
   wire _GEN_764 ;  
   wire _T_893 ;  
   wire _GEN_785 ;  
   wire _GEN_786 ;  
   wire _GEN_787 ;  
   wire _GEN_788 ;  
   wire _GEN_789 ;  
   wire _GEN_790 ;  
   wire _GEN_791 ;  
   wire _GEN_792 ;  
   wire _T_1032 ;  
   wire _GEN_813 ;  
   wire _GEN_814 ;  
   wire _GEN_815 ;  
   wire _GEN_816 ;  
   wire _GEN_817 ;  
   wire _GEN_818 ;  
   wire _GEN_819 ;  
   wire _GEN_820 ;  
   wire _GEN_826 ;  
   wire _GEN_827 ;  
   wire _GEN_830 ;  
   wire _GEN_831 ;  
   wire _GEN_834 ;  
   wire _GEN_835 ;  
   wire _GEN_838 ;  
   wire _GEN_839 ;  
   wire _GEN_842 ;  
   wire _GEN_843 ;  
   wire _T_1326 ;  
   reg [19:0] TLB_1_state ;  
   reg [31:0] _RAND_100 ;  
   reg TLB_1_cov[0:1048575] ;  
   reg [31:0] _RAND_101 ;  
   wire TLB_1_cov_read_data ;  
   wire [19:0] TLB_1_cov_read_addr ;  
   wire TLB_1_cov_write_data ;  
   wire [19:0] TLB_1_cov_write_addr ;  
   wire TLB_1_cov_write_mask ;  
   wire TLB_1_cov_write_en ;  
   reg [29:0] TLB_1_covSum ;  
   reg [31:0] _RAND_102 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire mux_cond_4 ;  
   wire mux_cond_5 ;  
   wire mux_cond_6 ;  
   wire mux_cond_7 ;  
   wire mux_cond_8 ;  
   wire mux_cond_9 ;  
   wire mux_cond_10 ;  
   wire mux_cond_11 ;  
   wire mux_cond_12 ;  
   wire mux_cond_13 ;  
   wire mux_cond_14 ;  
   wire mux_cond_15 ;  
   wire mux_cond_16 ;  
   wire mux_cond_17 ;  
   wire mux_cond_18 ;  
   wire mux_cond_19 ;  
   wire mux_cond_20 ;  
   wire mux_cond_21 ;  
   wire mux_cond_22 ;  
   wire mux_cond_23 ;  
   wire mux_cond_24 ;  
   wire mux_cond_25 ;  
   wire mux_cond_26 ;  
   wire mux_cond_27 ;  
   wire mux_cond_28 ;  
   wire mux_cond_29 ;  
   wire mux_cond_30 ;  
   wire mux_cond_31 ;  
   wire mux_cond_32 ;  
   wire mux_cond_33 ;  
   wire mux_cond_34 ;  
   wire mux_cond_35 ;  
   wire mux_cond_36 ;  
   wire mux_cond_37 ;  
   wire mux_cond_38 ;  
   wire mux_cond_39 ;  
   wire mux_cond_40 ;  
   wire mux_cond_41 ;  
   wire mux_cond_42 ;  
   wire mux_cond_43 ;  
   wire mux_cond_44 ;  
   wire mux_cond_45 ;  
   wire mux_cond_46 ;  
   wire mux_cond_47 ;  
   wire mux_cond_48 ;  
   wire mux_cond_49 ;  
   wire mux_cond_50 ;  
   wire mux_cond_51 ;  
   wire mux_cond_52 ;  
   wire mux_cond_53 ;  
   wire mux_cond_54 ;  
   wire mux_cond_55 ;  
   wire mux_cond_56 ;  
   wire mux_cond_57 ;  
   wire mux_cond_58 ;  
   wire mux_cond_59 ;  
   wire mux_cond_60 ;  
   wire mux_cond_61 ;  
   wire mux_cond_62 ;  
   wire mux_cond_63 ;  
   wire mux_cond_64 ;  
   wire mux_cond_65 ;  
   wire mux_cond_66 ;  
   wire mux_cond_67 ;  
   wire mux_cond_68 ;  
   wire r_sectored_hit_shl ;  
   wire [19:0] r_sectored_hit_pad ;  
   wire [10:0] r_sectored_repl_addr_shl ;  
   wire [19:0] r_sectored_repl_addr_pad ;  
   wire [1:0] r_superpage_repl_addr_shl ;  
   wire [19:0] r_superpage_repl_addr_pad ;  
   wire [13:0] special_entry_valid_0_shl ;  
   wire [19:0] special_entry_valid_0_pad ;  
   wire [13:0] special_entry_level_shl ;  
   wire [19:0] special_entry_level_pad ;  
   wire [13:0] state_shl ;  
   wire [19:0] state_pad ;  
   wire [3:0] r_sectored_hit_addr_shl ;  
   wire [19:0] r_sectored_hit_addr_pad ;  
   wire [16:0] mux_cond_0_shl ;  
   wire [19:0] mux_cond_0_pad ;  
   wire [10:0] mux_cond_1_shl ;  
   wire [19:0] mux_cond_1_pad ;  
   wire [2:0] mux_cond_2_shl ;  
   wire [19:0] mux_cond_2_pad ;  
   wire [15:0] mux_cond_3_shl ;  
   wire [19:0] mux_cond_3_pad ;  
   wire [4:0] mux_cond_4_shl ;  
   wire [19:0] mux_cond_4_pad ;  
   wire [13:0] mux_cond_5_shl ;  
   wire [19:0] mux_cond_5_pad ;  
   wire [9:0] mux_cond_6_shl ;  
   wire [19:0] mux_cond_6_pad ;  
   wire [8:0] mux_cond_7_shl ;  
   wire [19:0] mux_cond_7_pad ;  
   wire [12:0] mux_cond_8_shl ;  
   wire [19:0] mux_cond_8_pad ;  
   wire [19:0] mux_cond_9_shl ;  
   wire [19:0] mux_cond_9_pad ;  
   wire [18:0] mux_cond_10_shl ;  
   wire [19:0] mux_cond_10_pad ;  
   wire [9:0] mux_cond_11_shl ;  
   wire [19:0] mux_cond_11_pad ;  
   wire [19:0] mux_cond_12_shl ;  
   wire [19:0] mux_cond_12_pad ;  
   wire [7:0] mux_cond_13_shl ;  
   wire [19:0] mux_cond_13_pad ;  
   wire [11:0] mux_cond_14_shl ;  
   wire [19:0] mux_cond_14_pad ;  
   wire mux_cond_15_shl ;  
   wire [19:0] mux_cond_15_pad ;  
   wire [4:0] mux_cond_16_shl ;  
   wire [19:0] mux_cond_16_pad ;  
   wire [19:0] mux_cond_17_shl ;  
   wire [19:0] mux_cond_17_pad ;  
   wire [9:0] mux_cond_18_shl ;  
   wire [19:0] mux_cond_18_pad ;  
   wire [8:0] mux_cond_19_shl ;  
   wire [19:0] mux_cond_19_pad ;  
   wire [4:0] mux_cond_20_shl ;  
   wire [19:0] mux_cond_20_pad ;  
   wire [6:0] mux_cond_21_shl ;  
   wire [19:0] mux_cond_21_pad ;  
   wire [11:0] mux_cond_22_shl ;  
   wire [19:0] mux_cond_22_pad ;  
   wire [14:0] mux_cond_23_shl ;  
   wire [19:0] mux_cond_23_pad ;  
   wire [7:0] mux_cond_24_shl ;  
   wire [19:0] mux_cond_24_pad ;  
   wire [7:0] mux_cond_25_shl ;  
   wire [19:0] mux_cond_25_pad ;  
   wire [19:0] mux_cond_26_shl ;  
   wire [19:0] mux_cond_26_pad ;  
   wire [10:0] mux_cond_27_shl ;  
   wire [19:0] mux_cond_27_pad ;  
   wire [17:0] mux_cond_28_shl ;  
   wire [19:0] mux_cond_28_pad ;  
   wire [3:0] mux_cond_29_shl ;  
   wire [19:0] mux_cond_29_pad ;  
   wire [9:0] mux_cond_30_shl ;  
   wire [19:0] mux_cond_30_pad ;  
   wire [15:0] mux_cond_31_shl ;  
   wire [19:0] mux_cond_31_pad ;  
   wire mux_cond_32_shl ;  
   wire [19:0] mux_cond_32_pad ;  
   wire [12:0] mux_cond_33_shl ;  
   wire [19:0] mux_cond_33_pad ;  
   wire [17:0] mux_cond_34_shl ;  
   wire [19:0] mux_cond_34_pad ;  
   wire [9:0] mux_cond_35_shl ;  
   wire [19:0] mux_cond_35_pad ;  
   wire [12:0] mux_cond_36_shl ;  
   wire [19:0] mux_cond_36_pad ;  
   wire mux_cond_37_shl ;  
   wire [19:0] mux_cond_37_pad ;  
   wire [5:0] mux_cond_38_shl ;  
   wire [19:0] mux_cond_38_pad ;  
   wire [2:0] mux_cond_39_shl ;  
   wire [19:0] mux_cond_39_pad ;  
   wire [18:0] mux_cond_40_shl ;  
   wire [19:0] mux_cond_40_pad ;  
   wire [13:0] mux_cond_41_shl ;  
   wire [19:0] mux_cond_41_pad ;  
   wire [5:0] mux_cond_42_shl ;  
   wire [19:0] mux_cond_42_pad ;  
   wire [18:0] mux_cond_43_shl ;  
   wire [19:0] mux_cond_43_pad ;  
   wire [18:0] mux_cond_44_shl ;  
   wire [19:0] mux_cond_44_pad ;  
   wire [2:0] mux_cond_45_shl ;  
   wire [19:0] mux_cond_45_pad ;  
   wire [12:0] mux_cond_46_shl ;  
   wire [19:0] mux_cond_46_pad ;  
   wire [18:0] mux_cond_47_shl ;  
   wire [19:0] mux_cond_47_pad ;  
   wire [16:0] mux_cond_48_shl ;  
   wire [19:0] mux_cond_48_pad ;  
   wire mux_cond_49_shl ;  
   wire [19:0] mux_cond_49_pad ;  
   wire [4:0] mux_cond_50_shl ;  
   wire [19:0] mux_cond_50_pad ;  
   wire [9:0] mux_cond_51_shl ;  
   wire [19:0] mux_cond_51_pad ;  
   wire [13:0] mux_cond_52_shl ;  
   wire [19:0] mux_cond_52_pad ;  
   wire [4:0] mux_cond_53_shl ;  
   wire [19:0] mux_cond_53_pad ;  
   wire [5:0] mux_cond_54_shl ;  
   wire [19:0] mux_cond_54_pad ;  
   wire [10:0] mux_cond_55_shl ;  
   wire [19:0] mux_cond_55_pad ;  
   wire [12:0] mux_cond_56_shl ;  
   wire [19:0] mux_cond_56_pad ;  
   wire [4:0] mux_cond_57_shl ;  
   wire [19:0] mux_cond_57_pad ;  
   wire [19:0] mux_cond_58_shl ;  
   wire [19:0] mux_cond_58_pad ;  
   wire [8:0] mux_cond_59_shl ;  
   wire [19:0] mux_cond_59_pad ;  
   wire [12:0] mux_cond_60_shl ;  
   wire [19:0] mux_cond_60_pad ;  
   wire [13:0] mux_cond_61_shl ;  
   wire [19:0] mux_cond_61_pad ;  
   wire [19:0] mux_cond_62_shl ;  
   wire [19:0] mux_cond_62_pad ;  
   wire [7:0] mux_cond_63_shl ;  
   wire [19:0] mux_cond_63_pad ;  
   wire [1:0] mux_cond_64_shl ;  
   wire [19:0] mux_cond_64_pad ;  
   wire [3:0] mux_cond_65_shl ;  
   wire [19:0] mux_cond_65_pad ;  
   wire [1:0] mux_cond_66_shl ;  
   wire [19:0] mux_cond_66_pad ;  
   wire [15:0] mux_cond_67_shl ;  
   wire [19:0] mux_cond_67_pad ;  
   wire [15:0] mux_cond_68_shl ;  
   wire [19:0] mux_cond_68_pad ;  
   wire [5:0] sectored_entries_0_0_valid_3_shl ;  
   wire [19:0] sectored_entries_0_0_valid_3_pad ;  
   wire [4:0] sectored_entries_0_0_valid_2_shl ;  
   wire [19:0] sectored_entries_0_0_valid_2_pad ;  
   wire [5:0] sectored_entries_0_2_valid_0_shl ;  
   wire [19:0] sectored_entries_0_2_valid_0_pad ;  
   wire [5:0] sectored_entries_0_3_valid_0_shl ;  
   wire [19:0] sectored_entries_0_3_valid_0_pad ;  
   wire [14:0] superpage_entries_2_level_shl ;  
   wire [19:0] superpage_entries_2_level_pad ;  
   wire [4:0] sectored_entries_0_7_valid_1_shl ;  
   wire [19:0] sectored_entries_0_7_valid_1_pad ;  
   wire [5:0] sectored_entries_0_4_valid_0_shl ;  
   wire [19:0] sectored_entries_0_4_valid_0_pad ;  
   wire [5:0] sectored_entries_0_1_valid_3_shl ;  
   wire [19:0] sectored_entries_0_1_valid_3_pad ;  
   wire [4:0] sectored_entries_0_1_valid_1_shl ;  
   wire [19:0] sectored_entries_0_1_valid_1_pad ;  
   wire [5:0] sectored_entries_0_2_valid_3_shl ;  
   wire [19:0] sectored_entries_0_2_valid_3_pad ;  
   wire [4:0] sectored_entries_0_2_valid_1_shl ;  
   wire [19:0] sectored_entries_0_2_valid_1_pad ;  
   wire [1:0] superpage_entries_1_valid_0_shl ;  
   wire [19:0] superpage_entries_1_valid_0_pad ;  
   wire [5:0] sectored_entries_0_7_valid_0_shl ;  
   wire [19:0] sectored_entries_0_7_valid_0_pad ;  
   wire [1:0] superpage_entries_3_valid_0_shl ;  
   wire [19:0] superpage_entries_3_valid_0_pad ;  
   wire [5:0] sectored_entries_0_5_valid_3_shl ;  
   wire [19:0] sectored_entries_0_5_valid_3_pad ;  
   wire [4:0] sectored_entries_0_5_valid_1_shl ;  
   wire [19:0] sectored_entries_0_5_valid_1_pad ;  
   wire [5:0] sectored_entries_0_4_valid_3_shl ;  
   wire [19:0] sectored_entries_0_4_valid_3_pad ;  
   wire [4:0] sectored_entries_0_5_valid_2_shl ;  
   wire [19:0] sectored_entries_0_5_valid_2_pad ;  
   wire [4:0] sectored_entries_0_1_valid_2_shl ;  
   wire [19:0] sectored_entries_0_1_valid_2_pad ;  
   wire [4:0] sectored_entries_0_3_valid_1_shl ;  
   wire [19:0] sectored_entries_0_3_valid_1_pad ;  
   wire [5:0] sectored_entries_0_1_valid_0_shl ;  
   wire [19:0] sectored_entries_0_1_valid_0_pad ;  
   wire [4:0] sectored_entries_0_4_valid_2_shl ;  
   wire [19:0] sectored_entries_0_4_valid_2_pad ;  
   wire [4:0] sectored_entries_0_4_valid_1_shl ;  
   wire [19:0] sectored_entries_0_4_valid_1_pad ;  
   wire [14:0] superpage_entries_3_level_shl ;  
   wire [19:0] superpage_entries_3_level_pad ;  
   wire [4:0] sectored_entries_0_0_valid_1_shl ;  
   wire [19:0] sectored_entries_0_0_valid_1_pad ;  
   wire [4:0] sectored_entries_0_3_valid_2_shl ;  
   wire [19:0] sectored_entries_0_3_valid_2_pad ;  
   wire [4:0] sectored_entries_0_6_valid_1_shl ;  
   wire [19:0] sectored_entries_0_6_valid_1_pad ;  
   wire [5:0] sectored_entries_0_7_valid_3_shl ;  
   wire [19:0] sectored_entries_0_7_valid_3_pad ;  
   wire [5:0] sectored_entries_0_3_valid_3_shl ;  
   wire [19:0] sectored_entries_0_3_valid_3_pad ;  
   wire [5:0] sectored_entries_0_0_valid_0_shl ;  
   wire [19:0] sectored_entries_0_0_valid_0_pad ;  
   wire [1:0] superpage_entries_0_valid_0_shl ;  
   wire [19:0] superpage_entries_0_valid_0_pad ;  
   wire [4:0] sectored_entries_0_2_valid_2_shl ;  
   wire [19:0] sectored_entries_0_2_valid_2_pad ;  
   wire [4:0] sectored_entries_0_6_valid_2_shl ;  
   wire [19:0] sectored_entries_0_6_valid_2_pad ;  
   wire [1:0] superpage_entries_2_valid_0_shl ;  
   wire [19:0] superpage_entries_2_valid_0_pad ;  
   wire [5:0] sectored_entries_0_6_valid_3_shl ;  
   wire [19:0] sectored_entries_0_6_valid_3_pad ;  
   wire [5:0] sectored_entries_0_6_valid_0_shl ;  
   wire [19:0] sectored_entries_0_6_valid_0_pad ;  
   wire [4:0] sectored_entries_0_7_valid_2_shl ;  
   wire [19:0] sectored_entries_0_7_valid_2_pad ;  
   wire [14:0] superpage_entries_0_level_shl ;  
   wire [19:0] superpage_entries_0_level_pad ;  
   wire [14:0] superpage_entries_1_level_shl ;  
   wire [19:0] superpage_entries_1_level_pad ;  
   wire [5:0] sectored_entries_0_5_valid_0_shl ;  
   wire [19:0] sectored_entries_0_5_valid_0_pad ;  
   wire [19:0] TLB_1_xor64 ;  
   wire [19:0] TLB_1_xor31 ;  
   wire [19:0] TLB_1_xor65 ;  
   wire [19:0] TLB_1_xor66 ;  
   wire [19:0] TLB_1_xor32 ;  
   wire [19:0] TLB_1_xor15 ;  
   wire [19:0] TLB_1_xor68 ;  
   wire [19:0] TLB_1_xor33 ;  
   wire [19:0] TLB_1_xor69 ;  
   wire [19:0] TLB_1_xor70 ;  
   wire [19:0] TLB_1_xor34 ;  
   wire [19:0] TLB_1_xor16 ;  
   wire [19:0] TLB_1_xor7 ;  
   wire [19:0] TLB_1_xor72 ;  
   wire [19:0] TLB_1_xor35 ;  
   wire [19:0] TLB_1_xor73 ;  
   wire [19:0] TLB_1_xor74 ;  
   wire [19:0] TLB_1_xor36 ;  
   wire [19:0] TLB_1_xor17 ;  
   wire [19:0] TLB_1_xor75 ;  
   wire [19:0] TLB_1_xor76 ;  
   wire [19:0] TLB_1_xor37 ;  
   wire [19:0] TLB_1_xor77 ;  
   wire [19:0] TLB_1_xor78 ;  
   wire [19:0] TLB_1_xor38 ;  
   wire [19:0] TLB_1_xor18 ;  
   wire [19:0] TLB_1_xor8 ;  
   wire [19:0] TLB_1_xor3 ;  
   wire [19:0] TLB_1_xor80 ;  
   wire [19:0] TLB_1_xor39 ;  
   wire [19:0] TLB_1_xor81 ;  
   wire [19:0] TLB_1_xor82 ;  
   wire [19:0] TLB_1_xor40 ;  
   wire [19:0] TLB_1_xor19 ;  
   wire [19:0] TLB_1_xor84 ;  
   wire [19:0] TLB_1_xor41 ;  
   wire [19:0] TLB_1_xor85 ;  
   wire [19:0] TLB_1_xor86 ;  
   wire [19:0] TLB_1_xor42 ;  
   wire [19:0] TLB_1_xor20 ;  
   wire [19:0] TLB_1_xor9 ;  
   wire [19:0] TLB_1_xor88 ;  
   wire [19:0] TLB_1_xor43 ;  
   wire [19:0] TLB_1_xor89 ;  
   wire [19:0] TLB_1_xor90 ;  
   wire [19:0] TLB_1_xor44 ;  
   wire [19:0] TLB_1_xor21 ;  
   wire [19:0] TLB_1_xor91 ;  
   wire [19:0] TLB_1_xor92 ;  
   wire [19:0] TLB_1_xor45 ;  
   wire [19:0] TLB_1_xor93 ;  
   wire [19:0] TLB_1_xor94 ;  
   wire [19:0] TLB_1_xor46 ;  
   wire [19:0] TLB_1_xor22 ;  
   wire [19:0] TLB_1_xor10 ;  
   wire [19:0] TLB_1_xor4 ;  
   wire [19:0] TLB_1_xor1 ;  
   wire [19:0] TLB_1_xor96 ;  
   wire [19:0] TLB_1_xor47 ;  
   wire [19:0] TLB_1_xor97 ;  
   wire [19:0] TLB_1_xor98 ;  
   wire [19:0] TLB_1_xor48 ;  
   wire [19:0] TLB_1_xor23 ;  
   wire [19:0] TLB_1_xor100 ;  
   wire [19:0] TLB_1_xor49 ;  
   wire [19:0] TLB_1_xor101 ;  
   wire [19:0] TLB_1_xor102 ;  
   wire [19:0] TLB_1_xor50 ;  
   wire [19:0] TLB_1_xor24 ;  
   wire [19:0] TLB_1_xor11 ;  
   wire [19:0] TLB_1_xor104 ;  
   wire [19:0] TLB_1_xor51 ;  
   wire [19:0] TLB_1_xor105 ;  
   wire [19:0] TLB_1_xor106 ;  
   wire [19:0] TLB_1_xor52 ;  
   wire [19:0] TLB_1_xor25 ;  
   wire [19:0] TLB_1_xor107 ;  
   wire [19:0] TLB_1_xor108 ;  
   wire [19:0] TLB_1_xor53 ;  
   wire [19:0] TLB_1_xor109 ;  
   wire [19:0] TLB_1_xor110 ;  
   wire [19:0] TLB_1_xor54 ;  
   wire [19:0] TLB_1_xor26 ;  
   wire [19:0] TLB_1_xor12 ;  
   wire [19:0] TLB_1_xor5 ;  
   wire [19:0] TLB_1_xor112 ;  
   wire [19:0] TLB_1_xor55 ;  
   wire [19:0] TLB_1_xor113 ;  
   wire [19:0] TLB_1_xor114 ;  
   wire [19:0] TLB_1_xor56 ;  
   wire [19:0] TLB_1_xor27 ;  
   wire [19:0] TLB_1_xor116 ;  
   wire [19:0] TLB_1_xor57 ;  
   wire [19:0] TLB_1_xor117 ;  
   wire [19:0] TLB_1_xor118 ;  
   wire [19:0] TLB_1_xor58 ;  
   wire [19:0] TLB_1_xor28 ;  
   wire [19:0] TLB_1_xor13 ;  
   wire [19:0] TLB_1_xor120 ;  
   wire [19:0] TLB_1_xor59 ;  
   wire [19:0] TLB_1_xor121 ;  
   wire [19:0] TLB_1_xor122 ;  
   wire [19:0] TLB_1_xor60 ;  
   wire [19:0] TLB_1_xor29 ;  
   wire [19:0] TLB_1_xor123 ;  
   wire [19:0] TLB_1_xor124 ;  
   wire [19:0] TLB_1_xor61 ;  
   wire [19:0] TLB_1_xor125 ;  
   wire [19:0] TLB_1_xor126 ;  
   wire [19:0] TLB_1_xor62 ;  
   wire [19:0] TLB_1_xor30 ;  
   wire [19:0] TLB_1_xor14 ;  
   wire [19:0] TLB_1_xor6 ;  
   wire [19:0] TLB_1_xor2 ;  
   wire [19:0] TLB_1_xor0 ;  
   wire [29:0] mpu_ppn_barrier_sum ;  
   wire [29:0] entries_barrier_10_sum ;  
   wire [29:0] entries_barrier_9_sum ;  
   wire [29:0] entries_barrier_7_sum ;  
   wire [29:0] entries_barrier_sum ;  
   wire [29:0] pmp_sum ;  
   wire [29:0] entries_barrier_6_sum ;  
   wire [29:0] entries_barrier_12_sum ;  
   wire [29:0] entries_barrier_1_sum ;  
   wire [29:0] entries_barrier_11_sum ;  
   wire [29:0] entries_barrier_8_sum ;  
   wire [29:0] entries_barrier_2_sum ;  
   wire [29:0] entries_barrier_4_sum ;  
   wire [29:0] entries_barrier_5_sum ;  
   wire [29:0] entries_barrier_3_sum ;  
   wire stopEn0 ;  
   wire entries_barrier_11_metaAssert_wire ;  
   wire entries_barrier_8_metaAssert_wire ;  
   wire entries_barrier_3_metaAssert_wire ;  
   wire pmp_metaAssert_wire ;  
   wire entries_barrier_6_metaAssert_wire ;  
   wire entries_barrier_12_metaAssert_wire ;  
   wire entries_barrier_9_metaAssert_wire ;  
   wire mpu_ppn_barrier_metaAssert_wire ;  
   wire entries_barrier_7_metaAssert_wire ;  
   wire entries_barrier_metaAssert_wire ;  
   wire entries_barrier_5_metaAssert_wire ;  
   wire entries_barrier_2_metaAssert_wire ;  
   wire entries_barrier_4_metaAssert_wire ;  
   wire entries_barrier_1_metaAssert_wire ;  
   wire entries_barrier_10_metaAssert_wire ;  
   wire TLB_1_or7 ;  
   wire TLB_1_or8 ;  
   wire TLB_1_or3 ;  
   wire TLB_1_or9 ;  
   wire TLB_1_or10 ;  
   wire TLB_1_or4 ;  
   wire TLB_1_or1 ;  
   wire TLB_1_or11 ;  
   wire TLB_1_or12 ;  
   wire TLB_1_or5 ;  
   wire TLB_1_or13 ;  
   wire TLB_1_or14 ;  
   wire TLB_1_or6 ;  
   wire TLB_1_or2 ;  
   wire TLB_1_or0 ;  
   reg TLB_1_metaAssert ;  
   reg [31:0] _RAND_103 ;  
  OptimizationBarrier mpu_ppn_barrier(.io_x_ppn(mpu_ppn_barrier_io_x_ppn),.io_x_u(mpu_ppn_barrier_io_x_u),.io_x_ae(mpu_ppn_barrier_io_x_ae),.io_x_sw(mpu_ppn_barrier_io_x_sw),.io_x_sx(mpu_ppn_barrier_io_x_sx),.io_x_sr(mpu_ppn_barrier_io_x_sr),.io_x_pw(mpu_ppn_barrier_io_x_pw),.io_x_px(mpu_ppn_barrier_io_x_px),.io_x_pr(mpu_ppn_barrier_io_x_pr),.io_x_ppp(mpu_ppn_barrier_io_x_ppp),.io_x_pal(mpu_ppn_barrier_io_x_pal),.io_x_paa(mpu_ppn_barrier_io_x_paa),.io_x_eff(mpu_ppn_barrier_io_x_eff),.io_x_c(mpu_ppn_barrier_io_x_c),.io_y_ppn(mpu_ppn_barrier_io_y_ppn),.io_y_u(mpu_ppn_barrier_io_y_u),.io_y_ae(mpu_ppn_barrier_io_y_ae),.io_y_sw(mpu_ppn_barrier_io_y_sw),.io_y_sx(mpu_ppn_barrier_io_y_sx),.io_y_sr(mpu_ppn_barrier_io_y_sr),.io_y_pw(mpu_ppn_barrier_io_y_pw),.io_y_px(mpu_ppn_barrier_io_y_px),.io_y_pr(mpu_ppn_barrier_io_y_pr),.io_y_ppp(mpu_ppn_barrier_io_y_ppp),.io_y_pal(mpu_ppn_barrier_io_y_pal),.io_y_paa(mpu_ppn_barrier_io_y_paa),.io_y_eff(mpu_ppn_barrier_io_y_eff),.io_y_c(mpu_ppn_barrier_io_y_c),.io_covSum(mpu_ppn_barrier_io_covSum),.metaAssert(mpu_ppn_barrier_metaAssert)); 
  PMPChecker_2 pmp(.io_prv(pmp_io_prv),.io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),.io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),.io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),.io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),.io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),.io_pmp_0_addr(pmp_io_pmp_0_addr),.io_pmp_0_mask(pmp_io_pmp_0_mask),.io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),.io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),.io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),.io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),.io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),.io_pmp_1_addr(pmp_io_pmp_1_addr),.io_pmp_1_mask(pmp_io_pmp_1_mask),.io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),.io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),.io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),.io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),.io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),.io_pmp_2_addr(pmp_io_pmp_2_addr),.io_pmp_2_mask(pmp_io_pmp_2_mask),.io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),.io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),.io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),.io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),.io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),.io_pmp_3_addr(pmp_io_pmp_3_addr),.io_pmp_3_mask(pmp_io_pmp_3_mask),.io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),.io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),.io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),.io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),.io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),.io_pmp_4_addr(pmp_io_pmp_4_addr),.io_pmp_4_mask(pmp_io_pmp_4_mask),.io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),.io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),.io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),.io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),.io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),.io_pmp_5_addr(pmp_io_pmp_5_addr),.io_pmp_5_mask(pmp_io_pmp_5_mask),.io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),.io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),.io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),.io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),.io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),.io_pmp_6_addr(pmp_io_pmp_6_addr),.io_pmp_6_mask(pmp_io_pmp_6_mask),.io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),.io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),.io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),.io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),.io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),.io_pmp_7_addr(pmp_io_pmp_7_addr),.io_pmp_7_mask(pmp_io_pmp_7_mask),.io_addr(pmp_io_addr),.io_r(pmp_io_r),.io_w(pmp_io_w),.io_x(pmp_io_x),.io_covSum(pmp_io_covSum),.metaAssert(pmp_metaAssert)); 
  OptimizationBarrier entries_barrier(.io_x_ppn(entries_barrier_io_x_ppn),.io_x_u(entries_barrier_io_x_u),.io_x_ae(entries_barrier_io_x_ae),.io_x_sw(entries_barrier_io_x_sw),.io_x_sx(entries_barrier_io_x_sx),.io_x_sr(entries_barrier_io_x_sr),.io_x_pw(entries_barrier_io_x_pw),.io_x_px(entries_barrier_io_x_px),.io_x_pr(entries_barrier_io_x_pr),.io_x_ppp(entries_barrier_io_x_ppp),.io_x_pal(entries_barrier_io_x_pal),.io_x_paa(entries_barrier_io_x_paa),.io_x_eff(entries_barrier_io_x_eff),.io_x_c(entries_barrier_io_x_c),.io_y_ppn(entries_barrier_io_y_ppn),.io_y_u(entries_barrier_io_y_u),.io_y_ae(entries_barrier_io_y_ae),.io_y_sw(entries_barrier_io_y_sw),.io_y_sx(entries_barrier_io_y_sx),.io_y_sr(entries_barrier_io_y_sr),.io_y_pw(entries_barrier_io_y_pw),.io_y_px(entries_barrier_io_y_px),.io_y_pr(entries_barrier_io_y_pr),.io_y_ppp(entries_barrier_io_y_ppp),.io_y_pal(entries_barrier_io_y_pal),.io_y_paa(entries_barrier_io_y_paa),.io_y_eff(entries_barrier_io_y_eff),.io_y_c(entries_barrier_io_y_c),.io_covSum(entries_barrier_io_covSum),.metaAssert(entries_barrier_metaAssert)); 
  OptimizationBarrier entries_barrier_1(.io_x_ppn(entries_barrier_1_io_x_ppn),.io_x_u(entries_barrier_1_io_x_u),.io_x_ae(entries_barrier_1_io_x_ae),.io_x_sw(entries_barrier_1_io_x_sw),.io_x_sx(entries_barrier_1_io_x_sx),.io_x_sr(entries_barrier_1_io_x_sr),.io_x_pw(entries_barrier_1_io_x_pw),.io_x_px(entries_barrier_1_io_x_px),.io_x_pr(entries_barrier_1_io_x_pr),.io_x_ppp(entries_barrier_1_io_x_ppp),.io_x_pal(entries_barrier_1_io_x_pal),.io_x_paa(entries_barrier_1_io_x_paa),.io_x_eff(entries_barrier_1_io_x_eff),.io_x_c(entries_barrier_1_io_x_c),.io_y_ppn(entries_barrier_1_io_y_ppn),.io_y_u(entries_barrier_1_io_y_u),.io_y_ae(entries_barrier_1_io_y_ae),.io_y_sw(entries_barrier_1_io_y_sw),.io_y_sx(entries_barrier_1_io_y_sx),.io_y_sr(entries_barrier_1_io_y_sr),.io_y_pw(entries_barrier_1_io_y_pw),.io_y_px(entries_barrier_1_io_y_px),.io_y_pr(entries_barrier_1_io_y_pr),.io_y_ppp(entries_barrier_1_io_y_ppp),.io_y_pal(entries_barrier_1_io_y_pal),.io_y_paa(entries_barrier_1_io_y_paa),.io_y_eff(entries_barrier_1_io_y_eff),.io_y_c(entries_barrier_1_io_y_c),.io_covSum(entries_barrier_1_io_covSum),.metaAssert(entries_barrier_1_metaAssert)); 
  OptimizationBarrier entries_barrier_2(.io_x_ppn(entries_barrier_2_io_x_ppn),.io_x_u(entries_barrier_2_io_x_u),.io_x_ae(entries_barrier_2_io_x_ae),.io_x_sw(entries_barrier_2_io_x_sw),.io_x_sx(entries_barrier_2_io_x_sx),.io_x_sr(entries_barrier_2_io_x_sr),.io_x_pw(entries_barrier_2_io_x_pw),.io_x_px(entries_barrier_2_io_x_px),.io_x_pr(entries_barrier_2_io_x_pr),.io_x_ppp(entries_barrier_2_io_x_ppp),.io_x_pal(entries_barrier_2_io_x_pal),.io_x_paa(entries_barrier_2_io_x_paa),.io_x_eff(entries_barrier_2_io_x_eff),.io_x_c(entries_barrier_2_io_x_c),.io_y_ppn(entries_barrier_2_io_y_ppn),.io_y_u(entries_barrier_2_io_y_u),.io_y_ae(entries_barrier_2_io_y_ae),.io_y_sw(entries_barrier_2_io_y_sw),.io_y_sx(entries_barrier_2_io_y_sx),.io_y_sr(entries_barrier_2_io_y_sr),.io_y_pw(entries_barrier_2_io_y_pw),.io_y_px(entries_barrier_2_io_y_px),.io_y_pr(entries_barrier_2_io_y_pr),.io_y_ppp(entries_barrier_2_io_y_ppp),.io_y_pal(entries_barrier_2_io_y_pal),.io_y_paa(entries_barrier_2_io_y_paa),.io_y_eff(entries_barrier_2_io_y_eff),.io_y_c(entries_barrier_2_io_y_c),.io_covSum(entries_barrier_2_io_covSum),.metaAssert(entries_barrier_2_metaAssert)); 
  OptimizationBarrier entries_barrier_3(.io_x_ppn(entries_barrier_3_io_x_ppn),.io_x_u(entries_barrier_3_io_x_u),.io_x_ae(entries_barrier_3_io_x_ae),.io_x_sw(entries_barrier_3_io_x_sw),.io_x_sx(entries_barrier_3_io_x_sx),.io_x_sr(entries_barrier_3_io_x_sr),.io_x_pw(entries_barrier_3_io_x_pw),.io_x_px(entries_barrier_3_io_x_px),.io_x_pr(entries_barrier_3_io_x_pr),.io_x_ppp(entries_barrier_3_io_x_ppp),.io_x_pal(entries_barrier_3_io_x_pal),.io_x_paa(entries_barrier_3_io_x_paa),.io_x_eff(entries_barrier_3_io_x_eff),.io_x_c(entries_barrier_3_io_x_c),.io_y_ppn(entries_barrier_3_io_y_ppn),.io_y_u(entries_barrier_3_io_y_u),.io_y_ae(entries_barrier_3_io_y_ae),.io_y_sw(entries_barrier_3_io_y_sw),.io_y_sx(entries_barrier_3_io_y_sx),.io_y_sr(entries_barrier_3_io_y_sr),.io_y_pw(entries_barrier_3_io_y_pw),.io_y_px(entries_barrier_3_io_y_px),.io_y_pr(entries_barrier_3_io_y_pr),.io_y_ppp(entries_barrier_3_io_y_ppp),.io_y_pal(entries_barrier_3_io_y_pal),.io_y_paa(entries_barrier_3_io_y_paa),.io_y_eff(entries_barrier_3_io_y_eff),.io_y_c(entries_barrier_3_io_y_c),.io_covSum(entries_barrier_3_io_covSum),.metaAssert(entries_barrier_3_metaAssert)); 
  OptimizationBarrier entries_barrier_4(.io_x_ppn(entries_barrier_4_io_x_ppn),.io_x_u(entries_barrier_4_io_x_u),.io_x_ae(entries_barrier_4_io_x_ae),.io_x_sw(entries_barrier_4_io_x_sw),.io_x_sx(entries_barrier_4_io_x_sx),.io_x_sr(entries_barrier_4_io_x_sr),.io_x_pw(entries_barrier_4_io_x_pw),.io_x_px(entries_barrier_4_io_x_px),.io_x_pr(entries_barrier_4_io_x_pr),.io_x_ppp(entries_barrier_4_io_x_ppp),.io_x_pal(entries_barrier_4_io_x_pal),.io_x_paa(entries_barrier_4_io_x_paa),.io_x_eff(entries_barrier_4_io_x_eff),.io_x_c(entries_barrier_4_io_x_c),.io_y_ppn(entries_barrier_4_io_y_ppn),.io_y_u(entries_barrier_4_io_y_u),.io_y_ae(entries_barrier_4_io_y_ae),.io_y_sw(entries_barrier_4_io_y_sw),.io_y_sx(entries_barrier_4_io_y_sx),.io_y_sr(entries_barrier_4_io_y_sr),.io_y_pw(entries_barrier_4_io_y_pw),.io_y_px(entries_barrier_4_io_y_px),.io_y_pr(entries_barrier_4_io_y_pr),.io_y_ppp(entries_barrier_4_io_y_ppp),.io_y_pal(entries_barrier_4_io_y_pal),.io_y_paa(entries_barrier_4_io_y_paa),.io_y_eff(entries_barrier_4_io_y_eff),.io_y_c(entries_barrier_4_io_y_c),.io_covSum(entries_barrier_4_io_covSum),.metaAssert(entries_barrier_4_metaAssert)); 
  OptimizationBarrier entries_barrier_5(.io_x_ppn(entries_barrier_5_io_x_ppn),.io_x_u(entries_barrier_5_io_x_u),.io_x_ae(entries_barrier_5_io_x_ae),.io_x_sw(entries_barrier_5_io_x_sw),.io_x_sx(entries_barrier_5_io_x_sx),.io_x_sr(entries_barrier_5_io_x_sr),.io_x_pw(entries_barrier_5_io_x_pw),.io_x_px(entries_barrier_5_io_x_px),.io_x_pr(entries_barrier_5_io_x_pr),.io_x_ppp(entries_barrier_5_io_x_ppp),.io_x_pal(entries_barrier_5_io_x_pal),.io_x_paa(entries_barrier_5_io_x_paa),.io_x_eff(entries_barrier_5_io_x_eff),.io_x_c(entries_barrier_5_io_x_c),.io_y_ppn(entries_barrier_5_io_y_ppn),.io_y_u(entries_barrier_5_io_y_u),.io_y_ae(entries_barrier_5_io_y_ae),.io_y_sw(entries_barrier_5_io_y_sw),.io_y_sx(entries_barrier_5_io_y_sx),.io_y_sr(entries_barrier_5_io_y_sr),.io_y_pw(entries_barrier_5_io_y_pw),.io_y_px(entries_barrier_5_io_y_px),.io_y_pr(entries_barrier_5_io_y_pr),.io_y_ppp(entries_barrier_5_io_y_ppp),.io_y_pal(entries_barrier_5_io_y_pal),.io_y_paa(entries_barrier_5_io_y_paa),.io_y_eff(entries_barrier_5_io_y_eff),.io_y_c(entries_barrier_5_io_y_c),.io_covSum(entries_barrier_5_io_covSum),.metaAssert(entries_barrier_5_metaAssert)); 
  OptimizationBarrier entries_barrier_6(.io_x_ppn(entries_barrier_6_io_x_ppn),.io_x_u(entries_barrier_6_io_x_u),.io_x_ae(entries_barrier_6_io_x_ae),.io_x_sw(entries_barrier_6_io_x_sw),.io_x_sx(entries_barrier_6_io_x_sx),.io_x_sr(entries_barrier_6_io_x_sr),.io_x_pw(entries_barrier_6_io_x_pw),.io_x_px(entries_barrier_6_io_x_px),.io_x_pr(entries_barrier_6_io_x_pr),.io_x_ppp(entries_barrier_6_io_x_ppp),.io_x_pal(entries_barrier_6_io_x_pal),.io_x_paa(entries_barrier_6_io_x_paa),.io_x_eff(entries_barrier_6_io_x_eff),.io_x_c(entries_barrier_6_io_x_c),.io_y_ppn(entries_barrier_6_io_y_ppn),.io_y_u(entries_barrier_6_io_y_u),.io_y_ae(entries_barrier_6_io_y_ae),.io_y_sw(entries_barrier_6_io_y_sw),.io_y_sx(entries_barrier_6_io_y_sx),.io_y_sr(entries_barrier_6_io_y_sr),.io_y_pw(entries_barrier_6_io_y_pw),.io_y_px(entries_barrier_6_io_y_px),.io_y_pr(entries_barrier_6_io_y_pr),.io_y_ppp(entries_barrier_6_io_y_ppp),.io_y_pal(entries_barrier_6_io_y_pal),.io_y_paa(entries_barrier_6_io_y_paa),.io_y_eff(entries_barrier_6_io_y_eff),.io_y_c(entries_barrier_6_io_y_c),.io_covSum(entries_barrier_6_io_covSum),.metaAssert(entries_barrier_6_metaAssert)); 
  OptimizationBarrier entries_barrier_7(.io_x_ppn(entries_barrier_7_io_x_ppn),.io_x_u(entries_barrier_7_io_x_u),.io_x_ae(entries_barrier_7_io_x_ae),.io_x_sw(entries_barrier_7_io_x_sw),.io_x_sx(entries_barrier_7_io_x_sx),.io_x_sr(entries_barrier_7_io_x_sr),.io_x_pw(entries_barrier_7_io_x_pw),.io_x_px(entries_barrier_7_io_x_px),.io_x_pr(entries_barrier_7_io_x_pr),.io_x_ppp(entries_barrier_7_io_x_ppp),.io_x_pal(entries_barrier_7_io_x_pal),.io_x_paa(entries_barrier_7_io_x_paa),.io_x_eff(entries_barrier_7_io_x_eff),.io_x_c(entries_barrier_7_io_x_c),.io_y_ppn(entries_barrier_7_io_y_ppn),.io_y_u(entries_barrier_7_io_y_u),.io_y_ae(entries_barrier_7_io_y_ae),.io_y_sw(entries_barrier_7_io_y_sw),.io_y_sx(entries_barrier_7_io_y_sx),.io_y_sr(entries_barrier_7_io_y_sr),.io_y_pw(entries_barrier_7_io_y_pw),.io_y_px(entries_barrier_7_io_y_px),.io_y_pr(entries_barrier_7_io_y_pr),.io_y_ppp(entries_barrier_7_io_y_ppp),.io_y_pal(entries_barrier_7_io_y_pal),.io_y_paa(entries_barrier_7_io_y_paa),.io_y_eff(entries_barrier_7_io_y_eff),.io_y_c(entries_barrier_7_io_y_c),.io_covSum(entries_barrier_7_io_covSum),.metaAssert(entries_barrier_7_metaAssert)); 
  OptimizationBarrier entries_barrier_8(.io_x_ppn(entries_barrier_8_io_x_ppn),.io_x_u(entries_barrier_8_io_x_u),.io_x_ae(entries_barrier_8_io_x_ae),.io_x_sw(entries_barrier_8_io_x_sw),.io_x_sx(entries_barrier_8_io_x_sx),.io_x_sr(entries_barrier_8_io_x_sr),.io_x_pw(entries_barrier_8_io_x_pw),.io_x_px(entries_barrier_8_io_x_px),.io_x_pr(entries_barrier_8_io_x_pr),.io_x_ppp(entries_barrier_8_io_x_ppp),.io_x_pal(entries_barrier_8_io_x_pal),.io_x_paa(entries_barrier_8_io_x_paa),.io_x_eff(entries_barrier_8_io_x_eff),.io_x_c(entries_barrier_8_io_x_c),.io_y_ppn(entries_barrier_8_io_y_ppn),.io_y_u(entries_barrier_8_io_y_u),.io_y_ae(entries_barrier_8_io_y_ae),.io_y_sw(entries_barrier_8_io_y_sw),.io_y_sx(entries_barrier_8_io_y_sx),.io_y_sr(entries_barrier_8_io_y_sr),.io_y_pw(entries_barrier_8_io_y_pw),.io_y_px(entries_barrier_8_io_y_px),.io_y_pr(entries_barrier_8_io_y_pr),.io_y_ppp(entries_barrier_8_io_y_ppp),.io_y_pal(entries_barrier_8_io_y_pal),.io_y_paa(entries_barrier_8_io_y_paa),.io_y_eff(entries_barrier_8_io_y_eff),.io_y_c(entries_barrier_8_io_y_c),.io_covSum(entries_barrier_8_io_covSum),.metaAssert(entries_barrier_8_metaAssert)); 
  OptimizationBarrier entries_barrier_9(.io_x_ppn(entries_barrier_9_io_x_ppn),.io_x_u(entries_barrier_9_io_x_u),.io_x_ae(entries_barrier_9_io_x_ae),.io_x_sw(entries_barrier_9_io_x_sw),.io_x_sx(entries_barrier_9_io_x_sx),.io_x_sr(entries_barrier_9_io_x_sr),.io_x_pw(entries_barrier_9_io_x_pw),.io_x_px(entries_barrier_9_io_x_px),.io_x_pr(entries_barrier_9_io_x_pr),.io_x_ppp(entries_barrier_9_io_x_ppp),.io_x_pal(entries_barrier_9_io_x_pal),.io_x_paa(entries_barrier_9_io_x_paa),.io_x_eff(entries_barrier_9_io_x_eff),.io_x_c(entries_barrier_9_io_x_c),.io_y_ppn(entries_barrier_9_io_y_ppn),.io_y_u(entries_barrier_9_io_y_u),.io_y_ae(entries_barrier_9_io_y_ae),.io_y_sw(entries_barrier_9_io_y_sw),.io_y_sx(entries_barrier_9_io_y_sx),.io_y_sr(entries_barrier_9_io_y_sr),.io_y_pw(entries_barrier_9_io_y_pw),.io_y_px(entries_barrier_9_io_y_px),.io_y_pr(entries_barrier_9_io_y_pr),.io_y_ppp(entries_barrier_9_io_y_ppp),.io_y_pal(entries_barrier_9_io_y_pal),.io_y_paa(entries_barrier_9_io_y_paa),.io_y_eff(entries_barrier_9_io_y_eff),.io_y_c(entries_barrier_9_io_y_c),.io_covSum(entries_barrier_9_io_covSum),.metaAssert(entries_barrier_9_metaAssert)); 
  OptimizationBarrier entries_barrier_10(.io_x_ppn(entries_barrier_10_io_x_ppn),.io_x_u(entries_barrier_10_io_x_u),.io_x_ae(entries_barrier_10_io_x_ae),.io_x_sw(entries_barrier_10_io_x_sw),.io_x_sx(entries_barrier_10_io_x_sx),.io_x_sr(entries_barrier_10_io_x_sr),.io_x_pw(entries_barrier_10_io_x_pw),.io_x_px(entries_barrier_10_io_x_px),.io_x_pr(entries_barrier_10_io_x_pr),.io_x_ppp(entries_barrier_10_io_x_ppp),.io_x_pal(entries_barrier_10_io_x_pal),.io_x_paa(entries_barrier_10_io_x_paa),.io_x_eff(entries_barrier_10_io_x_eff),.io_x_c(entries_barrier_10_io_x_c),.io_y_ppn(entries_barrier_10_io_y_ppn),.io_y_u(entries_barrier_10_io_y_u),.io_y_ae(entries_barrier_10_io_y_ae),.io_y_sw(entries_barrier_10_io_y_sw),.io_y_sx(entries_barrier_10_io_y_sx),.io_y_sr(entries_barrier_10_io_y_sr),.io_y_pw(entries_barrier_10_io_y_pw),.io_y_px(entries_barrier_10_io_y_px),.io_y_pr(entries_barrier_10_io_y_pr),.io_y_ppp(entries_barrier_10_io_y_ppp),.io_y_pal(entries_barrier_10_io_y_pal),.io_y_paa(entries_barrier_10_io_y_paa),.io_y_eff(entries_barrier_10_io_y_eff),.io_y_c(entries_barrier_10_io_y_c),.io_covSum(entries_barrier_10_io_covSum),.metaAssert(entries_barrier_10_metaAssert)); 
  OptimizationBarrier entries_barrier_11(.io_x_ppn(entries_barrier_11_io_x_ppn),.io_x_u(entries_barrier_11_io_x_u),.io_x_ae(entries_barrier_11_io_x_ae),.io_x_sw(entries_barrier_11_io_x_sw),.io_x_sx(entries_barrier_11_io_x_sx),.io_x_sr(entries_barrier_11_io_x_sr),.io_x_pw(entries_barrier_11_io_x_pw),.io_x_px(entries_barrier_11_io_x_px),.io_x_pr(entries_barrier_11_io_x_pr),.io_x_ppp(entries_barrier_11_io_x_ppp),.io_x_pal(entries_barrier_11_io_x_pal),.io_x_paa(entries_barrier_11_io_x_paa),.io_x_eff(entries_barrier_11_io_x_eff),.io_x_c(entries_barrier_11_io_x_c),.io_y_ppn(entries_barrier_11_io_y_ppn),.io_y_u(entries_barrier_11_io_y_u),.io_y_ae(entries_barrier_11_io_y_ae),.io_y_sw(entries_barrier_11_io_y_sw),.io_y_sx(entries_barrier_11_io_y_sx),.io_y_sr(entries_barrier_11_io_y_sr),.io_y_pw(entries_barrier_11_io_y_pw),.io_y_px(entries_barrier_11_io_y_px),.io_y_pr(entries_barrier_11_io_y_pr),.io_y_ppp(entries_barrier_11_io_y_ppp),.io_y_pal(entries_barrier_11_io_y_pal),.io_y_paa(entries_barrier_11_io_y_paa),.io_y_eff(entries_barrier_11_io_y_eff),.io_y_c(entries_barrier_11_io_y_c),.io_covSum(entries_barrier_11_io_covSum),.metaAssert(entries_barrier_11_metaAssert)); 
  OptimizationBarrier entries_barrier_12(.io_x_ppn(entries_barrier_12_io_x_ppn),.io_x_u(entries_barrier_12_io_x_u),.io_x_ae(entries_barrier_12_io_x_ae),.io_x_sw(entries_barrier_12_io_x_sw),.io_x_sx(entries_barrier_12_io_x_sx),.io_x_sr(entries_barrier_12_io_x_sr),.io_x_pw(entries_barrier_12_io_x_pw),.io_x_px(entries_barrier_12_io_x_px),.io_x_pr(entries_barrier_12_io_x_pr),.io_x_ppp(entries_barrier_12_io_x_ppp),.io_x_pal(entries_barrier_12_io_x_pal),.io_x_paa(entries_barrier_12_io_x_paa),.io_x_eff(entries_barrier_12_io_x_eff),.io_x_c(entries_barrier_12_io_x_c),.io_y_ppn(entries_barrier_12_io_y_ppn),.io_y_u(entries_barrier_12_io_y_u),.io_y_ae(entries_barrier_12_io_y_ae),.io_y_sw(entries_barrier_12_io_y_sw),.io_y_sx(entries_barrier_12_io_y_sx),.io_y_sr(entries_barrier_12_io_y_sr),.io_y_pw(entries_barrier_12_io_y_pw),.io_y_px(entries_barrier_12_io_y_px),.io_y_pr(entries_barrier_12_io_y_pr),.io_y_ppp(entries_barrier_12_io_y_ppp),.io_y_pal(entries_barrier_12_io_y_pal),.io_y_paa(entries_barrier_12_io_y_paa),.io_y_eff(entries_barrier_12_io_y_eff),.io_y_c(entries_barrier_12_io_y_c),.io_covSum(entries_barrier_12_io_covSum),.metaAssert(entries_barrier_12_metaAssert)); 
  assign vpn=io_req_bits_vaddr[38:12]; 
  assign priv_s=io_ptw_status_prv[0]; 
  assign priv_uses_vm=io_ptw_status_prv<=2'h1; 
  assign vm_enabled=io_ptw_ptbr_mode[3]&priv_uses_vm; 
  assign refill_ppn=io_ptw_resp_bits_pte_ppn[19:0]; 
  assign _invalidate_refill_T=state==2'h1; 
  assign _invalidate_refill_T_1=state==2'h3; 
  assign _invalidate_refill_T_2=_invalidate_refill_T|_invalidate_refill_T_1; 
  assign invalidate_refill=_invalidate_refill_T_2|io_sfence_valid; 
  assign mpu_ppn_hi=mpu_ppn_barrier_io_y_ppn[19:18]; 
  assign mpu_ppn_ignore=special_entry_level<2'h1; 
  assign _mpu_ppn_T_17=mpu_ppn_ignore ? vpn:27'h0; 
  assign _GEN_919={7'b0,mpu_ppn_barrier_io_y_ppn}; 
  assign _mpu_ppn_T_18=_mpu_ppn_T_17|_GEN_919; 
  assign mpu_ppn_lo=_mpu_ppn_T_18[17:9]; 
  assign mpu_ppn_ignore_1=special_entry_level<2'h2; 
  assign _mpu_ppn_T_19=mpu_ppn_ignore_1 ? vpn:27'h0; 
  assign _mpu_ppn_T_20=_mpu_ppn_T_19|_GEN_919; 
  assign mpu_ppn_lo_1=_mpu_ppn_T_20[8:0]; 
  assign _mpu_ppn_T_21={mpu_ppn_hi,mpu_ppn_lo,mpu_ppn_lo_1}; 
  assign _mpu_ppn_T_23=vm_enabled ? {8'b0,_mpu_ppn_T_21}:io_req_bits_vaddr[39:12]; 
  assign mpu_ppn=io_ptw_resp_valid ? {8'b0,refill_ppn}:_mpu_ppn_T_23; 
  assign mpu_physaddr_lo=io_req_bits_vaddr[11:0]; 
  assign mpu_physaddr={mpu_ppn,mpu_physaddr_lo}; 
  assign _mpu_priv_T_2={io_ptw_status_debug,io_ptw_status_prv}; 
  assign mpu_priv=io_ptw_resp_valid ? 3'h1:_mpu_priv_T_2; 
  assign _legal_address_T=mpu_physaddr^40'h3000; 
  assign _legal_address_T_1={1'b0,$signed(_legal_address_T)}; 
  assign _legal_address_T_3=$signed(_legal_address_T_1)&-41'sh1000; 
  assign _legal_address_T_4=$signed(_legal_address_T_3)==41'sh0; 
  assign _legal_address_T_5=mpu_physaddr^40'hc000000; 
  assign _legal_address_T_6={1'b0,$signed(_legal_address_T_5)}; 
  assign _legal_address_T_8=$signed(_legal_address_T_6)&-41'sh4000000; 
  assign _legal_address_T_9=$signed(_legal_address_T_8)==41'sh0; 
  assign _legal_address_T_10=mpu_physaddr^40'h2000000; 
  assign _legal_address_T_11={1'b0,$signed(_legal_address_T_10)}; 
  assign _legal_address_T_13=$signed(_legal_address_T_11)&-41'sh10000; 
  assign _legal_address_T_14=$signed(_legal_address_T_13)==41'sh0; 
  assign _legal_address_T_16={1'b0,$signed(mpu_physaddr)}; 
  assign _legal_address_T_18=$signed(_legal_address_T_16)&-41'sh1000; 
  assign _legal_address_T_19=$signed(_legal_address_T_18)==41'sh0; 
  assign _legal_address_T_20=mpu_physaddr^40'h10000; 
  assign _legal_address_T_21={1'b0,$signed(_legal_address_T_20)}; 
  assign _legal_address_T_23=$signed(_legal_address_T_21)&-41'sh10000; 
  assign _legal_address_T_24=$signed(_legal_address_T_23)==41'sh0; 
  assign _legal_address_T_25=mpu_physaddr^40'h80000000; 
  assign _legal_address_T_26={1'b0,$signed(_legal_address_T_25)}; 
  assign _legal_address_T_28=$signed(_legal_address_T_26)&-41'sh10000000; 
  assign _legal_address_T_29=$signed(_legal_address_T_28)==41'sh0; 
  assign _legal_address_T_30=mpu_physaddr^40'h60000000; 
  assign _legal_address_T_31={1'b0,$signed(_legal_address_T_30)}; 
  assign _legal_address_T_33=$signed(_legal_address_T_31)&-41'sh20000000; 
  assign _legal_address_T_34=$signed(_legal_address_T_33)==41'sh0; 
  assign _legal_address_T_35=_legal_address_T_4|_legal_address_T_9; 
  assign _legal_address_T_36=_legal_address_T_35|_legal_address_T_14; 
  assign _legal_address_T_37=_legal_address_T_36|_legal_address_T_19; 
  assign _legal_address_T_38=_legal_address_T_37|_legal_address_T_24; 
  assign _legal_address_T_39=_legal_address_T_38|_legal_address_T_29; 
  assign legal_address=_legal_address_T_39|_legal_address_T_34; 
  assign _cacheable_T_8=$signed(_legal_address_T_26)&41'sh80000000; 
  assign _cacheable_T_9=$signed(_cacheable_T_8)==41'sh0; 
  assign cacheable=legal_address&_cacheable_T_9; 
  assign _homogeneous_T_54=mpu_physaddr^40'h8000000; 
  assign _homogeneous_T_55={1'b0,$signed(_homogeneous_T_54)}; 
  assign _homogeneous_T_57=$signed(_homogeneous_T_55)&41'shc8000000; 
  assign _homogeneous_T_58=$signed(_homogeneous_T_57)==41'sh0; 
  assign _homogeneous_T_71=$signed(_legal_address_T_16)&41'shc8010000; 
  assign _homogeneous_T_72=$signed(_homogeneous_T_71)==41'sh0; 
  assign _homogeneous_T_79=_homogeneous_T_72|_homogeneous_T_58; 
  assign _deny_access_to_debug_T=mpu_priv<=3'h3; 
  assign deny_access_to_debug=_deny_access_to_debug_T&_legal_address_T_19; 
  assign _prot_r_T_7=legal_address&~deny_access_to_debug; 
  assign prot_r=_prot_r_T_7&pmp_io_r; 
  assign _prot_w_T_10=mpu_physaddr^40'h40000000; 
  assign _prot_w_T_11={1'b0,$signed(_prot_w_T_10)}; 
  assign _prot_w_T_13=$signed(_prot_w_T_11)&41'shc0000000; 
  assign _prot_w_T_14=$signed(_prot_w_T_13)==41'sh0; 
  assign _prot_w_T_18=$signed(_legal_address_T_26)&41'shc0000000; 
  assign _prot_w_T_19=$signed(_prot_w_T_18)==41'sh0; 
  assign _prot_w_T_21=_homogeneous_T_79|_prot_w_T_14; 
  assign _prot_w_T_22=_prot_w_T_21|_prot_w_T_19; 
  assign _prot_w_T_31=legal_address&_prot_w_T_22; 
  assign _prot_w_T_33=_prot_w_T_31&~deny_access_to_debug; 
  assign prot_w=_prot_w_T_33&pmp_io_w; 
  assign prot_al=legal_address&_homogeneous_T_79; 
  assign _prot_x_T_3=$signed(_legal_address_T_16)&41'shca000000; 
  assign _prot_x_T_4=$signed(_prot_x_T_3)==41'sh0; 
  assign _prot_x_T_15=_prot_x_T_4|_prot_w_T_14; 
  assign _prot_x_T_16=_prot_x_T_15|_prot_w_T_19; 
  assign _prot_x_T_31=legal_address&_prot_x_T_16; 
  assign _prot_x_T_33=_prot_x_T_31&~deny_access_to_debug; 
  assign prot_x=_prot_x_T_33&pmp_io_x; 
  assign _prot_eff_T_20=$signed(_legal_address_T_16)&41'shca012000; 
  assign _prot_eff_T_21=$signed(_prot_eff_T_20)==41'sh0; 
  assign _prot_eff_T_25=$signed(_legal_address_T_11)&41'shca010000; 
  assign _prot_eff_T_26=$signed(_prot_eff_T_25)==41'sh0; 
  assign _prot_eff_T_37=_prot_eff_T_21|_prot_eff_T_26; 
  assign _prot_eff_T_38=_prot_eff_T_37|_homogeneous_T_58; 
  assign _prot_eff_T_39=_prot_eff_T_38|_prot_w_T_14; 
  assign prot_eff=legal_address&_prot_eff_T_39; 
  assign _sector_hits_T=sectored_entries_0_0_valid_0|sectored_entries_0_0_valid_1; 
  assign _sector_hits_T_1=_sector_hits_T|sectored_entries_0_0_valid_2; 
  assign _sector_hits_T_2=_sector_hits_T_1|sectored_entries_0_0_valid_3; 
  assign _sector_hits_T_3=sectored_entries_0_0_tag^vpn; 
  assign _sector_hits_T_5=_sector_hits_T_3[26:2]==25'h0; 
  assign sector_hits_0=_sector_hits_T_2&_sector_hits_T_5; 
  assign _sector_hits_T_6=sectored_entries_0_1_valid_0|sectored_entries_0_1_valid_1; 
  assign _sector_hits_T_7=_sector_hits_T_6|sectored_entries_0_1_valid_2; 
  assign _sector_hits_T_8=_sector_hits_T_7|sectored_entries_0_1_valid_3; 
  assign _sector_hits_T_9=sectored_entries_0_1_tag^vpn; 
  assign _sector_hits_T_11=_sector_hits_T_9[26:2]==25'h0; 
  assign sector_hits_1=_sector_hits_T_8&_sector_hits_T_11; 
  assign _sector_hits_T_12=sectored_entries_0_2_valid_0|sectored_entries_0_2_valid_1; 
  assign _sector_hits_T_13=_sector_hits_T_12|sectored_entries_0_2_valid_2; 
  assign _sector_hits_T_14=_sector_hits_T_13|sectored_entries_0_2_valid_3; 
  assign _sector_hits_T_15=sectored_entries_0_2_tag^vpn; 
  assign _sector_hits_T_17=_sector_hits_T_15[26:2]==25'h0; 
  assign sector_hits_2=_sector_hits_T_14&_sector_hits_T_17; 
  assign _sector_hits_T_18=sectored_entries_0_3_valid_0|sectored_entries_0_3_valid_1; 
  assign _sector_hits_T_19=_sector_hits_T_18|sectored_entries_0_3_valid_2; 
  assign _sector_hits_T_20=_sector_hits_T_19|sectored_entries_0_3_valid_3; 
  assign _sector_hits_T_21=sectored_entries_0_3_tag^vpn; 
  assign _sector_hits_T_23=_sector_hits_T_21[26:2]==25'h0; 
  assign sector_hits_3=_sector_hits_T_20&_sector_hits_T_23; 
  assign _sector_hits_T_24=sectored_entries_0_4_valid_0|sectored_entries_0_4_valid_1; 
  assign _sector_hits_T_25=_sector_hits_T_24|sectored_entries_0_4_valid_2; 
  assign _sector_hits_T_26=_sector_hits_T_25|sectored_entries_0_4_valid_3; 
  assign _sector_hits_T_27=sectored_entries_0_4_tag^vpn; 
  assign _sector_hits_T_29=_sector_hits_T_27[26:2]==25'h0; 
  assign sector_hits_4=_sector_hits_T_26&_sector_hits_T_29; 
  assign _sector_hits_T_30=sectored_entries_0_5_valid_0|sectored_entries_0_5_valid_1; 
  assign _sector_hits_T_31=_sector_hits_T_30|sectored_entries_0_5_valid_2; 
  assign _sector_hits_T_32=_sector_hits_T_31|sectored_entries_0_5_valid_3; 
  assign _sector_hits_T_33=sectored_entries_0_5_tag^vpn; 
  assign _sector_hits_T_35=_sector_hits_T_33[26:2]==25'h0; 
  assign sector_hits_5=_sector_hits_T_32&_sector_hits_T_35; 
  assign _sector_hits_T_36=sectored_entries_0_6_valid_0|sectored_entries_0_6_valid_1; 
  assign _sector_hits_T_37=_sector_hits_T_36|sectored_entries_0_6_valid_2; 
  assign _sector_hits_T_38=_sector_hits_T_37|sectored_entries_0_6_valid_3; 
  assign _sector_hits_T_39=sectored_entries_0_6_tag^vpn; 
  assign _sector_hits_T_41=_sector_hits_T_39[26:2]==25'h0; 
  assign sector_hits_6=_sector_hits_T_38&_sector_hits_T_41; 
  assign _sector_hits_T_42=sectored_entries_0_7_valid_0|sectored_entries_0_7_valid_1; 
  assign _sector_hits_T_43=_sector_hits_T_42|sectored_entries_0_7_valid_2; 
  assign _sector_hits_T_44=_sector_hits_T_43|sectored_entries_0_7_valid_3; 
  assign _sector_hits_T_45=sectored_entries_0_7_tag^vpn; 
  assign _sector_hits_T_47=_sector_hits_T_45[26:2]==25'h0; 
  assign sector_hits_7=_sector_hits_T_44&_sector_hits_T_47; 
  assign _superpage_hits_T_2=superpage_entries_0_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_4=superpage_entries_0_valid_0&_superpage_hits_T_2; 
  assign superpage_hits_ignore_1=superpage_entries_0_level<2'h1; 
  assign _superpage_hits_T_7=superpage_entries_0_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_8=superpage_hits_ignore_1|_superpage_hits_T_7; 
  assign superpage_hits_0=_superpage_hits_T_4&_superpage_hits_T_8; 
  assign _superpage_hits_T_16=superpage_entries_1_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_18=superpage_entries_1_valid_0&_superpage_hits_T_16; 
  assign superpage_hits_ignore_4=superpage_entries_1_level<2'h1; 
  assign _superpage_hits_T_21=superpage_entries_1_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_22=superpage_hits_ignore_4|_superpage_hits_T_21; 
  assign superpage_hits_1=_superpage_hits_T_18&_superpage_hits_T_22; 
  assign _superpage_hits_T_30=superpage_entries_2_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_32=superpage_entries_2_valid_0&_superpage_hits_T_30; 
  assign superpage_hits_ignore_7=superpage_entries_2_level<2'h1; 
  assign _superpage_hits_T_35=superpage_entries_2_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_36=superpage_hits_ignore_7|_superpage_hits_T_35; 
  assign superpage_hits_2=_superpage_hits_T_32&_superpage_hits_T_36; 
  assign _superpage_hits_T_44=superpage_entries_3_tag[26:18]==vpn[26:18]; 
  assign _superpage_hits_T_46=superpage_entries_3_valid_0&_superpage_hits_T_44; 
  assign superpage_hits_ignore_10=superpage_entries_3_level<2'h1; 
  assign _superpage_hits_T_49=superpage_entries_3_tag[17:9]==vpn[17:9]; 
  assign _superpage_hits_T_50=superpage_hits_ignore_10|_superpage_hits_T_49; 
  assign superpage_hits_3=_superpage_hits_T_46&_superpage_hits_T_50; 
  assign hitsVec_idx=vpn[1:0]; 
  assign _GEN_1=2'h1==hitsVec_idx ? sectored_entries_0_0_valid_1:sectored_entries_0_0_valid_0; 
  assign _GEN_2=2'h2==hitsVec_idx ? sectored_entries_0_0_valid_2:_GEN_1; 
  assign _GEN_3=2'h3==hitsVec_idx ? sectored_entries_0_0_valid_3:_GEN_2; 
  assign _hitsVec_T_3=_GEN_3&_sector_hits_T_5; 
  assign hitsVec_0=vm_enabled&_hitsVec_T_3; 
  assign _GEN_5=2'h1==hitsVec_idx ? sectored_entries_0_1_valid_1:sectored_entries_0_1_valid_0; 
  assign _GEN_6=2'h2==hitsVec_idx ? sectored_entries_0_1_valid_2:_GEN_5; 
  assign _GEN_7=2'h3==hitsVec_idx ? sectored_entries_0_1_valid_3:_GEN_6; 
  assign _hitsVec_T_7=_GEN_7&_sector_hits_T_11; 
  assign hitsVec_1=vm_enabled&_hitsVec_T_7; 
  assign _GEN_9=2'h1==hitsVec_idx ? sectored_entries_0_2_valid_1:sectored_entries_0_2_valid_0; 
  assign _GEN_10=2'h2==hitsVec_idx ? sectored_entries_0_2_valid_2:_GEN_9; 
  assign _GEN_11=2'h3==hitsVec_idx ? sectored_entries_0_2_valid_3:_GEN_10; 
  assign _hitsVec_T_11=_GEN_11&_sector_hits_T_17; 
  assign hitsVec_2=vm_enabled&_hitsVec_T_11; 
  assign _GEN_13=2'h1==hitsVec_idx ? sectored_entries_0_3_valid_1:sectored_entries_0_3_valid_0; 
  assign _GEN_14=2'h2==hitsVec_idx ? sectored_entries_0_3_valid_2:_GEN_13; 
  assign _GEN_15=2'h3==hitsVec_idx ? sectored_entries_0_3_valid_3:_GEN_14; 
  assign _hitsVec_T_15=_GEN_15&_sector_hits_T_23; 
  assign hitsVec_3=vm_enabled&_hitsVec_T_15; 
  assign _GEN_17=2'h1==hitsVec_idx ? sectored_entries_0_4_valid_1:sectored_entries_0_4_valid_0; 
  assign _GEN_18=2'h2==hitsVec_idx ? sectored_entries_0_4_valid_2:_GEN_17; 
  assign _GEN_19=2'h3==hitsVec_idx ? sectored_entries_0_4_valid_3:_GEN_18; 
  assign _hitsVec_T_19=_GEN_19&_sector_hits_T_29; 
  assign hitsVec_4=vm_enabled&_hitsVec_T_19; 
  assign _GEN_21=2'h1==hitsVec_idx ? sectored_entries_0_5_valid_1:sectored_entries_0_5_valid_0; 
  assign _GEN_22=2'h2==hitsVec_idx ? sectored_entries_0_5_valid_2:_GEN_21; 
  assign _GEN_23=2'h3==hitsVec_idx ? sectored_entries_0_5_valid_3:_GEN_22; 
  assign _hitsVec_T_23=_GEN_23&_sector_hits_T_35; 
  assign hitsVec_5=vm_enabled&_hitsVec_T_23; 
  assign _GEN_25=2'h1==hitsVec_idx ? sectored_entries_0_6_valid_1:sectored_entries_0_6_valid_0; 
  assign _GEN_26=2'h2==hitsVec_idx ? sectored_entries_0_6_valid_2:_GEN_25; 
  assign _GEN_27=2'h3==hitsVec_idx ? sectored_entries_0_6_valid_3:_GEN_26; 
  assign _hitsVec_T_27=_GEN_27&_sector_hits_T_41; 
  assign hitsVec_6=vm_enabled&_hitsVec_T_27; 
  assign _GEN_29=2'h1==hitsVec_idx ? sectored_entries_0_7_valid_1:sectored_entries_0_7_valid_0; 
  assign _GEN_30=2'h2==hitsVec_idx ? sectored_entries_0_7_valid_2:_GEN_29; 
  assign _GEN_31=2'h3==hitsVec_idx ? sectored_entries_0_7_valid_3:_GEN_30; 
  assign _hitsVec_T_31=_GEN_31&_sector_hits_T_47; 
  assign hitsVec_7=vm_enabled&_hitsVec_T_31; 
  assign hitsVec_8=vm_enabled&superpage_hits_0; 
  assign hitsVec_9=vm_enabled&superpage_hits_1; 
  assign hitsVec_10=vm_enabled&superpage_hits_2; 
  assign hitsVec_11=vm_enabled&superpage_hits_3; 
  assign _hitsVec_T_94=special_entry_tag[26:18]==vpn[26:18]; 
  assign _hitsVec_T_96=special_entry_valid_0&_hitsVec_T_94; 
  assign _hitsVec_T_99=special_entry_tag[17:9]==vpn[17:9]; 
  assign _hitsVec_T_100=mpu_ppn_ignore|_hitsVec_T_99; 
  assign _hitsVec_T_101=_hitsVec_T_96&_hitsVec_T_100; 
  assign _hitsVec_T_104=special_entry_tag[8:0]==vpn[8:0]; 
  assign _hitsVec_T_105=mpu_ppn_ignore_1|_hitsVec_T_104; 
  assign _hitsVec_T_106=_hitsVec_T_101&_hitsVec_T_105; 
  assign hitsVec_12=vm_enabled&_hitsVec_T_106; 
  assign real_hits_lo={hitsVec_5,hitsVec_4,hitsVec_3,hitsVec_2,hitsVec_1,hitsVec_0}; 
  assign real_hits={hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; 
  assign hits_hi=~vm_enabled; 
  assign hits={hits_hi,hitsVec_12,hitsVec_11,hitsVec_10,hitsVec_9,hitsVec_8,hitsVec_7,hitsVec_6,real_hits_lo}; 
  assign newEntry_g=io_ptw_resp_bits_pte_g&io_ptw_resp_bits_pte_v; 
  assign _newEntry_sr_T_1=io_ptw_resp_bits_pte_x&~io_ptw_resp_bits_pte_w; 
  assign _newEntry_sr_T_2=io_ptw_resp_bits_pte_r|_newEntry_sr_T_1; 
  assign _newEntry_sr_T_3=io_ptw_resp_bits_pte_v&_newEntry_sr_T_2; 
  assign _newEntry_sr_T_4=_newEntry_sr_T_3&io_ptw_resp_bits_pte_a; 
  assign newEntry_sr=_newEntry_sr_T_4&io_ptw_resp_bits_pte_r; 
  assign _newEntry_sw_T_5=_newEntry_sr_T_4&io_ptw_resp_bits_pte_w; 
  assign newEntry_sw=_newEntry_sw_T_5&io_ptw_resp_bits_pte_d; 
  assign newEntry_sx=_newEntry_sr_T_4&io_ptw_resp_bits_pte_x; 
  assign special_entry_data_0_lo={prot_x,prot_r,_prot_w_T_31,prot_al,prot_al,prot_eff,cacheable,1'h0}; 
  assign _special_entry_data_0_T={refill_ppn,io_ptw_resp_bits_pte_u,newEntry_g,io_ptw_resp_bits_ae,newEntry_sw,newEntry_sx,newEntry_sr,prot_w,special_entry_data_0_lo}; 
  assign _GEN_32=invalidate_refill ? 1'h0:1'h1; 
  assign _T_2=io_ptw_resp_bits_level<2'h2; 
  assign _T_3=r_superpage_repl_addr==2'h0; 
  assign _GEN_35=_T_3 ? _GEN_32:superpage_entries_0_valid_0; 
  assign _T_4=r_superpage_repl_addr==2'h1; 
  assign _GEN_39=_T_4 ? _GEN_32:superpage_entries_1_valid_0; 
  assign _T_5=r_superpage_repl_addr==2'h2; 
  assign _GEN_43=_T_5 ? _GEN_32:superpage_entries_2_valid_0; 
  assign _T_6=r_superpage_repl_addr==2'h3; 
  assign _GEN_47=_T_6 ? _GEN_32:superpage_entries_3_valid_0; 
  assign waddr=r_sectored_hit ? r_sectored_hit_addr:r_sectored_repl_addr; 
  assign _T_7=waddr==3'h0; 
  assign _GEN_49=r_sectored_hit ? sectored_entries_0_0_valid_0:1'h0; 
  assign _GEN_50=r_sectored_hit ? sectored_entries_0_0_valid_1:1'h0; 
  assign _GEN_51=r_sectored_hit ? sectored_entries_0_0_valid_2:1'h0; 
  assign _GEN_52=r_sectored_hit ? sectored_entries_0_0_valid_3:1'h0; 
  assign idx=r_refill_tag[1:0]; 
  assign _GEN_921=2'h0==idx; 
  assign _GEN_53=_GEN_921|_GEN_49; 
  assign _GEN_922=2'h1==idx; 
  assign _GEN_54=_GEN_922|_GEN_50; 
  assign _GEN_923=2'h2==idx; 
  assign _GEN_55=_GEN_923|_GEN_51; 
  assign _GEN_924=2'h3==idx; 
  assign _GEN_56=_GEN_924|_GEN_52; 
  assign _GEN_61=invalidate_refill ? 1'h0:_GEN_53; 
  assign _GEN_62=invalidate_refill ? 1'h0:_GEN_54; 
  assign _GEN_63=invalidate_refill ? 1'h0:_GEN_55; 
  assign _GEN_64=invalidate_refill ? 1'h0:_GEN_56; 
  assign _GEN_65=_T_7 ? _GEN_61:sectored_entries_0_0_valid_0; 
  assign _GEN_66=_T_7 ? _GEN_62:sectored_entries_0_0_valid_1; 
  assign _GEN_67=_T_7 ? _GEN_63:sectored_entries_0_0_valid_2; 
  assign _GEN_68=_T_7 ? _GEN_64:sectored_entries_0_0_valid_3; 
  assign _T_9=waddr==3'h1; 
  assign _GEN_75=r_sectored_hit ? sectored_entries_0_1_valid_0:1'h0; 
  assign _GEN_76=r_sectored_hit ? sectored_entries_0_1_valid_1:1'h0; 
  assign _GEN_77=r_sectored_hit ? sectored_entries_0_1_valid_2:1'h0; 
  assign _GEN_78=r_sectored_hit ? sectored_entries_0_1_valid_3:1'h0; 
  assign _GEN_79=_GEN_921|_GEN_75; 
  assign _GEN_80=_GEN_922|_GEN_76; 
  assign _GEN_81=_GEN_923|_GEN_77; 
  assign _GEN_82=_GEN_924|_GEN_78; 
  assign _GEN_87=invalidate_refill ? 1'h0:_GEN_79; 
  assign _GEN_88=invalidate_refill ? 1'h0:_GEN_80; 
  assign _GEN_89=invalidate_refill ? 1'h0:_GEN_81; 
  assign _GEN_90=invalidate_refill ? 1'h0:_GEN_82; 
  assign _GEN_91=_T_9 ? _GEN_87:sectored_entries_0_1_valid_0; 
  assign _GEN_92=_T_9 ? _GEN_88:sectored_entries_0_1_valid_1; 
  assign _GEN_93=_T_9 ? _GEN_89:sectored_entries_0_1_valid_2; 
  assign _GEN_94=_T_9 ? _GEN_90:sectored_entries_0_1_valid_3; 
  assign _T_11=waddr==3'h2; 
  assign _GEN_101=r_sectored_hit ? sectored_entries_0_2_valid_0:1'h0; 
  assign _GEN_102=r_sectored_hit ? sectored_entries_0_2_valid_1:1'h0; 
  assign _GEN_103=r_sectored_hit ? sectored_entries_0_2_valid_2:1'h0; 
  assign _GEN_104=r_sectored_hit ? sectored_entries_0_2_valid_3:1'h0; 
  assign _GEN_105=_GEN_921|_GEN_101; 
  assign _GEN_106=_GEN_922|_GEN_102; 
  assign _GEN_107=_GEN_923|_GEN_103; 
  assign _GEN_108=_GEN_924|_GEN_104; 
  assign _GEN_113=invalidate_refill ? 1'h0:_GEN_105; 
  assign _GEN_114=invalidate_refill ? 1'h0:_GEN_106; 
  assign _GEN_115=invalidate_refill ? 1'h0:_GEN_107; 
  assign _GEN_116=invalidate_refill ? 1'h0:_GEN_108; 
  assign _GEN_117=_T_11 ? _GEN_113:sectored_entries_0_2_valid_0; 
  assign _GEN_118=_T_11 ? _GEN_114:sectored_entries_0_2_valid_1; 
  assign _GEN_119=_T_11 ? _GEN_115:sectored_entries_0_2_valid_2; 
  assign _GEN_120=_T_11 ? _GEN_116:sectored_entries_0_2_valid_3; 
  assign _T_13=waddr==3'h3; 
  assign _GEN_127=r_sectored_hit ? sectored_entries_0_3_valid_0:1'h0; 
  assign _GEN_128=r_sectored_hit ? sectored_entries_0_3_valid_1:1'h0; 
  assign _GEN_129=r_sectored_hit ? sectored_entries_0_3_valid_2:1'h0; 
  assign _GEN_130=r_sectored_hit ? sectored_entries_0_3_valid_3:1'h0; 
  assign _GEN_131=_GEN_921|_GEN_127; 
  assign _GEN_132=_GEN_922|_GEN_128; 
  assign _GEN_133=_GEN_923|_GEN_129; 
  assign _GEN_134=_GEN_924|_GEN_130; 
  assign _GEN_139=invalidate_refill ? 1'h0:_GEN_131; 
  assign _GEN_140=invalidate_refill ? 1'h0:_GEN_132; 
  assign _GEN_141=invalidate_refill ? 1'h0:_GEN_133; 
  assign _GEN_142=invalidate_refill ? 1'h0:_GEN_134; 
  assign _GEN_143=_T_13 ? _GEN_139:sectored_entries_0_3_valid_0; 
  assign _GEN_144=_T_13 ? _GEN_140:sectored_entries_0_3_valid_1; 
  assign _GEN_145=_T_13 ? _GEN_141:sectored_entries_0_3_valid_2; 
  assign _GEN_146=_T_13 ? _GEN_142:sectored_entries_0_3_valid_3; 
  assign _T_15=waddr==3'h4; 
  assign _GEN_153=r_sectored_hit ? sectored_entries_0_4_valid_0:1'h0; 
  assign _GEN_154=r_sectored_hit ? sectored_entries_0_4_valid_1:1'h0; 
  assign _GEN_155=r_sectored_hit ? sectored_entries_0_4_valid_2:1'h0; 
  assign _GEN_156=r_sectored_hit ? sectored_entries_0_4_valid_3:1'h0; 
  assign _GEN_157=_GEN_921|_GEN_153; 
  assign _GEN_158=_GEN_922|_GEN_154; 
  assign _GEN_159=_GEN_923|_GEN_155; 
  assign _GEN_160=_GEN_924|_GEN_156; 
  assign _GEN_165=invalidate_refill ? 1'h0:_GEN_157; 
  assign _GEN_166=invalidate_refill ? 1'h0:_GEN_158; 
  assign _GEN_167=invalidate_refill ? 1'h0:_GEN_159; 
  assign _GEN_168=invalidate_refill ? 1'h0:_GEN_160; 
  assign _GEN_169=_T_15 ? _GEN_165:sectored_entries_0_4_valid_0; 
  assign _GEN_170=_T_15 ? _GEN_166:sectored_entries_0_4_valid_1; 
  assign _GEN_171=_T_15 ? _GEN_167:sectored_entries_0_4_valid_2; 
  assign _GEN_172=_T_15 ? _GEN_168:sectored_entries_0_4_valid_3; 
  assign _T_17=waddr==3'h5; 
  assign _GEN_179=r_sectored_hit ? sectored_entries_0_5_valid_0:1'h0; 
  assign _GEN_180=r_sectored_hit ? sectored_entries_0_5_valid_1:1'h0; 
  assign _GEN_181=r_sectored_hit ? sectored_entries_0_5_valid_2:1'h0; 
  assign _GEN_182=r_sectored_hit ? sectored_entries_0_5_valid_3:1'h0; 
  assign _GEN_183=_GEN_921|_GEN_179; 
  assign _GEN_184=_GEN_922|_GEN_180; 
  assign _GEN_185=_GEN_923|_GEN_181; 
  assign _GEN_186=_GEN_924|_GEN_182; 
  assign _GEN_191=invalidate_refill ? 1'h0:_GEN_183; 
  assign _GEN_192=invalidate_refill ? 1'h0:_GEN_184; 
  assign _GEN_193=invalidate_refill ? 1'h0:_GEN_185; 
  assign _GEN_194=invalidate_refill ? 1'h0:_GEN_186; 
  assign _GEN_195=_T_17 ? _GEN_191:sectored_entries_0_5_valid_0; 
  assign _GEN_196=_T_17 ? _GEN_192:sectored_entries_0_5_valid_1; 
  assign _GEN_197=_T_17 ? _GEN_193:sectored_entries_0_5_valid_2; 
  assign _GEN_198=_T_17 ? _GEN_194:sectored_entries_0_5_valid_3; 
  assign _T_19=waddr==3'h6; 
  assign _GEN_205=r_sectored_hit ? sectored_entries_0_6_valid_0:1'h0; 
  assign _GEN_206=r_sectored_hit ? sectored_entries_0_6_valid_1:1'h0; 
  assign _GEN_207=r_sectored_hit ? sectored_entries_0_6_valid_2:1'h0; 
  assign _GEN_208=r_sectored_hit ? sectored_entries_0_6_valid_3:1'h0; 
  assign _GEN_209=_GEN_921|_GEN_205; 
  assign _GEN_210=_GEN_922|_GEN_206; 
  assign _GEN_211=_GEN_923|_GEN_207; 
  assign _GEN_212=_GEN_924|_GEN_208; 
  assign _GEN_217=invalidate_refill ? 1'h0:_GEN_209; 
  assign _GEN_218=invalidate_refill ? 1'h0:_GEN_210; 
  assign _GEN_219=invalidate_refill ? 1'h0:_GEN_211; 
  assign _GEN_220=invalidate_refill ? 1'h0:_GEN_212; 
  assign _GEN_221=_T_19 ? _GEN_217:sectored_entries_0_6_valid_0; 
  assign _GEN_222=_T_19 ? _GEN_218:sectored_entries_0_6_valid_1; 
  assign _GEN_223=_T_19 ? _GEN_219:sectored_entries_0_6_valid_2; 
  assign _GEN_224=_T_19 ? _GEN_220:sectored_entries_0_6_valid_3; 
  assign _T_21=waddr==3'h7; 
  assign _GEN_231=r_sectored_hit ? sectored_entries_0_7_valid_0:1'h0; 
  assign _GEN_232=r_sectored_hit ? sectored_entries_0_7_valid_1:1'h0; 
  assign _GEN_233=r_sectored_hit ? sectored_entries_0_7_valid_2:1'h0; 
  assign _GEN_234=r_sectored_hit ? sectored_entries_0_7_valid_3:1'h0; 
  assign _GEN_235=_GEN_921|_GEN_231; 
  assign _GEN_236=_GEN_922|_GEN_232; 
  assign _GEN_237=_GEN_923|_GEN_233; 
  assign _GEN_238=_GEN_924|_GEN_234; 
  assign _GEN_243=invalidate_refill ? 1'h0:_GEN_235; 
  assign _GEN_244=invalidate_refill ? 1'h0:_GEN_236; 
  assign _GEN_245=invalidate_refill ? 1'h0:_GEN_237; 
  assign _GEN_246=invalidate_refill ? 1'h0:_GEN_238; 
  assign _GEN_247=_T_21 ? _GEN_243:sectored_entries_0_7_valid_0; 
  assign _GEN_248=_T_21 ? _GEN_244:sectored_entries_0_7_valid_1; 
  assign _GEN_249=_T_21 ? _GEN_245:sectored_entries_0_7_valid_2; 
  assign _GEN_250=_T_21 ? _GEN_246:sectored_entries_0_7_valid_3; 
  assign _GEN_259=_T_2 ? _GEN_35:superpage_entries_0_valid_0; 
  assign _GEN_263=_T_2 ? _GEN_39:superpage_entries_1_valid_0; 
  assign _GEN_267=_T_2 ? _GEN_43:superpage_entries_2_valid_0; 
  assign _GEN_271=_T_2 ? _GEN_47:superpage_entries_3_valid_0; 
  assign _GEN_273=_T_2 ? sectored_entries_0_0_valid_0:_GEN_65; 
  assign _GEN_274=_T_2 ? sectored_entries_0_0_valid_1:_GEN_66; 
  assign _GEN_275=_T_2 ? sectored_entries_0_0_valid_2:_GEN_67; 
  assign _GEN_276=_T_2 ? sectored_entries_0_0_valid_3:_GEN_68; 
  assign _GEN_283=_T_2 ? sectored_entries_0_1_valid_0:_GEN_91; 
  assign _GEN_284=_T_2 ? sectored_entries_0_1_valid_1:_GEN_92; 
  assign _GEN_285=_T_2 ? sectored_entries_0_1_valid_2:_GEN_93; 
  assign _GEN_286=_T_2 ? sectored_entries_0_1_valid_3:_GEN_94; 
  assign _GEN_293=_T_2 ? sectored_entries_0_2_valid_0:_GEN_117; 
  assign _GEN_294=_T_2 ? sectored_entries_0_2_valid_1:_GEN_118; 
  assign _GEN_295=_T_2 ? sectored_entries_0_2_valid_2:_GEN_119; 
  assign _GEN_296=_T_2 ? sectored_entries_0_2_valid_3:_GEN_120; 
  assign _GEN_303=_T_2 ? sectored_entries_0_3_valid_0:_GEN_143; 
  assign _GEN_304=_T_2 ? sectored_entries_0_3_valid_1:_GEN_144; 
  assign _GEN_305=_T_2 ? sectored_entries_0_3_valid_2:_GEN_145; 
  assign _GEN_306=_T_2 ? sectored_entries_0_3_valid_3:_GEN_146; 
  assign _GEN_313=_T_2 ? sectored_entries_0_4_valid_0:_GEN_169; 
  assign _GEN_314=_T_2 ? sectored_entries_0_4_valid_1:_GEN_170; 
  assign _GEN_315=_T_2 ? sectored_entries_0_4_valid_2:_GEN_171; 
  assign _GEN_316=_T_2 ? sectored_entries_0_4_valid_3:_GEN_172; 
  assign _GEN_323=_T_2 ? sectored_entries_0_5_valid_0:_GEN_195; 
  assign _GEN_324=_T_2 ? sectored_entries_0_5_valid_1:_GEN_196; 
  assign _GEN_325=_T_2 ? sectored_entries_0_5_valid_2:_GEN_197; 
  assign _GEN_326=_T_2 ? sectored_entries_0_5_valid_3:_GEN_198; 
  assign _GEN_333=_T_2 ? sectored_entries_0_6_valid_0:_GEN_221; 
  assign _GEN_334=_T_2 ? sectored_entries_0_6_valid_1:_GEN_222; 
  assign _GEN_335=_T_2 ? sectored_entries_0_6_valid_2:_GEN_223; 
  assign _GEN_336=_T_2 ? sectored_entries_0_6_valid_3:_GEN_224; 
  assign _GEN_343=_T_2 ? sectored_entries_0_7_valid_0:_GEN_247; 
  assign _GEN_344=_T_2 ? sectored_entries_0_7_valid_1:_GEN_248; 
  assign _GEN_345=_T_2 ? sectored_entries_0_7_valid_2:_GEN_249; 
  assign _GEN_346=_T_2 ? sectored_entries_0_7_valid_3:_GEN_250; 
  assign _GEN_355=io_ptw_resp_bits_homogeneous ? special_entry_valid_0:_GEN_32; 
  assign _GEN_359=io_ptw_resp_bits_homogeneous ? _GEN_259:superpage_entries_0_valid_0; 
  assign _GEN_363=io_ptw_resp_bits_homogeneous ? _GEN_263:superpage_entries_1_valid_0; 
  assign _GEN_367=io_ptw_resp_bits_homogeneous ? _GEN_267:superpage_entries_2_valid_0; 
  assign _GEN_371=io_ptw_resp_bits_homogeneous ? _GEN_271:superpage_entries_3_valid_0; 
  assign _GEN_373=io_ptw_resp_bits_homogeneous ? _GEN_273:sectored_entries_0_0_valid_0; 
  assign _GEN_374=io_ptw_resp_bits_homogeneous ? _GEN_274:sectored_entries_0_0_valid_1; 
  assign _GEN_375=io_ptw_resp_bits_homogeneous ? _GEN_275:sectored_entries_0_0_valid_2; 
  assign _GEN_376=io_ptw_resp_bits_homogeneous ? _GEN_276:sectored_entries_0_0_valid_3; 
  assign _GEN_383=io_ptw_resp_bits_homogeneous ? _GEN_283:sectored_entries_0_1_valid_0; 
  assign _GEN_384=io_ptw_resp_bits_homogeneous ? _GEN_284:sectored_entries_0_1_valid_1; 
  assign _GEN_385=io_ptw_resp_bits_homogeneous ? _GEN_285:sectored_entries_0_1_valid_2; 
  assign _GEN_386=io_ptw_resp_bits_homogeneous ? _GEN_286:sectored_entries_0_1_valid_3; 
  assign _GEN_393=io_ptw_resp_bits_homogeneous ? _GEN_293:sectored_entries_0_2_valid_0; 
  assign _GEN_394=io_ptw_resp_bits_homogeneous ? _GEN_294:sectored_entries_0_2_valid_1; 
  assign _GEN_395=io_ptw_resp_bits_homogeneous ? _GEN_295:sectored_entries_0_2_valid_2; 
  assign _GEN_396=io_ptw_resp_bits_homogeneous ? _GEN_296:sectored_entries_0_2_valid_3; 
  assign _GEN_403=io_ptw_resp_bits_homogeneous ? _GEN_303:sectored_entries_0_3_valid_0; 
  assign _GEN_404=io_ptw_resp_bits_homogeneous ? _GEN_304:sectored_entries_0_3_valid_1; 
  assign _GEN_405=io_ptw_resp_bits_homogeneous ? _GEN_305:sectored_entries_0_3_valid_2; 
  assign _GEN_406=io_ptw_resp_bits_homogeneous ? _GEN_306:sectored_entries_0_3_valid_3; 
  assign _GEN_413=io_ptw_resp_bits_homogeneous ? _GEN_313:sectored_entries_0_4_valid_0; 
  assign _GEN_414=io_ptw_resp_bits_homogeneous ? _GEN_314:sectored_entries_0_4_valid_1; 
  assign _GEN_415=io_ptw_resp_bits_homogeneous ? _GEN_315:sectored_entries_0_4_valid_2; 
  assign _GEN_416=io_ptw_resp_bits_homogeneous ? _GEN_316:sectored_entries_0_4_valid_3; 
  assign _GEN_423=io_ptw_resp_bits_homogeneous ? _GEN_323:sectored_entries_0_5_valid_0; 
  assign _GEN_424=io_ptw_resp_bits_homogeneous ? _GEN_324:sectored_entries_0_5_valid_1; 
  assign _GEN_425=io_ptw_resp_bits_homogeneous ? _GEN_325:sectored_entries_0_5_valid_2; 
  assign _GEN_426=io_ptw_resp_bits_homogeneous ? _GEN_326:sectored_entries_0_5_valid_3; 
  assign _GEN_433=io_ptw_resp_bits_homogeneous ? _GEN_333:sectored_entries_0_6_valid_0; 
  assign _GEN_434=io_ptw_resp_bits_homogeneous ? _GEN_334:sectored_entries_0_6_valid_1; 
  assign _GEN_435=io_ptw_resp_bits_homogeneous ? _GEN_335:sectored_entries_0_6_valid_2; 
  assign _GEN_436=io_ptw_resp_bits_homogeneous ? _GEN_336:sectored_entries_0_6_valid_3; 
  assign _GEN_443=io_ptw_resp_bits_homogeneous ? _GEN_343:sectored_entries_0_7_valid_0; 
  assign _GEN_444=io_ptw_resp_bits_homogeneous ? _GEN_344:sectored_entries_0_7_valid_1; 
  assign _GEN_445=io_ptw_resp_bits_homogeneous ? _GEN_345:sectored_entries_0_7_valid_2; 
  assign _GEN_446=io_ptw_resp_bits_homogeneous ? _GEN_346:sectored_entries_0_7_valid_3; 
  assign _GEN_455=io_ptw_resp_valid ? _GEN_355:special_entry_valid_0; 
  assign _GEN_459=io_ptw_resp_valid ? _GEN_359:superpage_entries_0_valid_0; 
  assign _GEN_463=io_ptw_resp_valid ? _GEN_363:superpage_entries_1_valid_0; 
  assign _GEN_467=io_ptw_resp_valid ? _GEN_367:superpage_entries_2_valid_0; 
  assign _GEN_471=io_ptw_resp_valid ? _GEN_371:superpage_entries_3_valid_0; 
  assign _GEN_473=io_ptw_resp_valid ? _GEN_373:sectored_entries_0_0_valid_0; 
  assign _GEN_474=io_ptw_resp_valid ? _GEN_374:sectored_entries_0_0_valid_1; 
  assign _GEN_475=io_ptw_resp_valid ? _GEN_375:sectored_entries_0_0_valid_2; 
  assign _GEN_476=io_ptw_resp_valid ? _GEN_376:sectored_entries_0_0_valid_3; 
  assign _GEN_483=io_ptw_resp_valid ? _GEN_383:sectored_entries_0_1_valid_0; 
  assign _GEN_484=io_ptw_resp_valid ? _GEN_384:sectored_entries_0_1_valid_1; 
  assign _GEN_485=io_ptw_resp_valid ? _GEN_385:sectored_entries_0_1_valid_2; 
  assign _GEN_486=io_ptw_resp_valid ? _GEN_386:sectored_entries_0_1_valid_3; 
  assign _GEN_493=io_ptw_resp_valid ? _GEN_393:sectored_entries_0_2_valid_0; 
  assign _GEN_494=io_ptw_resp_valid ? _GEN_394:sectored_entries_0_2_valid_1; 
  assign _GEN_495=io_ptw_resp_valid ? _GEN_395:sectored_entries_0_2_valid_2; 
  assign _GEN_496=io_ptw_resp_valid ? _GEN_396:sectored_entries_0_2_valid_3; 
  assign _GEN_503=io_ptw_resp_valid ? _GEN_403:sectored_entries_0_3_valid_0; 
  assign _GEN_504=io_ptw_resp_valid ? _GEN_404:sectored_entries_0_3_valid_1; 
  assign _GEN_505=io_ptw_resp_valid ? _GEN_405:sectored_entries_0_3_valid_2; 
  assign _GEN_506=io_ptw_resp_valid ? _GEN_406:sectored_entries_0_3_valid_3; 
  assign _GEN_513=io_ptw_resp_valid ? _GEN_413:sectored_entries_0_4_valid_0; 
  assign _GEN_514=io_ptw_resp_valid ? _GEN_414:sectored_entries_0_4_valid_1; 
  assign _GEN_515=io_ptw_resp_valid ? _GEN_415:sectored_entries_0_4_valid_2; 
  assign _GEN_516=io_ptw_resp_valid ? _GEN_416:sectored_entries_0_4_valid_3; 
  assign _GEN_523=io_ptw_resp_valid ? _GEN_423:sectored_entries_0_5_valid_0; 
  assign _GEN_524=io_ptw_resp_valid ? _GEN_424:sectored_entries_0_5_valid_1; 
  assign _GEN_525=io_ptw_resp_valid ? _GEN_425:sectored_entries_0_5_valid_2; 
  assign _GEN_526=io_ptw_resp_valid ? _GEN_426:sectored_entries_0_5_valid_3; 
  assign _GEN_533=io_ptw_resp_valid ? _GEN_433:sectored_entries_0_6_valid_0; 
  assign _GEN_534=io_ptw_resp_valid ? _GEN_434:sectored_entries_0_6_valid_1; 
  assign _GEN_535=io_ptw_resp_valid ? _GEN_435:sectored_entries_0_6_valid_2; 
  assign _GEN_536=io_ptw_resp_valid ? _GEN_436:sectored_entries_0_6_valid_3; 
  assign _GEN_543=io_ptw_resp_valid ? _GEN_443:sectored_entries_0_7_valid_0; 
  assign _GEN_544=io_ptw_resp_valid ? _GEN_444:sectored_entries_0_7_valid_1; 
  assign _GEN_545=io_ptw_resp_valid ? _GEN_445:sectored_entries_0_7_valid_2; 
  assign _GEN_546=io_ptw_resp_valid ? _GEN_446:sectored_entries_0_7_valid_3; 
  assign _GEN_554=2'h1==hitsVec_idx ? sectored_entries_0_0_data_1:sectored_entries_0_0_data_0; 
  assign _GEN_555=2'h2==hitsVec_idx ? sectored_entries_0_0_data_2:_GEN_554; 
  assign _GEN_556=2'h3==hitsVec_idx ? sectored_entries_0_0_data_3:_GEN_555; 
  assign _GEN_558=2'h1==hitsVec_idx ? sectored_entries_0_1_data_1:sectored_entries_0_1_data_0; 
  assign _GEN_559=2'h2==hitsVec_idx ? sectored_entries_0_1_data_2:_GEN_558; 
  assign _GEN_560=2'h3==hitsVec_idx ? sectored_entries_0_1_data_3:_GEN_559; 
  assign _GEN_562=2'h1==hitsVec_idx ? sectored_entries_0_2_data_1:sectored_entries_0_2_data_0; 
  assign _GEN_563=2'h2==hitsVec_idx ? sectored_entries_0_2_data_2:_GEN_562; 
  assign _GEN_564=2'h3==hitsVec_idx ? sectored_entries_0_2_data_3:_GEN_563; 
  assign _GEN_566=2'h1==hitsVec_idx ? sectored_entries_0_3_data_1:sectored_entries_0_3_data_0; 
  assign _GEN_567=2'h2==hitsVec_idx ? sectored_entries_0_3_data_2:_GEN_566; 
  assign _GEN_568=2'h3==hitsVec_idx ? sectored_entries_0_3_data_3:_GEN_567; 
  assign _GEN_570=2'h1==hitsVec_idx ? sectored_entries_0_4_data_1:sectored_entries_0_4_data_0; 
  assign _GEN_571=2'h2==hitsVec_idx ? sectored_entries_0_4_data_2:_GEN_570; 
  assign _GEN_572=2'h3==hitsVec_idx ? sectored_entries_0_4_data_3:_GEN_571; 
  assign _GEN_574=2'h1==hitsVec_idx ? sectored_entries_0_5_data_1:sectored_entries_0_5_data_0; 
  assign _GEN_575=2'h2==hitsVec_idx ? sectored_entries_0_5_data_2:_GEN_574; 
  assign _GEN_576=2'h3==hitsVec_idx ? sectored_entries_0_5_data_3:_GEN_575; 
  assign _GEN_578=2'h1==hitsVec_idx ? sectored_entries_0_6_data_1:sectored_entries_0_6_data_0; 
  assign _GEN_579=2'h2==hitsVec_idx ? sectored_entries_0_6_data_2:_GEN_578; 
  assign _GEN_580=2'h3==hitsVec_idx ? sectored_entries_0_6_data_3:_GEN_579; 
  assign _GEN_582=2'h1==hitsVec_idx ? sectored_entries_0_7_data_1:sectored_entries_0_7_data_0; 
  assign _GEN_583=2'h2==hitsVec_idx ? sectored_entries_0_7_data_2:_GEN_582; 
  assign _GEN_584=2'h3==hitsVec_idx ? sectored_entries_0_7_data_3:_GEN_583; 
  assign ppn_hi=entries_barrier_8_io_y_ppn[19:18]; 
  assign _ppn_T_1=superpage_hits_ignore_1 ? vpn:27'h0; 
  assign _GEN_953={7'b0,entries_barrier_8_io_y_ppn}; 
  assign _ppn_T_2=_ppn_T_1|_GEN_953; 
  assign ppn_lo=_ppn_T_2[17:9]; 
  assign _ppn_T_4=vpn|_GEN_953; 
  assign ppn_lo_1=_ppn_T_4[8:0]; 
  assign _ppn_T_5={ppn_hi,ppn_lo,ppn_lo_1}; 
  assign ppn_hi_2=entries_barrier_9_io_y_ppn[19:18]; 
  assign _ppn_T_6=superpage_hits_ignore_4 ? vpn:27'h0; 
  assign _GEN_955={7'b0,entries_barrier_9_io_y_ppn}; 
  assign _ppn_T_7=_ppn_T_6|_GEN_955; 
  assign ppn_lo_2=_ppn_T_7[17:9]; 
  assign _ppn_T_9=vpn|_GEN_955; 
  assign ppn_lo_3=_ppn_T_9[8:0]; 
  assign _ppn_T_10={ppn_hi_2,ppn_lo_2,ppn_lo_3}; 
  assign ppn_hi_4=entries_barrier_10_io_y_ppn[19:18]; 
  assign _ppn_T_11=superpage_hits_ignore_7 ? vpn:27'h0; 
  assign _GEN_957={7'b0,entries_barrier_10_io_y_ppn}; 
  assign _ppn_T_12=_ppn_T_11|_GEN_957; 
  assign ppn_lo_4=_ppn_T_12[17:9]; 
  assign _ppn_T_14=vpn|_GEN_957; 
  assign ppn_lo_5=_ppn_T_14[8:0]; 
  assign _ppn_T_15={ppn_hi_4,ppn_lo_4,ppn_lo_5}; 
  assign ppn_hi_6=entries_barrier_11_io_y_ppn[19:18]; 
  assign _ppn_T_16=superpage_hits_ignore_10 ? vpn:27'h0; 
  assign _GEN_959={7'b0,entries_barrier_11_io_y_ppn}; 
  assign _ppn_T_17=_ppn_T_16|_GEN_959; 
  assign ppn_lo_6=_ppn_T_17[17:9]; 
  assign _ppn_T_19=vpn|_GEN_959; 
  assign ppn_lo_7=_ppn_T_19[8:0]; 
  assign _ppn_T_20={ppn_hi_6,ppn_lo_6,ppn_lo_7}; 
  assign ppn_hi_8=entries_barrier_12_io_y_ppn[19:18]; 
  assign _GEN_961={7'b0,entries_barrier_12_io_y_ppn}; 
  assign _ppn_T_22=_mpu_ppn_T_17|_GEN_961; 
  assign ppn_lo_8=_ppn_T_22[17:9]; 
  assign _ppn_T_24=_mpu_ppn_T_19|_GEN_961; 
  assign ppn_lo_9=_ppn_T_24[8:0]; 
  assign _ppn_T_25={ppn_hi_8,ppn_lo_8,ppn_lo_9}; 
  assign _ppn_T_27=hitsVec_0 ? entries_barrier_io_y_ppn:20'h0; 
  assign _ppn_T_28=hitsVec_1 ? entries_barrier_1_io_y_ppn:20'h0; 
  assign _ppn_T_29=hitsVec_2 ? entries_barrier_2_io_y_ppn:20'h0; 
  assign _ppn_T_30=hitsVec_3 ? entries_barrier_3_io_y_ppn:20'h0; 
  assign _ppn_T_31=hitsVec_4 ? entries_barrier_4_io_y_ppn:20'h0; 
  assign _ppn_T_32=hitsVec_5 ? entries_barrier_5_io_y_ppn:20'h0; 
  assign _ppn_T_33=hitsVec_6 ? entries_barrier_6_io_y_ppn:20'h0; 
  assign _ppn_T_34=hitsVec_7 ? entries_barrier_7_io_y_ppn:20'h0; 
  assign _ppn_T_35=hitsVec_8 ? _ppn_T_5:20'h0; 
  assign _ppn_T_36=hitsVec_9 ? _ppn_T_10:20'h0; 
  assign _ppn_T_37=hitsVec_10 ? _ppn_T_15:20'h0; 
  assign _ppn_T_38=hitsVec_11 ? _ppn_T_20:20'h0; 
  assign _ppn_T_39=hitsVec_12 ? _ppn_T_25:20'h0; 
  assign _ppn_T_40=hits_hi ? vpn[19:0]:20'h0; 
  assign _ppn_T_41=_ppn_T_27|_ppn_T_28; 
  assign _ppn_T_42=_ppn_T_41|_ppn_T_29; 
  assign _ppn_T_43=_ppn_T_42|_ppn_T_30; 
  assign _ppn_T_44=_ppn_T_43|_ppn_T_31; 
  assign _ppn_T_45=_ppn_T_44|_ppn_T_32; 
  assign _ppn_T_46=_ppn_T_45|_ppn_T_33; 
  assign _ppn_T_47=_ppn_T_46|_ppn_T_34; 
  assign _ppn_T_48=_ppn_T_47|_ppn_T_35; 
  assign _ppn_T_49=_ppn_T_48|_ppn_T_36; 
  assign _ppn_T_50=_ppn_T_49|_ppn_T_37; 
  assign _ppn_T_51=_ppn_T_50|_ppn_T_38; 
  assign _ppn_T_52=_ppn_T_51|_ppn_T_39; 
  assign ppn=_ppn_T_52|_ppn_T_40; 
  assign ptw_ae_array_lo={entries_barrier_5_io_y_ae,entries_barrier_4_io_y_ae,entries_barrier_3_io_y_ae,entries_barrier_2_io_y_ae,entries_barrier_1_io_y_ae,entries_barrier_io_y_ae}; 
  assign ptw_ae_array={1'h0,entries_barrier_12_io_y_ae,entries_barrier_11_io_y_ae,entries_barrier_10_io_y_ae,entries_barrier_9_io_y_ae,entries_barrier_8_io_y_ae,entries_barrier_7_io_y_ae,entries_barrier_6_io_y_ae,ptw_ae_array_lo}; 
  assign priv_rw_ok_lo={entries_barrier_5_io_y_u,entries_barrier_4_io_y_u,entries_barrier_3_io_y_u,entries_barrier_2_io_y_u,entries_barrier_1_io_y_u,entries_barrier_io_y_u}; 
  assign _priv_rw_ok_T_2={entries_barrier_12_io_y_u,entries_barrier_11_io_y_u,entries_barrier_10_io_y_u,entries_barrier_9_io_y_u,entries_barrier_8_io_y_u,entries_barrier_7_io_y_u,entries_barrier_6_io_y_u,priv_rw_ok_lo}; 
  assign priv_x_ok=priv_s ? ~_priv_rw_ok_T_2:_priv_rw_ok_T_2; 
  assign r_array_lo_1={entries_barrier_5_io_y_sx,entries_barrier_4_io_y_sx,entries_barrier_3_io_y_sx,entries_barrier_2_io_y_sx,entries_barrier_1_io_y_sx,entries_barrier_io_y_sx}; 
  assign _r_array_T_1={entries_barrier_12_io_y_sx,entries_barrier_11_io_y_sx,entries_barrier_10_io_y_sx,entries_barrier_9_io_y_sx,entries_barrier_8_io_y_sx,entries_barrier_7_io_y_sx,entries_barrier_6_io_y_sx,r_array_lo_1}; 
  assign x_array_lo_1=priv_x_ok&_r_array_T_1; 
  assign x_array={1'h1,x_array_lo_1}; 
  assign px_array_hi=prot_x ? 2'h3:2'h0; 
  assign px_array_lo={entries_barrier_5_io_y_px,entries_barrier_4_io_y_px,entries_barrier_3_io_y_px,entries_barrier_2_io_y_px,entries_barrier_1_io_y_px,entries_barrier_io_y_px}; 
  assign _px_array_T_1={px_array_hi,entries_barrier_11_io_y_px,entries_barrier_10_io_y_px,entries_barrier_9_io_y_px,entries_barrier_8_io_y_px,entries_barrier_7_io_y_px,entries_barrier_6_io_y_px,px_array_lo}; 
  assign px_array=_px_array_T_1&~ptw_ae_array; 
  assign c_array_hi=cacheable ? 2'h3:2'h0; 
  assign c_array_lo={entries_barrier_5_io_y_c,entries_barrier_4_io_y_c,entries_barrier_3_io_y_c,entries_barrier_2_io_y_c,entries_barrier_1_io_y_c,entries_barrier_io_y_c}; 
  assign c_array={c_array_hi,entries_barrier_11_io_y_c,entries_barrier_10_io_y_c,entries_barrier_9_io_y_c,entries_barrier_8_io_y_c,entries_barrier_7_io_y_c,entries_barrier_6_io_y_c,c_array_lo}; 
  assign bad_va_maskedVAddr=io_req_bits_vaddr&40'hc000000000; 
  assign _bad_va_T_1=bad_va_maskedVAddr==40'h0; 
  assign _bad_va_T_2=bad_va_maskedVAddr==40'hc000000000; 
  assign _bad_va_T_3=_bad_va_T_1|_bad_va_T_2; 
  assign bad_va=vm_enabled&~_bad_va_T_3; 
  assign _pf_inst_array_T=x_array|ptw_ae_array; 
  assign pf_inst_array=~_pf_inst_array_T; 
  assign tlb_hit=|real_hits; 
  assign _tlb_miss_T_1=vm_enabled&~bad_va; 
  assign tlb_miss=_tlb_miss_T_1&~tlb_hit; 
  assign _T_23=io_req_valid&vm_enabled; 
  assign _T_24=sector_hits_0|sector_hits_1; 
  assign _T_25=_T_24|sector_hits_2; 
  assign _T_26=_T_25|sector_hits_3; 
  assign _T_27=_T_26|sector_hits_4; 
  assign _T_28=_T_27|sector_hits_5; 
  assign _T_29=_T_28|sector_hits_6; 
  assign _T_30=_T_29|sector_hits_7; 
  assign _T_31={sector_hits_7,sector_hits_6,sector_hits_5,sector_hits_4,sector_hits_3,sector_hits_2,sector_hits_1,sector_hits_0}; 
  assign hi_1=_T_31[7:4]; 
  assign lo_1=_T_31[3:0]; 
  assign hi_2=|hi_1; 
  assign _T_32=hi_1|lo_1; 
  assign hi_3=_T_32[3:2]; 
  assign lo_2=_T_32[1:0]; 
  assign hi_4=|hi_3; 
  assign _T_33=hi_3|lo_2; 
  assign lo_3=_T_33[1]; 
  assign state_vec_0_touch_way_sized={hi_2,hi_4,lo_3}; 
  assign state_vec_0_hi_hi=~state_vec_0_touch_way_sized[2]; 
  assign state_vec_0_left_subtree_state=state_vec_0[5:3]; 
  assign state_vec_0_right_subtree_state=state_vec_0[2:0]; 
  assign state_vec_0_hi_hi_1=~state_vec_0_touch_way_sized[1]; 
  assign state_vec_0_left_subtree_state_1=state_vec_0_left_subtree_state[1]; 
  assign state_vec_0_right_subtree_state_1=state_vec_0_left_subtree_state[0]; 
  assign state_vec_0_hi_lo=state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_1:~state_vec_0_touch_way_sized[0]; 
  assign state_vec_0_lo=state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0]:state_vec_0_right_subtree_state_1; 
  assign _state_vec_0_T_7={state_vec_0_hi_hi_1,state_vec_0_hi_lo,state_vec_0_lo}; 
  assign state_vec_0_hi_lo_1=state_vec_0_hi_hi ? state_vec_0_left_subtree_state:_state_vec_0_T_7; 
  assign state_vec_0_left_subtree_state_2=state_vec_0_right_subtree_state[1]; 
  assign state_vec_0_right_subtree_state_2=state_vec_0_right_subtree_state[0]; 
  assign state_vec_0_hi_lo_2=state_vec_0_hi_hi_1 ? state_vec_0_left_subtree_state_2:~state_vec_0_touch_way_sized[0]; 
  assign state_vec_0_lo_1=state_vec_0_hi_hi_1 ? ~state_vec_0_touch_way_sized[0]:state_vec_0_right_subtree_state_2; 
  assign _state_vec_0_T_15={state_vec_0_hi_hi_1,state_vec_0_hi_lo_2,state_vec_0_lo_1}; 
  assign state_vec_0_lo_2=state_vec_0_hi_hi ? _state_vec_0_T_15:state_vec_0_right_subtree_state; 
  assign _state_vec_0_T_16={state_vec_0_hi_hi,state_vec_0_hi_lo_1,state_vec_0_lo_2}; 
  assign _T_35=superpage_hits_0|superpage_hits_1; 
  assign _T_36=_T_35|superpage_hits_2; 
  assign _T_37=_T_36|superpage_hits_3; 
  assign _T_38={superpage_hits_3,superpage_hits_2,superpage_hits_1,superpage_hits_0}; 
  assign hi_6=_T_38[3:2]; 
  assign lo_6=_T_38[1:0]; 
  assign hi_7=|hi_6; 
  assign _T_39=hi_6|lo_6; 
  assign lo_7=_T_39[1]; 
  assign state_reg_touch_way_sized={hi_7,lo_7}; 
  assign state_reg_hi_hi=~state_reg_touch_way_sized[1]; 
  assign state_reg_left_subtree_state=state_reg_1[1]; 
  assign state_reg_right_subtree_state=state_reg_1[0]; 
  assign state_reg_hi_lo=state_reg_hi_hi ? state_reg_left_subtree_state:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo=state_reg_hi_hi ? ~state_reg_touch_way_sized[0]:state_reg_right_subtree_state; 
  assign _state_reg_T_6={state_reg_hi_hi,state_reg_hi_lo,state_reg_lo}; 
  assign multipleHits_leftOne=real_hits[0]; 
  assign multipleHits_leftOne_1=real_hits[1]; 
  assign multipleHits_rightOne=real_hits[2]; 
  assign multipleHits_rightOne_1=multipleHits_leftOne_1|multipleHits_rightOne; 
  assign multipleHits_rightTwo=multipleHits_leftOne_1&multipleHits_rightOne; 
  assign multipleHits_leftOne_2=multipleHits_leftOne|multipleHits_rightOne_1; 
  assign _multipleHits_T_9=multipleHits_leftOne&multipleHits_rightOne_1; 
  assign multipleHits_leftTwo=multipleHits_rightTwo|_multipleHits_T_9; 
  assign multipleHits_leftOne_3=real_hits[3]; 
  assign multipleHits_leftOne_4=real_hits[4]; 
  assign multipleHits_rightOne_2=real_hits[5]; 
  assign multipleHits_rightOne_3=multipleHits_leftOne_4|multipleHits_rightOne_2; 
  assign multipleHits_rightTwo_1=multipleHits_leftOne_4&multipleHits_rightOne_2; 
  assign multipleHits_rightOne_4=multipleHits_leftOne_3|multipleHits_rightOne_3; 
  assign _multipleHits_T_18=multipleHits_leftOne_3&multipleHits_rightOne_3; 
  assign multipleHits_rightTwo_2=multipleHits_rightTwo_1|_multipleHits_T_18; 
  assign multipleHits_leftOne_5=multipleHits_leftOne_2|multipleHits_rightOne_4; 
  assign _multipleHits_T_19=multipleHits_leftTwo|multipleHits_rightTwo_2; 
  assign _multipleHits_T_20=multipleHits_leftOne_2&multipleHits_rightOne_4; 
  assign multipleHits_leftTwo_1=_multipleHits_T_19|_multipleHits_T_20; 
  assign multipleHits_leftOne_6=real_hits[6]; 
  assign multipleHits_leftOne_7=real_hits[7]; 
  assign multipleHits_rightOne_5=real_hits[8]; 
  assign multipleHits_rightOne_6=multipleHits_leftOne_7|multipleHits_rightOne_5; 
  assign multipleHits_rightTwo_3=multipleHits_leftOne_7&multipleHits_rightOne_5; 
  assign multipleHits_leftOne_8=multipleHits_leftOne_6|multipleHits_rightOne_6; 
  assign _multipleHits_T_30=multipleHits_leftOne_6&multipleHits_rightOne_6; 
  assign multipleHits_leftTwo_2=multipleHits_rightTwo_3|_multipleHits_T_30; 
  assign multipleHits_leftOne_9=real_hits[9]; 
  assign multipleHits_rightOne_7=real_hits[10]; 
  assign multipleHits_leftOne_10=multipleHits_leftOne_9|multipleHits_rightOne_7; 
  assign multipleHits_leftTwo_3=multipleHits_leftOne_9&multipleHits_rightOne_7; 
  assign multipleHits_leftOne_11=real_hits[11]; 
  assign multipleHits_rightOne_8=real_hits[12]; 
  assign multipleHits_rightOne_9=multipleHits_leftOne_11|multipleHits_rightOne_8; 
  assign multipleHits_rightTwo_4=multipleHits_leftOne_11&multipleHits_rightOne_8; 
  assign multipleHits_rightOne_10=multipleHits_leftOne_10|multipleHits_rightOne_9; 
  assign _multipleHits_T_42=multipleHits_leftTwo_3|multipleHits_rightTwo_4; 
  assign _multipleHits_T_43=multipleHits_leftOne_10&multipleHits_rightOne_9; 
  assign multipleHits_rightTwo_5=_multipleHits_T_42|_multipleHits_T_43; 
  assign multipleHits_rightOne_11=multipleHits_leftOne_8|multipleHits_rightOne_10; 
  assign _multipleHits_T_44=multipleHits_leftTwo_2|multipleHits_rightTwo_5; 
  assign _multipleHits_T_45=multipleHits_leftOne_8&multipleHits_rightOne_10; 
  assign multipleHits_rightTwo_6=_multipleHits_T_44|_multipleHits_T_45; 
  assign _multipleHits_T_47=multipleHits_leftTwo_1|multipleHits_rightTwo_6; 
  assign _multipleHits_T_48=multipleHits_leftOne_5&multipleHits_rightOne_11; 
  assign multipleHits=_multipleHits_T_47|_multipleHits_T_48; 
  assign _io_resp_pf_inst_T=pf_inst_array&hits; 
  assign _io_resp_pf_inst_T_1=|_io_resp_pf_inst_T; 
  assign _io_resp_ae_inst_T_1=~px_array&hits; 
  assign _io_resp_cacheable_T=c_array&hits; 
  assign _io_resp_miss_T=io_ptw_resp_valid|tlb_miss; 
  assign _T_41=io_req_ready&io_req_valid; 
  assign _T_42=_T_41&tlb_miss; 
  assign r_superpage_repl_addr_hi=state_reg_1[2]; 
  assign r_superpage_repl_addr_lo=r_superpage_repl_addr_hi ? state_reg_left_subtree_state:state_reg_right_subtree_state; 
  assign _r_superpage_repl_addr_T_2={r_superpage_repl_addr_hi,r_superpage_repl_addr_lo}; 
  assign r_superpage_repl_addr_valids={superpage_entries_3_valid_0,superpage_entries_2_valid_0,superpage_entries_1_valid_0,superpage_entries_0_valid_0}; 
  assign _r_superpage_repl_addr_T_3=&r_superpage_repl_addr_valids; 
  assign _r_superpage_repl_addr_T_5=~r_superpage_repl_addr_valids[0]; 
  assign _r_superpage_repl_addr_T_6=~r_superpage_repl_addr_valids[1]; 
  assign _r_superpage_repl_addr_T_7=~r_superpage_repl_addr_valids[2]; 
  assign r_sectored_repl_addr_hi=state_vec_0[6]; 
  assign r_sectored_repl_addr_hi_1=state_vec_0_left_subtree_state[2]; 
  assign r_sectored_repl_addr_lo=r_sectored_repl_addr_hi_1 ? state_vec_0_left_subtree_state_1:state_vec_0_right_subtree_state_1; 
  assign _r_sectored_repl_addr_T_2={r_sectored_repl_addr_hi_1,r_sectored_repl_addr_lo}; 
  assign r_sectored_repl_addr_hi_2=state_vec_0_right_subtree_state[2]; 
  assign r_sectored_repl_addr_lo_1=r_sectored_repl_addr_hi_2 ? state_vec_0_left_subtree_state_2:state_vec_0_right_subtree_state_2; 
  assign _r_sectored_repl_addr_T_5={r_sectored_repl_addr_hi_2,r_sectored_repl_addr_lo_1}; 
  assign r_sectored_repl_addr_lo_2=r_sectored_repl_addr_hi ? _r_sectored_repl_addr_T_2:_r_sectored_repl_addr_T_5; 
  assign _r_sectored_repl_addr_T_6={r_sectored_repl_addr_hi,r_sectored_repl_addr_lo_2}; 
  assign r_sectored_repl_addr_valids={_sector_hits_T_44,_sector_hits_T_38,_sector_hits_T_32,_sector_hits_T_26,_sector_hits_T_20,_sector_hits_T_14,_sector_hits_T_8,_sector_hits_T_2}; 
  assign _r_sectored_repl_addr_T_7=&r_sectored_repl_addr_valids; 
  assign _r_sectored_repl_addr_T_9=~r_sectored_repl_addr_valids[0]; 
  assign _r_sectored_repl_addr_T_10=~r_sectored_repl_addr_valids[1]; 
  assign _r_sectored_repl_addr_T_11=~r_sectored_repl_addr_valids[2]; 
  assign _r_sectored_repl_addr_T_12=~r_sectored_repl_addr_valids[3]; 
  assign _r_sectored_repl_addr_T_13=~r_sectored_repl_addr_valids[4]; 
  assign _r_sectored_repl_addr_T_14=~r_sectored_repl_addr_valids[5]; 
  assign _r_sectored_repl_addr_T_15=~r_sectored_repl_addr_valids[6]; 
  assign _T_44=state==2'h2; 
  assign _T_45=_T_44&io_sfence_valid; 
  assign _T_48=io_sfence_bits_addr[38:12]==vpn; 
  assign _T_49=~io_sfence_bits_rs1|_T_48; 
  assign _T_51=_T_49|reset; 
  assign _T_59=_sector_hits_T_3[26:18]==9'h0; 
  assign _GEN_617=sectored_entries_0_0_data_0[13] ? _GEN_473:1'h0; 
  assign _GEN_618=sectored_entries_0_0_data_1[13] ? _GEN_474:1'h0; 
  assign _GEN_619=sectored_entries_0_0_data_2[13] ? _GEN_475:1'h0; 
  assign _GEN_620=sectored_entries_0_0_data_3[13] ? _GEN_476:1'h0; 
  assign _GEN_621=io_sfence_bits_rs2&_GEN_617; 
  assign _GEN_622=io_sfence_bits_rs2&_GEN_618; 
  assign _GEN_623=io_sfence_bits_rs2&_GEN_619; 
  assign _GEN_624=io_sfence_bits_rs2&_GEN_620; 
  assign _T_198=_sector_hits_T_9[26:18]==9'h0; 
  assign _GEN_645=sectored_entries_0_1_data_0[13] ? _GEN_483:1'h0; 
  assign _GEN_646=sectored_entries_0_1_data_1[13] ? _GEN_484:1'h0; 
  assign _GEN_647=sectored_entries_0_1_data_2[13] ? _GEN_485:1'h0; 
  assign _GEN_648=sectored_entries_0_1_data_3[13] ? _GEN_486:1'h0; 
  assign _GEN_649=io_sfence_bits_rs2&_GEN_645; 
  assign _GEN_650=io_sfence_bits_rs2&_GEN_646; 
  assign _GEN_651=io_sfence_bits_rs2&_GEN_647; 
  assign _GEN_652=io_sfence_bits_rs2&_GEN_648; 
  assign _T_337=_sector_hits_T_15[26:18]==9'h0; 
  assign _GEN_673=sectored_entries_0_2_data_0[13] ? _GEN_493:1'h0; 
  assign _GEN_674=sectored_entries_0_2_data_1[13] ? _GEN_494:1'h0; 
  assign _GEN_675=sectored_entries_0_2_data_2[13] ? _GEN_495:1'h0; 
  assign _GEN_676=sectored_entries_0_2_data_3[13] ? _GEN_496:1'h0; 
  assign _GEN_677=io_sfence_bits_rs2&_GEN_673; 
  assign _GEN_678=io_sfence_bits_rs2&_GEN_674; 
  assign _GEN_679=io_sfence_bits_rs2&_GEN_675; 
  assign _GEN_680=io_sfence_bits_rs2&_GEN_676; 
  assign _T_476=_sector_hits_T_21[26:18]==9'h0; 
  assign _GEN_701=sectored_entries_0_3_data_0[13] ? _GEN_503:1'h0; 
  assign _GEN_702=sectored_entries_0_3_data_1[13] ? _GEN_504:1'h0; 
  assign _GEN_703=sectored_entries_0_3_data_2[13] ? _GEN_505:1'h0; 
  assign _GEN_704=sectored_entries_0_3_data_3[13] ? _GEN_506:1'h0; 
  assign _GEN_705=io_sfence_bits_rs2&_GEN_701; 
  assign _GEN_706=io_sfence_bits_rs2&_GEN_702; 
  assign _GEN_707=io_sfence_bits_rs2&_GEN_703; 
  assign _GEN_708=io_sfence_bits_rs2&_GEN_704; 
  assign _T_615=_sector_hits_T_27[26:18]==9'h0; 
  assign _GEN_729=sectored_entries_0_4_data_0[13] ? _GEN_513:1'h0; 
  assign _GEN_730=sectored_entries_0_4_data_1[13] ? _GEN_514:1'h0; 
  assign _GEN_731=sectored_entries_0_4_data_2[13] ? _GEN_515:1'h0; 
  assign _GEN_732=sectored_entries_0_4_data_3[13] ? _GEN_516:1'h0; 
  assign _GEN_733=io_sfence_bits_rs2&_GEN_729; 
  assign _GEN_734=io_sfence_bits_rs2&_GEN_730; 
  assign _GEN_735=io_sfence_bits_rs2&_GEN_731; 
  assign _GEN_736=io_sfence_bits_rs2&_GEN_732; 
  assign _T_754=_sector_hits_T_33[26:18]==9'h0; 
  assign _GEN_757=sectored_entries_0_5_data_0[13] ? _GEN_523:1'h0; 
  assign _GEN_758=sectored_entries_0_5_data_1[13] ? _GEN_524:1'h0; 
  assign _GEN_759=sectored_entries_0_5_data_2[13] ? _GEN_525:1'h0; 
  assign _GEN_760=sectored_entries_0_5_data_3[13] ? _GEN_526:1'h0; 
  assign _GEN_761=io_sfence_bits_rs2&_GEN_757; 
  assign _GEN_762=io_sfence_bits_rs2&_GEN_758; 
  assign _GEN_763=io_sfence_bits_rs2&_GEN_759; 
  assign _GEN_764=io_sfence_bits_rs2&_GEN_760; 
  assign _T_893=_sector_hits_T_39[26:18]==9'h0; 
  assign _GEN_785=sectored_entries_0_6_data_0[13] ? _GEN_533:1'h0; 
  assign _GEN_786=sectored_entries_0_6_data_1[13] ? _GEN_534:1'h0; 
  assign _GEN_787=sectored_entries_0_6_data_2[13] ? _GEN_535:1'h0; 
  assign _GEN_788=sectored_entries_0_6_data_3[13] ? _GEN_536:1'h0; 
  assign _GEN_789=io_sfence_bits_rs2&_GEN_785; 
  assign _GEN_790=io_sfence_bits_rs2&_GEN_786; 
  assign _GEN_791=io_sfence_bits_rs2&_GEN_787; 
  assign _GEN_792=io_sfence_bits_rs2&_GEN_788; 
  assign _T_1032=_sector_hits_T_45[26:18]==9'h0; 
  assign _GEN_813=sectored_entries_0_7_data_0[13] ? _GEN_543:1'h0; 
  assign _GEN_814=sectored_entries_0_7_data_1[13] ? _GEN_544:1'h0; 
  assign _GEN_815=sectored_entries_0_7_data_2[13] ? _GEN_545:1'h0; 
  assign _GEN_816=sectored_entries_0_7_data_3[13] ? _GEN_546:1'h0; 
  assign _GEN_817=io_sfence_bits_rs2&_GEN_813; 
  assign _GEN_818=io_sfence_bits_rs2&_GEN_814; 
  assign _GEN_819=io_sfence_bits_rs2&_GEN_815; 
  assign _GEN_820=io_sfence_bits_rs2&_GEN_816; 
  assign _GEN_826=superpage_entries_0_data_0[13] ? _GEN_459:1'h0; 
  assign _GEN_827=io_sfence_bits_rs2&_GEN_826; 
  assign _GEN_830=superpage_entries_1_data_0[13] ? _GEN_463:1'h0; 
  assign _GEN_831=io_sfence_bits_rs2&_GEN_830; 
  assign _GEN_834=superpage_entries_2_data_0[13] ? _GEN_467:1'h0; 
  assign _GEN_835=io_sfence_bits_rs2&_GEN_834; 
  assign _GEN_838=superpage_entries_3_data_0[13] ? _GEN_471:1'h0; 
  assign _GEN_839=io_sfence_bits_rs2&_GEN_838; 
  assign _GEN_842=special_entry_data_0[13] ? _GEN_455:1'h0; 
  assign _GEN_843=io_sfence_bits_rs2&_GEN_842; 
  assign _T_1326=multipleHits|reset; 
  assign io_req_ready=state==2'h0; 
  assign io_resp_miss=_io_resp_miss_T|multipleHits; 
  assign io_resp_paddr={ppn,mpu_physaddr_lo}; 
  assign io_resp_pf_inst=bad_va|_io_resp_pf_inst_T_1; 
  assign io_resp_ae_inst=|_io_resp_ae_inst_T_1; 
  assign io_resp_cacheable=|_io_resp_cacheable_T; 
  assign io_ptw_req_valid=state==2'h1; 
  assign io_ptw_req_bits_valid=~io_kill; 
  assign io_ptw_req_bits_bits_addr=r_refill_tag; 
  assign mpu_ppn_barrier_io_x_ppn=special_entry_data_0[34:15]; 
  assign mpu_ppn_barrier_io_x_u=special_entry_data_0[14]; 
  assign mpu_ppn_barrier_io_x_ae=special_entry_data_0[12]; 
  assign mpu_ppn_barrier_io_x_sw=special_entry_data_0[11]; 
  assign mpu_ppn_barrier_io_x_sx=special_entry_data_0[10]; 
  assign mpu_ppn_barrier_io_x_sr=special_entry_data_0[9]; 
  assign mpu_ppn_barrier_io_x_pw=special_entry_data_0[8]; 
  assign mpu_ppn_barrier_io_x_px=special_entry_data_0[7]; 
  assign mpu_ppn_barrier_io_x_pr=special_entry_data_0[6]; 
  assign mpu_ppn_barrier_io_x_ppp=special_entry_data_0[5]; 
  assign mpu_ppn_barrier_io_x_pal=special_entry_data_0[4]; 
  assign mpu_ppn_barrier_io_x_paa=special_entry_data_0[3]; 
  assign mpu_ppn_barrier_io_x_eff=special_entry_data_0[2]; 
  assign mpu_ppn_barrier_io_x_c=special_entry_data_0[1]; 
  assign pmp_io_prv=mpu_priv[1:0]; 
  assign pmp_io_pmp_0_cfg_l=io_ptw_pmp_0_cfg_l; 
  assign pmp_io_pmp_0_cfg_a=io_ptw_pmp_0_cfg_a; 
  assign pmp_io_pmp_0_cfg_x=io_ptw_pmp_0_cfg_x; 
  assign pmp_io_pmp_0_cfg_w=io_ptw_pmp_0_cfg_w; 
  assign pmp_io_pmp_0_cfg_r=io_ptw_pmp_0_cfg_r; 
  assign pmp_io_pmp_0_addr=io_ptw_pmp_0_addr; 
  assign pmp_io_pmp_0_mask=io_ptw_pmp_0_mask; 
  assign pmp_io_pmp_1_cfg_l=io_ptw_pmp_1_cfg_l; 
  assign pmp_io_pmp_1_cfg_a=io_ptw_pmp_1_cfg_a; 
  assign pmp_io_pmp_1_cfg_x=io_ptw_pmp_1_cfg_x; 
  assign pmp_io_pmp_1_cfg_w=io_ptw_pmp_1_cfg_w; 
  assign pmp_io_pmp_1_cfg_r=io_ptw_pmp_1_cfg_r; 
  assign pmp_io_pmp_1_addr=io_ptw_pmp_1_addr; 
  assign pmp_io_pmp_1_mask=io_ptw_pmp_1_mask; 
  assign pmp_io_pmp_2_cfg_l=io_ptw_pmp_2_cfg_l; 
  assign pmp_io_pmp_2_cfg_a=io_ptw_pmp_2_cfg_a; 
  assign pmp_io_pmp_2_cfg_x=io_ptw_pmp_2_cfg_x; 
  assign pmp_io_pmp_2_cfg_w=io_ptw_pmp_2_cfg_w; 
  assign pmp_io_pmp_2_cfg_r=io_ptw_pmp_2_cfg_r; 
  assign pmp_io_pmp_2_addr=io_ptw_pmp_2_addr; 
  assign pmp_io_pmp_2_mask=io_ptw_pmp_2_mask; 
  assign pmp_io_pmp_3_cfg_l=io_ptw_pmp_3_cfg_l; 
  assign pmp_io_pmp_3_cfg_a=io_ptw_pmp_3_cfg_a; 
  assign pmp_io_pmp_3_cfg_x=io_ptw_pmp_3_cfg_x; 
  assign pmp_io_pmp_3_cfg_w=io_ptw_pmp_3_cfg_w; 
  assign pmp_io_pmp_3_cfg_r=io_ptw_pmp_3_cfg_r; 
  assign pmp_io_pmp_3_addr=io_ptw_pmp_3_addr; 
  assign pmp_io_pmp_3_mask=io_ptw_pmp_3_mask; 
  assign pmp_io_pmp_4_cfg_l=io_ptw_pmp_4_cfg_l; 
  assign pmp_io_pmp_4_cfg_a=io_ptw_pmp_4_cfg_a; 
  assign pmp_io_pmp_4_cfg_x=io_ptw_pmp_4_cfg_x; 
  assign pmp_io_pmp_4_cfg_w=io_ptw_pmp_4_cfg_w; 
  assign pmp_io_pmp_4_cfg_r=io_ptw_pmp_4_cfg_r; 
  assign pmp_io_pmp_4_addr=io_ptw_pmp_4_addr; 
  assign pmp_io_pmp_4_mask=io_ptw_pmp_4_mask; 
  assign pmp_io_pmp_5_cfg_l=io_ptw_pmp_5_cfg_l; 
  assign pmp_io_pmp_5_cfg_a=io_ptw_pmp_5_cfg_a; 
  assign pmp_io_pmp_5_cfg_x=io_ptw_pmp_5_cfg_x; 
  assign pmp_io_pmp_5_cfg_w=io_ptw_pmp_5_cfg_w; 
  assign pmp_io_pmp_5_cfg_r=io_ptw_pmp_5_cfg_r; 
  assign pmp_io_pmp_5_addr=io_ptw_pmp_5_addr; 
  assign pmp_io_pmp_5_mask=io_ptw_pmp_5_mask; 
  assign pmp_io_pmp_6_cfg_l=io_ptw_pmp_6_cfg_l; 
  assign pmp_io_pmp_6_cfg_a=io_ptw_pmp_6_cfg_a; 
  assign pmp_io_pmp_6_cfg_x=io_ptw_pmp_6_cfg_x; 
  assign pmp_io_pmp_6_cfg_w=io_ptw_pmp_6_cfg_w; 
  assign pmp_io_pmp_6_cfg_r=io_ptw_pmp_6_cfg_r; 
  assign pmp_io_pmp_6_addr=io_ptw_pmp_6_addr; 
  assign pmp_io_pmp_6_mask=io_ptw_pmp_6_mask; 
  assign pmp_io_pmp_7_cfg_l=io_ptw_pmp_7_cfg_l; 
  assign pmp_io_pmp_7_cfg_a=io_ptw_pmp_7_cfg_a; 
  assign pmp_io_pmp_7_cfg_x=io_ptw_pmp_7_cfg_x; 
  assign pmp_io_pmp_7_cfg_w=io_ptw_pmp_7_cfg_w; 
  assign pmp_io_pmp_7_cfg_r=io_ptw_pmp_7_cfg_r; 
  assign pmp_io_pmp_7_addr=io_ptw_pmp_7_addr; 
  assign pmp_io_pmp_7_mask=io_ptw_pmp_7_mask; 
  assign pmp_io_addr=mpu_physaddr[31:0]; 
  assign entries_barrier_io_x_ppn=_GEN_556[34:15]; 
  assign entries_barrier_io_x_u=_GEN_556[14]; 
  assign entries_barrier_io_x_ae=_GEN_556[12]; 
  assign entries_barrier_io_x_sw=_GEN_556[11]; 
  assign entries_barrier_io_x_sx=_GEN_556[10]; 
  assign entries_barrier_io_x_sr=_GEN_556[9]; 
  assign entries_barrier_io_x_pw=_GEN_556[8]; 
  assign entries_barrier_io_x_px=_GEN_556[7]; 
  assign entries_barrier_io_x_pr=_GEN_556[6]; 
  assign entries_barrier_io_x_ppp=_GEN_556[5]; 
  assign entries_barrier_io_x_pal=_GEN_556[4]; 
  assign entries_barrier_io_x_paa=_GEN_556[3]; 
  assign entries_barrier_io_x_eff=_GEN_556[2]; 
  assign entries_barrier_io_x_c=_GEN_556[1]; 
  assign entries_barrier_1_io_x_ppn=_GEN_560[34:15]; 
  assign entries_barrier_1_io_x_u=_GEN_560[14]; 
  assign entries_barrier_1_io_x_ae=_GEN_560[12]; 
  assign entries_barrier_1_io_x_sw=_GEN_560[11]; 
  assign entries_barrier_1_io_x_sx=_GEN_560[10]; 
  assign entries_barrier_1_io_x_sr=_GEN_560[9]; 
  assign entries_barrier_1_io_x_pw=_GEN_560[8]; 
  assign entries_barrier_1_io_x_px=_GEN_560[7]; 
  assign entries_barrier_1_io_x_pr=_GEN_560[6]; 
  assign entries_barrier_1_io_x_ppp=_GEN_560[5]; 
  assign entries_barrier_1_io_x_pal=_GEN_560[4]; 
  assign entries_barrier_1_io_x_paa=_GEN_560[3]; 
  assign entries_barrier_1_io_x_eff=_GEN_560[2]; 
  assign entries_barrier_1_io_x_c=_GEN_560[1]; 
  assign entries_barrier_2_io_x_ppn=_GEN_564[34:15]; 
  assign entries_barrier_2_io_x_u=_GEN_564[14]; 
  assign entries_barrier_2_io_x_ae=_GEN_564[12]; 
  assign entries_barrier_2_io_x_sw=_GEN_564[11]; 
  assign entries_barrier_2_io_x_sx=_GEN_564[10]; 
  assign entries_barrier_2_io_x_sr=_GEN_564[9]; 
  assign entries_barrier_2_io_x_pw=_GEN_564[8]; 
  assign entries_barrier_2_io_x_px=_GEN_564[7]; 
  assign entries_barrier_2_io_x_pr=_GEN_564[6]; 
  assign entries_barrier_2_io_x_ppp=_GEN_564[5]; 
  assign entries_barrier_2_io_x_pal=_GEN_564[4]; 
  assign entries_barrier_2_io_x_paa=_GEN_564[3]; 
  assign entries_barrier_2_io_x_eff=_GEN_564[2]; 
  assign entries_barrier_2_io_x_c=_GEN_564[1]; 
  assign entries_barrier_3_io_x_ppn=_GEN_568[34:15]; 
  assign entries_barrier_3_io_x_u=_GEN_568[14]; 
  assign entries_barrier_3_io_x_ae=_GEN_568[12]; 
  assign entries_barrier_3_io_x_sw=_GEN_568[11]; 
  assign entries_barrier_3_io_x_sx=_GEN_568[10]; 
  assign entries_barrier_3_io_x_sr=_GEN_568[9]; 
  assign entries_barrier_3_io_x_pw=_GEN_568[8]; 
  assign entries_barrier_3_io_x_px=_GEN_568[7]; 
  assign entries_barrier_3_io_x_pr=_GEN_568[6]; 
  assign entries_barrier_3_io_x_ppp=_GEN_568[5]; 
  assign entries_barrier_3_io_x_pal=_GEN_568[4]; 
  assign entries_barrier_3_io_x_paa=_GEN_568[3]; 
  assign entries_barrier_3_io_x_eff=_GEN_568[2]; 
  assign entries_barrier_3_io_x_c=_GEN_568[1]; 
  assign entries_barrier_4_io_x_ppn=_GEN_572[34:15]; 
  assign entries_barrier_4_io_x_u=_GEN_572[14]; 
  assign entries_barrier_4_io_x_ae=_GEN_572[12]; 
  assign entries_barrier_4_io_x_sw=_GEN_572[11]; 
  assign entries_barrier_4_io_x_sx=_GEN_572[10]; 
  assign entries_barrier_4_io_x_sr=_GEN_572[9]; 
  assign entries_barrier_4_io_x_pw=_GEN_572[8]; 
  assign entries_barrier_4_io_x_px=_GEN_572[7]; 
  assign entries_barrier_4_io_x_pr=_GEN_572[6]; 
  assign entries_barrier_4_io_x_ppp=_GEN_572[5]; 
  assign entries_barrier_4_io_x_pal=_GEN_572[4]; 
  assign entries_barrier_4_io_x_paa=_GEN_572[3]; 
  assign entries_barrier_4_io_x_eff=_GEN_572[2]; 
  assign entries_barrier_4_io_x_c=_GEN_572[1]; 
  assign entries_barrier_5_io_x_ppn=_GEN_576[34:15]; 
  assign entries_barrier_5_io_x_u=_GEN_576[14]; 
  assign entries_barrier_5_io_x_ae=_GEN_576[12]; 
  assign entries_barrier_5_io_x_sw=_GEN_576[11]; 
  assign entries_barrier_5_io_x_sx=_GEN_576[10]; 
  assign entries_barrier_5_io_x_sr=_GEN_576[9]; 
  assign entries_barrier_5_io_x_pw=_GEN_576[8]; 
  assign entries_barrier_5_io_x_px=_GEN_576[7]; 
  assign entries_barrier_5_io_x_pr=_GEN_576[6]; 
  assign entries_barrier_5_io_x_ppp=_GEN_576[5]; 
  assign entries_barrier_5_io_x_pal=_GEN_576[4]; 
  assign entries_barrier_5_io_x_paa=_GEN_576[3]; 
  assign entries_barrier_5_io_x_eff=_GEN_576[2]; 
  assign entries_barrier_5_io_x_c=_GEN_576[1]; 
  assign entries_barrier_6_io_x_ppn=_GEN_580[34:15]; 
  assign entries_barrier_6_io_x_u=_GEN_580[14]; 
  assign entries_barrier_6_io_x_ae=_GEN_580[12]; 
  assign entries_barrier_6_io_x_sw=_GEN_580[11]; 
  assign entries_barrier_6_io_x_sx=_GEN_580[10]; 
  assign entries_barrier_6_io_x_sr=_GEN_580[9]; 
  assign entries_barrier_6_io_x_pw=_GEN_580[8]; 
  assign entries_barrier_6_io_x_px=_GEN_580[7]; 
  assign entries_barrier_6_io_x_pr=_GEN_580[6]; 
  assign entries_barrier_6_io_x_ppp=_GEN_580[5]; 
  assign entries_barrier_6_io_x_pal=_GEN_580[4]; 
  assign entries_barrier_6_io_x_paa=_GEN_580[3]; 
  assign entries_barrier_6_io_x_eff=_GEN_580[2]; 
  assign entries_barrier_6_io_x_c=_GEN_580[1]; 
  assign entries_barrier_7_io_x_ppn=_GEN_584[34:15]; 
  assign entries_barrier_7_io_x_u=_GEN_584[14]; 
  assign entries_barrier_7_io_x_ae=_GEN_584[12]; 
  assign entries_barrier_7_io_x_sw=_GEN_584[11]; 
  assign entries_barrier_7_io_x_sx=_GEN_584[10]; 
  assign entries_barrier_7_io_x_sr=_GEN_584[9]; 
  assign entries_barrier_7_io_x_pw=_GEN_584[8]; 
  assign entries_barrier_7_io_x_px=_GEN_584[7]; 
  assign entries_barrier_7_io_x_pr=_GEN_584[6]; 
  assign entries_barrier_7_io_x_ppp=_GEN_584[5]; 
  assign entries_barrier_7_io_x_pal=_GEN_584[4]; 
  assign entries_barrier_7_io_x_paa=_GEN_584[3]; 
  assign entries_barrier_7_io_x_eff=_GEN_584[2]; 
  assign entries_barrier_7_io_x_c=_GEN_584[1]; 
  assign entries_barrier_8_io_x_ppn=superpage_entries_0_data_0[34:15]; 
  assign entries_barrier_8_io_x_u=superpage_entries_0_data_0[14]; 
  assign entries_barrier_8_io_x_ae=superpage_entries_0_data_0[12]; 
  assign entries_barrier_8_io_x_sw=superpage_entries_0_data_0[11]; 
  assign entries_barrier_8_io_x_sx=superpage_entries_0_data_0[10]; 
  assign entries_barrier_8_io_x_sr=superpage_entries_0_data_0[9]; 
  assign entries_barrier_8_io_x_pw=superpage_entries_0_data_0[8]; 
  assign entries_barrier_8_io_x_px=superpage_entries_0_data_0[7]; 
  assign entries_barrier_8_io_x_pr=superpage_entries_0_data_0[6]; 
  assign entries_barrier_8_io_x_ppp=superpage_entries_0_data_0[5]; 
  assign entries_barrier_8_io_x_pal=superpage_entries_0_data_0[4]; 
  assign entries_barrier_8_io_x_paa=superpage_entries_0_data_0[3]; 
  assign entries_barrier_8_io_x_eff=superpage_entries_0_data_0[2]; 
  assign entries_barrier_8_io_x_c=superpage_entries_0_data_0[1]; 
  assign entries_barrier_9_io_x_ppn=superpage_entries_1_data_0[34:15]; 
  assign entries_barrier_9_io_x_u=superpage_entries_1_data_0[14]; 
  assign entries_barrier_9_io_x_ae=superpage_entries_1_data_0[12]; 
  assign entries_barrier_9_io_x_sw=superpage_entries_1_data_0[11]; 
  assign entries_barrier_9_io_x_sx=superpage_entries_1_data_0[10]; 
  assign entries_barrier_9_io_x_sr=superpage_entries_1_data_0[9]; 
  assign entries_barrier_9_io_x_pw=superpage_entries_1_data_0[8]; 
  assign entries_barrier_9_io_x_px=superpage_entries_1_data_0[7]; 
  assign entries_barrier_9_io_x_pr=superpage_entries_1_data_0[6]; 
  assign entries_barrier_9_io_x_ppp=superpage_entries_1_data_0[5]; 
  assign entries_barrier_9_io_x_pal=superpage_entries_1_data_0[4]; 
  assign entries_barrier_9_io_x_paa=superpage_entries_1_data_0[3]; 
  assign entries_barrier_9_io_x_eff=superpage_entries_1_data_0[2]; 
  assign entries_barrier_9_io_x_c=superpage_entries_1_data_0[1]; 
  assign entries_barrier_10_io_x_ppn=superpage_entries_2_data_0[34:15]; 
  assign entries_barrier_10_io_x_u=superpage_entries_2_data_0[14]; 
  assign entries_barrier_10_io_x_ae=superpage_entries_2_data_0[12]; 
  assign entries_barrier_10_io_x_sw=superpage_entries_2_data_0[11]; 
  assign entries_barrier_10_io_x_sx=superpage_entries_2_data_0[10]; 
  assign entries_barrier_10_io_x_sr=superpage_entries_2_data_0[9]; 
  assign entries_barrier_10_io_x_pw=superpage_entries_2_data_0[8]; 
  assign entries_barrier_10_io_x_px=superpage_entries_2_data_0[7]; 
  assign entries_barrier_10_io_x_pr=superpage_entries_2_data_0[6]; 
  assign entries_barrier_10_io_x_ppp=superpage_entries_2_data_0[5]; 
  assign entries_barrier_10_io_x_pal=superpage_entries_2_data_0[4]; 
  assign entries_barrier_10_io_x_paa=superpage_entries_2_data_0[3]; 
  assign entries_barrier_10_io_x_eff=superpage_entries_2_data_0[2]; 
  assign entries_barrier_10_io_x_c=superpage_entries_2_data_0[1]; 
  assign entries_barrier_11_io_x_ppn=superpage_entries_3_data_0[34:15]; 
  assign entries_barrier_11_io_x_u=superpage_entries_3_data_0[14]; 
  assign entries_barrier_11_io_x_ae=superpage_entries_3_data_0[12]; 
  assign entries_barrier_11_io_x_sw=superpage_entries_3_data_0[11]; 
  assign entries_barrier_11_io_x_sx=superpage_entries_3_data_0[10]; 
  assign entries_barrier_11_io_x_sr=superpage_entries_3_data_0[9]; 
  assign entries_barrier_11_io_x_pw=superpage_entries_3_data_0[8]; 
  assign entries_barrier_11_io_x_px=superpage_entries_3_data_0[7]; 
  assign entries_barrier_11_io_x_pr=superpage_entries_3_data_0[6]; 
  assign entries_barrier_11_io_x_ppp=superpage_entries_3_data_0[5]; 
  assign entries_barrier_11_io_x_pal=superpage_entries_3_data_0[4]; 
  assign entries_barrier_11_io_x_paa=superpage_entries_3_data_0[3]; 
  assign entries_barrier_11_io_x_eff=superpage_entries_3_data_0[2]; 
  assign entries_barrier_11_io_x_c=superpage_entries_3_data_0[1]; 
  assign entries_barrier_12_io_x_ppn=special_entry_data_0[34:15]; 
  assign entries_barrier_12_io_x_u=special_entry_data_0[14]; 
  assign entries_barrier_12_io_x_ae=special_entry_data_0[12]; 
  assign entries_barrier_12_io_x_sw=special_entry_data_0[11]; 
  assign entries_barrier_12_io_x_sx=special_entry_data_0[10]; 
  assign entries_barrier_12_io_x_sr=special_entry_data_0[9]; 
  assign entries_barrier_12_io_x_pw=special_entry_data_0[8]; 
  assign entries_barrier_12_io_x_px=special_entry_data_0[7]; 
  assign entries_barrier_12_io_x_pr=special_entry_data_0[6]; 
  assign entries_barrier_12_io_x_ppp=special_entry_data_0[5]; 
  assign entries_barrier_12_io_x_pal=special_entry_data_0[4]; 
  assign entries_barrier_12_io_x_paa=special_entry_data_0[3]; 
  assign entries_barrier_12_io_x_eff=special_entry_data_0[2]; 
  assign entries_barrier_12_io_x_c=special_entry_data_0[1]; 
  assign TLB_1_cov_read_addr=TLB_1_state; 
  assign TLB_1_cov_read_data=TLB_1_cov[TLB_1_cov_read_addr]; 
  assign TLB_1_cov_write_data=1'h1; 
  assign TLB_1_cov_write_addr=TLB_1_state; 
  assign TLB_1_cov_write_mask=1'h1; 
  assign TLB_1_cov_write_en=1'h1; 
  assign mux_cond_0=sectored_entries_0_6_data_1[0]; 
  assign mux_cond_1=sectored_entries_0_7_data_1[0]; 
  assign mux_cond_2=~sectored_entries_0_2_data_0[13]; 
  assign mux_cond_3=~sectored_entries_0_7_data_1[13]; 
  assign mux_cond_4=sectored_entries_0_7_data_3[0]; 
  assign mux_cond_5=sectored_entries_0_4_data_0[0]; 
  assign mux_cond_6=sectored_entries_0_3_data_3[0]; 
  assign mux_cond_7=sectored_entries_0_2_data_3[0]; 
  assign mux_cond_8=sectored_entries_0_2_data_0[0]; 
  assign mux_cond_9=~sectored_entries_0_6_data_1[13]; 
  assign mux_cond_10=~sectored_entries_0_2_data_2[13]; 
  assign mux_cond_11=~superpage_entries_0_data_0[13]; 
  assign mux_cond_12=sectored_entries_0_3_data_1[0]; 
  assign mux_cond_13=sectored_entries_0_4_data_3[0]; 
  assign mux_cond_14=~sectored_entries_0_3_data_3[13]; 
  assign mux_cond_15=sectored_entries_0_3_data_2[0]; 
  assign mux_cond_16=~sectored_entries_0_4_data_3[13]; 
  assign mux_cond_17=~sectored_entries_0_4_data_0[13]; 
  assign mux_cond_18=~sectored_entries_0_4_data_1[13]; 
  assign mux_cond_19=sectored_entries_0_6_data_0[0]; 
  assign mux_cond_20=sectored_entries_0_5_data_0[0]; 
  assign mux_cond_21=sectored_entries_0_6_data_2[0]; 
  assign mux_cond_22=sectored_entries_0_0_data_3[0]; 
  assign mux_cond_23=~sectored_entries_0_3_data_1[13]; 
  assign mux_cond_24=~sectored_entries_0_7_data_0[13]; 
  assign mux_cond_25=sectored_entries_0_7_data_0[0]; 
  assign mux_cond_26=~sectored_entries_0_7_data_3[13]; 
  assign mux_cond_27=~sectored_entries_0_0_data_3[13]; 
  assign mux_cond_28=~superpage_entries_1_data_0[13]; 
  assign mux_cond_29=~sectored_entries_0_7_data_2[13]; 
  assign mux_cond_30=~sectored_entries_0_6_data_0[13]; 
  assign mux_cond_31=~sectored_entries_0_6_data_3[13]; 
  assign mux_cond_32=sectored_entries_0_2_data_2[0]; 
  assign mux_cond_33=sectored_entries_0_1_data_1[0]; 
  assign mux_cond_34=~sectored_entries_0_2_data_1[13]; 
  assign mux_cond_35=~sectored_entries_0_4_data_2[13]; 
  assign mux_cond_36=~sectored_entries_0_1_data_3[13]; 
  assign mux_cond_37=~sectored_entries_0_0_data_2[13]; 
  assign mux_cond_38=~sectored_entries_0_0_data_0[13]; 
  assign mux_cond_39=~sectored_entries_0_2_data_3[13]; 
  assign mux_cond_40=sectored_entries_0_7_data_2[0]; 
  assign mux_cond_41=sectored_entries_0_0_data_0[0]; 
  assign mux_cond_42=~sectored_entries_0_5_data_0[13]; 
  assign mux_cond_43=sectored_entries_0_4_data_1[0]; 
  assign mux_cond_44=sectored_entries_0_5_data_1[0]; 
  assign mux_cond_45=~sectored_entries_0_5_data_3[13]; 
  assign mux_cond_46=sectored_entries_0_1_data_0[0]; 
  assign mux_cond_47=sectored_entries_0_5_data_3[0]; 
  assign mux_cond_48=~sectored_entries_0_0_data_1[13]; 
  assign mux_cond_49=~special_entry_data_0[13]; 
  assign mux_cond_50=~superpage_entries_2_data_0[13]; 
  assign mux_cond_51=sectored_entries_0_0_data_2[0]; 
  assign mux_cond_52=sectored_entries_0_6_data_3[0]; 
  assign mux_cond_53=~sectored_entries_0_3_data_0[13]; 
  assign mux_cond_54=~sectored_entries_0_1_data_0[13]; 
  assign mux_cond_55=sectored_entries_0_1_data_2[0]; 
  assign mux_cond_56=~sectored_entries_0_5_data_2[13]; 
  assign mux_cond_57=~sectored_entries_0_6_data_2[13]; 
  assign mux_cond_58=sectored_entries_0_1_data_3[0]; 
  assign mux_cond_59=~sectored_entries_0_3_data_2[13]; 
  assign mux_cond_60=~sectored_entries_0_1_data_1[13]; 
  assign mux_cond_61=~sectored_entries_0_1_data_2[13]; 
  assign mux_cond_62=sectored_entries_0_3_data_0[0]; 
  assign mux_cond_63=sectored_entries_0_5_data_2[0]; 
  assign mux_cond_64=sectored_entries_0_0_data_1[0]; 
  assign mux_cond_65=sectored_entries_0_2_data_1[0]; 
  assign mux_cond_66=~sectored_entries_0_5_data_1[13]; 
  assign mux_cond_67=~superpage_entries_3_data_0[13]; 
  assign mux_cond_68=sectored_entries_0_4_data_2[0]; 
  assign r_sectored_hit_shl=r_sectored_hit; 
  assign r_sectored_hit_pad={19'h0,r_sectored_hit_shl}; 
  assign r_sectored_repl_addr_shl={r_sectored_repl_addr,8'h0}; 
  assign r_sectored_repl_addr_pad={9'h0,r_sectored_repl_addr_shl}; 
  assign r_superpage_repl_addr_shl=r_superpage_repl_addr; 
  assign r_superpage_repl_addr_pad={18'h0,r_superpage_repl_addr_shl}; 
  assign special_entry_valid_0_shl={special_entry_valid_0,13'h0}; 
  assign special_entry_valid_0_pad={6'h0,special_entry_valid_0_shl}; 
  assign special_entry_level_shl={special_entry_level,12'h0}; 
  assign special_entry_level_pad={6'h0,special_entry_level_shl}; 
  assign state_shl={state,12'h0}; 
  assign state_pad={6'h0,state_shl}; 
  assign r_sectored_hit_addr_shl={r_sectored_hit_addr,1'h0}; 
  assign r_sectored_hit_addr_pad={16'h0,r_sectored_hit_addr_shl}; 
  assign mux_cond_0_shl={mux_cond_0,16'h0}; 
  assign mux_cond_0_pad={3'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,10'h0}; 
  assign mux_cond_1_pad={9'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl={mux_cond_2,2'h0}; 
  assign mux_cond_2_pad={17'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,15'h0}; 
  assign mux_cond_3_pad={4'h0,mux_cond_3_shl}; 
  assign mux_cond_4_shl={mux_cond_4,4'h0}; 
  assign mux_cond_4_pad={15'h0,mux_cond_4_shl}; 
  assign mux_cond_5_shl={mux_cond_5,13'h0}; 
  assign mux_cond_5_pad={6'h0,mux_cond_5_shl}; 
  assign mux_cond_6_shl={mux_cond_6,9'h0}; 
  assign mux_cond_6_pad={10'h0,mux_cond_6_shl}; 
  assign mux_cond_7_shl={mux_cond_7,8'h0}; 
  assign mux_cond_7_pad={11'h0,mux_cond_7_shl}; 
  assign mux_cond_8_shl={mux_cond_8,12'h0}; 
  assign mux_cond_8_pad={7'h0,mux_cond_8_shl}; 
  assign mux_cond_9_shl={mux_cond_9,19'h0}; 
  assign mux_cond_9_pad=mux_cond_9_shl; 
  assign mux_cond_10_shl={mux_cond_10,18'h0}; 
  assign mux_cond_10_pad={1'h0,mux_cond_10_shl}; 
  assign mux_cond_11_shl={mux_cond_11,9'h0}; 
  assign mux_cond_11_pad={10'h0,mux_cond_11_shl}; 
  assign mux_cond_12_shl={mux_cond_12,19'h0}; 
  assign mux_cond_12_pad=mux_cond_12_shl; 
  assign mux_cond_13_shl={mux_cond_13,7'h0}; 
  assign mux_cond_13_pad={12'h0,mux_cond_13_shl}; 
  assign mux_cond_14_shl={mux_cond_14,11'h0}; 
  assign mux_cond_14_pad={8'h0,mux_cond_14_shl}; 
  assign mux_cond_15_shl=mux_cond_15; 
  assign mux_cond_15_pad={19'h0,mux_cond_15_shl}; 
  assign mux_cond_16_shl={mux_cond_16,4'h0}; 
  assign mux_cond_16_pad={15'h0,mux_cond_16_shl}; 
  assign mux_cond_17_shl={mux_cond_17,19'h0}; 
  assign mux_cond_17_pad=mux_cond_17_shl; 
  assign mux_cond_18_shl={mux_cond_18,9'h0}; 
  assign mux_cond_18_pad={10'h0,mux_cond_18_shl}; 
  assign mux_cond_19_shl={mux_cond_19,8'h0}; 
  assign mux_cond_19_pad={11'h0,mux_cond_19_shl}; 
  assign mux_cond_20_shl={mux_cond_20,4'h0}; 
  assign mux_cond_20_pad={15'h0,mux_cond_20_shl}; 
  assign mux_cond_21_shl={mux_cond_21,6'h0}; 
  assign mux_cond_21_pad={13'h0,mux_cond_21_shl}; 
  assign mux_cond_22_shl={mux_cond_22,11'h0}; 
  assign mux_cond_22_pad={8'h0,mux_cond_22_shl}; 
  assign mux_cond_23_shl={mux_cond_23,14'h0}; 
  assign mux_cond_23_pad={5'h0,mux_cond_23_shl}; 
  assign mux_cond_24_shl={mux_cond_24,7'h0}; 
  assign mux_cond_24_pad={12'h0,mux_cond_24_shl}; 
  assign mux_cond_25_shl={mux_cond_25,7'h0}; 
  assign mux_cond_25_pad={12'h0,mux_cond_25_shl}; 
  assign mux_cond_26_shl={mux_cond_26,19'h0}; 
  assign mux_cond_26_pad=mux_cond_26_shl; 
  assign mux_cond_27_shl={mux_cond_27,10'h0}; 
  assign mux_cond_27_pad={9'h0,mux_cond_27_shl}; 
  assign mux_cond_28_shl={mux_cond_28,17'h0}; 
  assign mux_cond_28_pad={2'h0,mux_cond_28_shl}; 
  assign mux_cond_29_shl={mux_cond_29,3'h0}; 
  assign mux_cond_29_pad={16'h0,mux_cond_29_shl}; 
  assign mux_cond_30_shl={mux_cond_30,9'h0}; 
  assign mux_cond_30_pad={10'h0,mux_cond_30_shl}; 
  assign mux_cond_31_shl={mux_cond_31,15'h0}; 
  assign mux_cond_31_pad={4'h0,mux_cond_31_shl}; 
  assign mux_cond_32_shl=mux_cond_32; 
  assign mux_cond_32_pad={19'h0,mux_cond_32_shl}; 
  assign mux_cond_33_shl={mux_cond_33,12'h0}; 
  assign mux_cond_33_pad={7'h0,mux_cond_33_shl}; 
  assign mux_cond_34_shl={mux_cond_34,17'h0}; 
  assign mux_cond_34_pad={2'h0,mux_cond_34_shl}; 
  assign mux_cond_35_shl={mux_cond_35,9'h0}; 
  assign mux_cond_35_pad={10'h0,mux_cond_35_shl}; 
  assign mux_cond_36_shl={mux_cond_36,12'h0}; 
  assign mux_cond_36_pad={7'h0,mux_cond_36_shl}; 
  assign mux_cond_37_shl=mux_cond_37; 
  assign mux_cond_37_pad={19'h0,mux_cond_37_shl}; 
  assign mux_cond_38_shl={mux_cond_38,5'h0}; 
  assign mux_cond_38_pad={14'h0,mux_cond_38_shl}; 
  assign mux_cond_39_shl={mux_cond_39,2'h0}; 
  assign mux_cond_39_pad={17'h0,mux_cond_39_shl}; 
  assign mux_cond_40_shl={mux_cond_40,18'h0}; 
  assign mux_cond_40_pad={1'h0,mux_cond_40_shl}; 
  assign mux_cond_41_shl={mux_cond_41,13'h0}; 
  assign mux_cond_41_pad={6'h0,mux_cond_41_shl}; 
  assign mux_cond_42_shl={mux_cond_42,5'h0}; 
  assign mux_cond_42_pad={14'h0,mux_cond_42_shl}; 
  assign mux_cond_43_shl={mux_cond_43,18'h0}; 
  assign mux_cond_43_pad={1'h0,mux_cond_43_shl}; 
  assign mux_cond_44_shl={mux_cond_44,18'h0}; 
  assign mux_cond_44_pad={1'h0,mux_cond_44_shl}; 
  assign mux_cond_45_shl={mux_cond_45,2'h0}; 
  assign mux_cond_45_pad={17'h0,mux_cond_45_shl}; 
  assign mux_cond_46_shl={mux_cond_46,12'h0}; 
  assign mux_cond_46_pad={7'h0,mux_cond_46_shl}; 
  assign mux_cond_47_shl={mux_cond_47,18'h0}; 
  assign mux_cond_47_pad={1'h0,mux_cond_47_shl}; 
  assign mux_cond_48_shl={mux_cond_48,16'h0}; 
  assign mux_cond_48_pad={3'h0,mux_cond_48_shl}; 
  assign mux_cond_49_shl=mux_cond_49; 
  assign mux_cond_49_pad={19'h0,mux_cond_49_shl}; 
  assign mux_cond_50_shl={mux_cond_50,4'h0}; 
  assign mux_cond_50_pad={15'h0,mux_cond_50_shl}; 
  assign mux_cond_51_shl={mux_cond_51,9'h0}; 
  assign mux_cond_51_pad={10'h0,mux_cond_51_shl}; 
  assign mux_cond_52_shl={mux_cond_52,13'h0}; 
  assign mux_cond_52_pad={6'h0,mux_cond_52_shl}; 
  assign mux_cond_53_shl={mux_cond_53,4'h0}; 
  assign mux_cond_53_pad={15'h0,mux_cond_53_shl}; 
  assign mux_cond_54_shl={mux_cond_54,5'h0}; 
  assign mux_cond_54_pad={14'h0,mux_cond_54_shl}; 
  assign mux_cond_55_shl={mux_cond_55,10'h0}; 
  assign mux_cond_55_pad={9'h0,mux_cond_55_shl}; 
  assign mux_cond_56_shl={mux_cond_56,12'h0}; 
  assign mux_cond_56_pad={7'h0,mux_cond_56_shl}; 
  assign mux_cond_57_shl={mux_cond_57,4'h0}; 
  assign mux_cond_57_pad={15'h0,mux_cond_57_shl}; 
  assign mux_cond_58_shl={mux_cond_58,19'h0}; 
  assign mux_cond_58_pad=mux_cond_58_shl; 
  assign mux_cond_59_shl={mux_cond_59,8'h0}; 
  assign mux_cond_59_pad={11'h0,mux_cond_59_shl}; 
  assign mux_cond_60_shl={mux_cond_60,12'h0}; 
  assign mux_cond_60_pad={7'h0,mux_cond_60_shl}; 
  assign mux_cond_61_shl={mux_cond_61,13'h0}; 
  assign mux_cond_61_pad={6'h0,mux_cond_61_shl}; 
  assign mux_cond_62_shl={mux_cond_62,19'h0}; 
  assign mux_cond_62_pad=mux_cond_62_shl; 
  assign mux_cond_63_shl={mux_cond_63,7'h0}; 
  assign mux_cond_63_pad={12'h0,mux_cond_63_shl}; 
  assign mux_cond_64_shl={mux_cond_64,1'h0}; 
  assign mux_cond_64_pad={18'h0,mux_cond_64_shl}; 
  assign mux_cond_65_shl={mux_cond_65,3'h0}; 
  assign mux_cond_65_pad={16'h0,mux_cond_65_shl}; 
  assign mux_cond_66_shl={mux_cond_66,1'h0}; 
  assign mux_cond_66_pad={18'h0,mux_cond_66_shl}; 
  assign mux_cond_67_shl={mux_cond_67,15'h0}; 
  assign mux_cond_67_pad={4'h0,mux_cond_67_shl}; 
  assign mux_cond_68_shl={mux_cond_68,15'h0}; 
  assign mux_cond_68_pad={4'h0,mux_cond_68_shl}; 
  assign sectored_entries_0_0_valid_3_shl={sectored_entries_0_0_valid_3,5'h0}; 
  assign sectored_entries_0_0_valid_3_pad={14'h0,sectored_entries_0_0_valid_3_shl}; 
  assign sectored_entries_0_0_valid_2_shl={sectored_entries_0_0_valid_2,4'h0}; 
  assign sectored_entries_0_0_valid_2_pad={15'h0,sectored_entries_0_0_valid_2_shl}; 
  assign sectored_entries_0_2_valid_0_shl={sectored_entries_0_2_valid_0,5'h0}; 
  assign sectored_entries_0_2_valid_0_pad={14'h0,sectored_entries_0_2_valid_0_shl}; 
  assign sectored_entries_0_3_valid_0_shl={sectored_entries_0_3_valid_0,5'h0}; 
  assign sectored_entries_0_3_valid_0_pad={14'h0,sectored_entries_0_3_valid_0_shl}; 
  assign superpage_entries_2_level_shl={superpage_entries_2_level,13'h0}; 
  assign superpage_entries_2_level_pad={5'h0,superpage_entries_2_level_shl}; 
  assign sectored_entries_0_7_valid_1_shl={sectored_entries_0_7_valid_1,4'h0}; 
  assign sectored_entries_0_7_valid_1_pad={15'h0,sectored_entries_0_7_valid_1_shl}; 
  assign sectored_entries_0_4_valid_0_shl={sectored_entries_0_4_valid_0,5'h0}; 
  assign sectored_entries_0_4_valid_0_pad={14'h0,sectored_entries_0_4_valid_0_shl}; 
  assign sectored_entries_0_1_valid_3_shl={sectored_entries_0_1_valid_3,5'h0}; 
  assign sectored_entries_0_1_valid_3_pad={14'h0,sectored_entries_0_1_valid_3_shl}; 
  assign sectored_entries_0_1_valid_1_shl={sectored_entries_0_1_valid_1,4'h0}; 
  assign sectored_entries_0_1_valid_1_pad={15'h0,sectored_entries_0_1_valid_1_shl}; 
  assign sectored_entries_0_2_valid_3_shl={sectored_entries_0_2_valid_3,5'h0}; 
  assign sectored_entries_0_2_valid_3_pad={14'h0,sectored_entries_0_2_valid_3_shl}; 
  assign sectored_entries_0_2_valid_1_shl={sectored_entries_0_2_valid_1,4'h0}; 
  assign sectored_entries_0_2_valid_1_pad={15'h0,sectored_entries_0_2_valid_1_shl}; 
  assign superpage_entries_1_valid_0_shl={superpage_entries_1_valid_0,1'h0}; 
  assign superpage_entries_1_valid_0_pad={18'h0,superpage_entries_1_valid_0_shl}; 
  assign sectored_entries_0_7_valid_0_shl={sectored_entries_0_7_valid_0,5'h0}; 
  assign sectored_entries_0_7_valid_0_pad={14'h0,sectored_entries_0_7_valid_0_shl}; 
  assign superpage_entries_3_valid_0_shl={superpage_entries_3_valid_0,1'h0}; 
  assign superpage_entries_3_valid_0_pad={18'h0,superpage_entries_3_valid_0_shl}; 
  assign sectored_entries_0_5_valid_3_shl={sectored_entries_0_5_valid_3,5'h0}; 
  assign sectored_entries_0_5_valid_3_pad={14'h0,sectored_entries_0_5_valid_3_shl}; 
  assign sectored_entries_0_5_valid_1_shl={sectored_entries_0_5_valid_1,4'h0}; 
  assign sectored_entries_0_5_valid_1_pad={15'h0,sectored_entries_0_5_valid_1_shl}; 
  assign sectored_entries_0_4_valid_3_shl={sectored_entries_0_4_valid_3,5'h0}; 
  assign sectored_entries_0_4_valid_3_pad={14'h0,sectored_entries_0_4_valid_3_shl}; 
  assign sectored_entries_0_5_valid_2_shl={sectored_entries_0_5_valid_2,4'h0}; 
  assign sectored_entries_0_5_valid_2_pad={15'h0,sectored_entries_0_5_valid_2_shl}; 
  assign sectored_entries_0_1_valid_2_shl={sectored_entries_0_1_valid_2,4'h0}; 
  assign sectored_entries_0_1_valid_2_pad={15'h0,sectored_entries_0_1_valid_2_shl}; 
  assign sectored_entries_0_3_valid_1_shl={sectored_entries_0_3_valid_1,4'h0}; 
  assign sectored_entries_0_3_valid_1_pad={15'h0,sectored_entries_0_3_valid_1_shl}; 
  assign sectored_entries_0_1_valid_0_shl={sectored_entries_0_1_valid_0,5'h0}; 
  assign sectored_entries_0_1_valid_0_pad={14'h0,sectored_entries_0_1_valid_0_shl}; 
  assign sectored_entries_0_4_valid_2_shl={sectored_entries_0_4_valid_2,4'h0}; 
  assign sectored_entries_0_4_valid_2_pad={15'h0,sectored_entries_0_4_valid_2_shl}; 
  assign sectored_entries_0_4_valid_1_shl={sectored_entries_0_4_valid_1,4'h0}; 
  assign sectored_entries_0_4_valid_1_pad={15'h0,sectored_entries_0_4_valid_1_shl}; 
  assign superpage_entries_3_level_shl={superpage_entries_3_level,13'h0}; 
  assign superpage_entries_3_level_pad={5'h0,superpage_entries_3_level_shl}; 
  assign sectored_entries_0_0_valid_1_shl={sectored_entries_0_0_valid_1,4'h0}; 
  assign sectored_entries_0_0_valid_1_pad={15'h0,sectored_entries_0_0_valid_1_shl}; 
  assign sectored_entries_0_3_valid_2_shl={sectored_entries_0_3_valid_2,4'h0}; 
  assign sectored_entries_0_3_valid_2_pad={15'h0,sectored_entries_0_3_valid_2_shl}; 
  assign sectored_entries_0_6_valid_1_shl={sectored_entries_0_6_valid_1,4'h0}; 
  assign sectored_entries_0_6_valid_1_pad={15'h0,sectored_entries_0_6_valid_1_shl}; 
  assign sectored_entries_0_7_valid_3_shl={sectored_entries_0_7_valid_3,5'h0}; 
  assign sectored_entries_0_7_valid_3_pad={14'h0,sectored_entries_0_7_valid_3_shl}; 
  assign sectored_entries_0_3_valid_3_shl={sectored_entries_0_3_valid_3,5'h0}; 
  assign sectored_entries_0_3_valid_3_pad={14'h0,sectored_entries_0_3_valid_3_shl}; 
  assign sectored_entries_0_0_valid_0_shl={sectored_entries_0_0_valid_0,5'h0}; 
  assign sectored_entries_0_0_valid_0_pad={14'h0,sectored_entries_0_0_valid_0_shl}; 
  assign superpage_entries_0_valid_0_shl={superpage_entries_0_valid_0,1'h0}; 
  assign superpage_entries_0_valid_0_pad={18'h0,superpage_entries_0_valid_0_shl}; 
  assign sectored_entries_0_2_valid_2_shl={sectored_entries_0_2_valid_2,4'h0}; 
  assign sectored_entries_0_2_valid_2_pad={15'h0,sectored_entries_0_2_valid_2_shl}; 
  assign sectored_entries_0_6_valid_2_shl={sectored_entries_0_6_valid_2,4'h0}; 
  assign sectored_entries_0_6_valid_2_pad={15'h0,sectored_entries_0_6_valid_2_shl}; 
  assign superpage_entries_2_valid_0_shl={superpage_entries_2_valid_0,1'h0}; 
  assign superpage_entries_2_valid_0_pad={18'h0,superpage_entries_2_valid_0_shl}; 
  assign sectored_entries_0_6_valid_3_shl={sectored_entries_0_6_valid_3,5'h0}; 
  assign sectored_entries_0_6_valid_3_pad={14'h0,sectored_entries_0_6_valid_3_shl}; 
  assign sectored_entries_0_6_valid_0_shl={sectored_entries_0_6_valid_0,5'h0}; 
  assign sectored_entries_0_6_valid_0_pad={14'h0,sectored_entries_0_6_valid_0_shl}; 
  assign sectored_entries_0_7_valid_2_shl={sectored_entries_0_7_valid_2,4'h0}; 
  assign sectored_entries_0_7_valid_2_pad={15'h0,sectored_entries_0_7_valid_2_shl}; 
  assign superpage_entries_0_level_shl={superpage_entries_0_level,13'h0}; 
  assign superpage_entries_0_level_pad={5'h0,superpage_entries_0_level_shl}; 
  assign superpage_entries_1_level_shl={superpage_entries_1_level,13'h0}; 
  assign superpage_entries_1_level_pad={5'h0,superpage_entries_1_level_shl}; 
  assign sectored_entries_0_5_valid_0_shl={sectored_entries_0_5_valid_0,5'h0}; 
  assign sectored_entries_0_5_valid_0_pad={14'h0,sectored_entries_0_5_valid_0_shl}; 
  assign TLB_1_xor64=r_sectored_repl_addr_pad^r_superpage_repl_addr_pad; 
  assign TLB_1_xor31=r_sectored_hit_pad^TLB_1_xor64; 
  assign TLB_1_xor65=special_entry_valid_0_pad^special_entry_level_pad; 
  assign TLB_1_xor66=state_pad^r_sectored_hit_addr_pad; 
  assign TLB_1_xor32=TLB_1_xor65^TLB_1_xor66; 
  assign TLB_1_xor15=TLB_1_xor31^TLB_1_xor32; 
  assign TLB_1_xor68=mux_cond_1_pad^mux_cond_2_pad; 
  assign TLB_1_xor33=mux_cond_0_pad^TLB_1_xor68; 
  assign TLB_1_xor69=mux_cond_3_pad^mux_cond_4_pad; 
  assign TLB_1_xor70=mux_cond_5_pad^mux_cond_6_pad; 
  assign TLB_1_xor34=TLB_1_xor69^TLB_1_xor70; 
  assign TLB_1_xor16=TLB_1_xor33^TLB_1_xor34; 
  assign TLB_1_xor7=TLB_1_xor15^TLB_1_xor16; 
  assign TLB_1_xor72=mux_cond_8_pad^mux_cond_9_pad; 
  assign TLB_1_xor35=mux_cond_7_pad^TLB_1_xor72; 
  assign TLB_1_xor73=mux_cond_10_pad^mux_cond_11_pad; 
  assign TLB_1_xor74=mux_cond_12_pad^mux_cond_13_pad; 
  assign TLB_1_xor36=TLB_1_xor73^TLB_1_xor74; 
  assign TLB_1_xor17=TLB_1_xor35^TLB_1_xor36; 
  assign TLB_1_xor75=mux_cond_14_pad^mux_cond_15_pad; 
  assign TLB_1_xor76=mux_cond_16_pad^mux_cond_17_pad; 
  assign TLB_1_xor37=TLB_1_xor75^TLB_1_xor76; 
  assign TLB_1_xor77=mux_cond_18_pad^mux_cond_19_pad; 
  assign TLB_1_xor78=mux_cond_20_pad^mux_cond_21_pad; 
  assign TLB_1_xor38=TLB_1_xor77^TLB_1_xor78; 
  assign TLB_1_xor18=TLB_1_xor37^TLB_1_xor38; 
  assign TLB_1_xor8=TLB_1_xor17^TLB_1_xor18; 
  assign TLB_1_xor3=TLB_1_xor7^TLB_1_xor8; 
  assign TLB_1_xor80=mux_cond_23_pad^mux_cond_24_pad; 
  assign TLB_1_xor39=mux_cond_22_pad^TLB_1_xor80; 
  assign TLB_1_xor81=mux_cond_25_pad^mux_cond_26_pad; 
  assign TLB_1_xor82=mux_cond_27_pad^mux_cond_28_pad; 
  assign TLB_1_xor40=TLB_1_xor81^TLB_1_xor82; 
  assign TLB_1_xor19=TLB_1_xor39^TLB_1_xor40; 
  assign TLB_1_xor84=mux_cond_30_pad^mux_cond_31_pad; 
  assign TLB_1_xor41=mux_cond_29_pad^TLB_1_xor84; 
  assign TLB_1_xor85=mux_cond_32_pad^mux_cond_33_pad; 
  assign TLB_1_xor86=mux_cond_34_pad^mux_cond_35_pad; 
  assign TLB_1_xor42=TLB_1_xor85^TLB_1_xor86; 
  assign TLB_1_xor20=TLB_1_xor41^TLB_1_xor42; 
  assign TLB_1_xor9=TLB_1_xor19^TLB_1_xor20; 
  assign TLB_1_xor88=mux_cond_37_pad^mux_cond_38_pad; 
  assign TLB_1_xor43=mux_cond_36_pad^TLB_1_xor88; 
  assign TLB_1_xor89=mux_cond_39_pad^mux_cond_40_pad; 
  assign TLB_1_xor90=mux_cond_41_pad^mux_cond_42_pad; 
  assign TLB_1_xor44=TLB_1_xor89^TLB_1_xor90; 
  assign TLB_1_xor21=TLB_1_xor43^TLB_1_xor44; 
  assign TLB_1_xor91=mux_cond_43_pad^mux_cond_44_pad; 
  assign TLB_1_xor92=mux_cond_45_pad^mux_cond_46_pad; 
  assign TLB_1_xor45=TLB_1_xor91^TLB_1_xor92; 
  assign TLB_1_xor93=mux_cond_47_pad^mux_cond_48_pad; 
  assign TLB_1_xor94=mux_cond_49_pad^mux_cond_50_pad; 
  assign TLB_1_xor46=TLB_1_xor93^TLB_1_xor94; 
  assign TLB_1_xor22=TLB_1_xor45^TLB_1_xor46; 
  assign TLB_1_xor10=TLB_1_xor21^TLB_1_xor22; 
  assign TLB_1_xor4=TLB_1_xor9^TLB_1_xor10; 
  assign TLB_1_xor1=TLB_1_xor3^TLB_1_xor4; 
  assign TLB_1_xor96=mux_cond_52_pad^mux_cond_53_pad; 
  assign TLB_1_xor47=mux_cond_51_pad^TLB_1_xor96; 
  assign TLB_1_xor97=mux_cond_54_pad^mux_cond_55_pad; 
  assign TLB_1_xor98=mux_cond_56_pad^mux_cond_57_pad; 
  assign TLB_1_xor48=TLB_1_xor97^TLB_1_xor98; 
  assign TLB_1_xor23=TLB_1_xor47^TLB_1_xor48; 
  assign TLB_1_xor100=mux_cond_59_pad^mux_cond_60_pad; 
  assign TLB_1_xor49=mux_cond_58_pad^TLB_1_xor100; 
  assign TLB_1_xor101=mux_cond_61_pad^mux_cond_62_pad; 
  assign TLB_1_xor102=mux_cond_63_pad^mux_cond_64_pad; 
  assign TLB_1_xor50=TLB_1_xor101^TLB_1_xor102; 
  assign TLB_1_xor24=TLB_1_xor49^TLB_1_xor50; 
  assign TLB_1_xor11=TLB_1_xor23^TLB_1_xor24; 
  assign TLB_1_xor104=mux_cond_66_pad^mux_cond_67_pad; 
  assign TLB_1_xor51=mux_cond_65_pad^TLB_1_xor104; 
  assign TLB_1_xor105=mux_cond_68_pad^sectored_entries_0_0_valid_3_pad; 
  assign TLB_1_xor106=sectored_entries_0_0_valid_2_pad^sectored_entries_0_2_valid_0_pad; 
  assign TLB_1_xor52=TLB_1_xor105^TLB_1_xor106; 
  assign TLB_1_xor25=TLB_1_xor51^TLB_1_xor52; 
  assign TLB_1_xor107=sectored_entries_0_3_valid_0_pad^superpage_entries_2_level_pad; 
  assign TLB_1_xor108=sectored_entries_0_7_valid_1_pad^sectored_entries_0_4_valid_0_pad; 
  assign TLB_1_xor53=TLB_1_xor107^TLB_1_xor108; 
  assign TLB_1_xor109=sectored_entries_0_1_valid_3_pad^sectored_entries_0_1_valid_1_pad; 
  assign TLB_1_xor110=sectored_entries_0_2_valid_3_pad^sectored_entries_0_2_valid_1_pad; 
  assign TLB_1_xor54=TLB_1_xor109^TLB_1_xor110; 
  assign TLB_1_xor26=TLB_1_xor53^TLB_1_xor54; 
  assign TLB_1_xor12=TLB_1_xor25^TLB_1_xor26; 
  assign TLB_1_xor5=TLB_1_xor11^TLB_1_xor12; 
  assign TLB_1_xor112=sectored_entries_0_7_valid_0_pad^superpage_entries_3_valid_0_pad; 
  assign TLB_1_xor55=superpage_entries_1_valid_0_pad^TLB_1_xor112; 
  assign TLB_1_xor113=sectored_entries_0_5_valid_3_pad^sectored_entries_0_5_valid_1_pad; 
  assign TLB_1_xor114=sectored_entries_0_4_valid_3_pad^sectored_entries_0_5_valid_2_pad; 
  assign TLB_1_xor56=TLB_1_xor113^TLB_1_xor114; 
  assign TLB_1_xor27=TLB_1_xor55^TLB_1_xor56; 
  assign TLB_1_xor116=sectored_entries_0_3_valid_1_pad^sectored_entries_0_1_valid_0_pad; 
  assign TLB_1_xor57=sectored_entries_0_1_valid_2_pad^TLB_1_xor116; 
  assign TLB_1_xor117=sectored_entries_0_4_valid_2_pad^sectored_entries_0_4_valid_1_pad; 
  assign TLB_1_xor118=superpage_entries_3_level_pad^sectored_entries_0_0_valid_1_pad; 
  assign TLB_1_xor58=TLB_1_xor117^TLB_1_xor118; 
  assign TLB_1_xor28=TLB_1_xor57^TLB_1_xor58; 
  assign TLB_1_xor13=TLB_1_xor27^TLB_1_xor28; 
  assign TLB_1_xor120=sectored_entries_0_6_valid_1_pad^sectored_entries_0_7_valid_3_pad; 
  assign TLB_1_xor59=sectored_entries_0_3_valid_2_pad^TLB_1_xor120; 
  assign TLB_1_xor121=sectored_entries_0_3_valid_3_pad^sectored_entries_0_0_valid_0_pad; 
  assign TLB_1_xor122=superpage_entries_0_valid_0_pad^sectored_entries_0_2_valid_2_pad; 
  assign TLB_1_xor60=TLB_1_xor121^TLB_1_xor122; 
  assign TLB_1_xor29=TLB_1_xor59^TLB_1_xor60; 
  assign TLB_1_xor123=sectored_entries_0_6_valid_2_pad^superpage_entries_2_valid_0_pad; 
  assign TLB_1_xor124=sectored_entries_0_6_valid_3_pad^sectored_entries_0_6_valid_0_pad; 
  assign TLB_1_xor61=TLB_1_xor123^TLB_1_xor124; 
  assign TLB_1_xor125=sectored_entries_0_7_valid_2_pad^superpage_entries_0_level_pad; 
  assign TLB_1_xor126=superpage_entries_1_level_pad^sectored_entries_0_5_valid_0_pad; 
  assign TLB_1_xor62=TLB_1_xor125^TLB_1_xor126; 
  assign TLB_1_xor30=TLB_1_xor61^TLB_1_xor62; 
  assign TLB_1_xor14=TLB_1_xor29^TLB_1_xor30; 
  assign TLB_1_xor6=TLB_1_xor13^TLB_1_xor14; 
  assign TLB_1_xor2=TLB_1_xor5^TLB_1_xor6; 
  assign TLB_1_xor0=TLB_1_xor1^TLB_1_xor2; 
  assign mpu_ppn_barrier_sum=TLB_1_covSum+mpu_ppn_barrier_io_covSum; 
  assign entries_barrier_10_sum=mpu_ppn_barrier_sum+entries_barrier_10_io_covSum; 
  assign entries_barrier_9_sum=entries_barrier_10_sum+entries_barrier_9_io_covSum; 
  assign entries_barrier_7_sum=entries_barrier_9_sum+entries_barrier_7_io_covSum; 
  assign entries_barrier_sum=entries_barrier_7_sum+entries_barrier_io_covSum; 
  assign pmp_sum=entries_barrier_sum+pmp_io_covSum; 
  assign entries_barrier_6_sum=pmp_sum+entries_barrier_6_io_covSum; 
  assign entries_barrier_12_sum=entries_barrier_6_sum+entries_barrier_12_io_covSum; 
  assign entries_barrier_1_sum=entries_barrier_12_sum+entries_barrier_1_io_covSum; 
  assign entries_barrier_11_sum=entries_barrier_1_sum+entries_barrier_11_io_covSum; 
  assign entries_barrier_8_sum=entries_barrier_11_sum+entries_barrier_8_io_covSum; 
  assign entries_barrier_2_sum=entries_barrier_8_sum+entries_barrier_2_io_covSum; 
  assign entries_barrier_4_sum=entries_barrier_2_sum+entries_barrier_4_io_covSum; 
  assign entries_barrier_5_sum=entries_barrier_4_sum+entries_barrier_5_io_covSum; 
  assign entries_barrier_3_sum=entries_barrier_5_sum+entries_barrier_3_io_covSum; 
  assign io_covSum=entries_barrier_3_sum; 
  assign stopEn0=io_sfence_valid&~_T_51; 
  assign entries_barrier_12_metaAssert_wire=entries_barrier_12_metaAssert; 
  assign entries_barrier_metaAssert_wire=entries_barrier_metaAssert; 
  assign entries_barrier_10_metaAssert_wire=entries_barrier_10_metaAssert; 
  assign entries_barrier_5_metaAssert_wire=entries_barrier_5_metaAssert; 
  assign entries_barrier_11_metaAssert_wire=entries_barrier_11_metaAssert; 
  assign entries_barrier_9_metaAssert_wire=entries_barrier_9_metaAssert; 
  assign entries_barrier_8_metaAssert_wire=entries_barrier_8_metaAssert; 
  assign entries_barrier_1_metaAssert_wire=entries_barrier_1_metaAssert; 
  assign mpu_ppn_barrier_metaAssert_wire=mpu_ppn_barrier_metaAssert; 
  assign entries_barrier_4_metaAssert_wire=entries_barrier_4_metaAssert; 
  assign entries_barrier_6_metaAssert_wire=entries_barrier_6_metaAssert; 
  assign entries_barrier_3_metaAssert_wire=entries_barrier_3_metaAssert; 
  assign pmp_metaAssert_wire=pmp_metaAssert; 
  assign entries_barrier_7_metaAssert_wire=entries_barrier_7_metaAssert; 
  assign entries_barrier_2_metaAssert_wire=entries_barrier_2_metaAssert; 
  assign TLB_1_or7=stopEn0|entries_barrier_6_metaAssert_wire; 
  assign TLB_1_or8=entries_barrier_10_metaAssert_wire|entries_barrier_7_metaAssert_wire; 
  assign TLB_1_or3=TLB_1_or7|TLB_1_or8; 
  assign TLB_1_or9=entries_barrier_4_metaAssert_wire|entries_barrier_11_metaAssert_wire; 
  assign TLB_1_or10=entries_barrier_8_metaAssert_wire|entries_barrier_9_metaAssert_wire; 
  assign TLB_1_or4=TLB_1_or9|TLB_1_or10; 
  assign TLB_1_or1=TLB_1_or3|TLB_1_or4; 
  assign TLB_1_or11=entries_barrier_metaAssert_wire|entries_barrier_3_metaAssert_wire; 
  assign TLB_1_or12=pmp_metaAssert_wire|mpu_ppn_barrier_metaAssert_wire; 
  assign TLB_1_or5=TLB_1_or11|TLB_1_or12; 
  assign TLB_1_or13=entries_barrier_12_metaAssert_wire|entries_barrier_5_metaAssert_wire; 
  assign TLB_1_or14=entries_barrier_2_metaAssert_wire|entries_barrier_1_metaAssert_wire; 
  assign TLB_1_or6=TLB_1_or13|TLB_1_or14; 
  assign TLB_1_or2=TLB_1_or5|TLB_1_or6; 
  assign TLB_1_or0=TLB_1_or1|TLB_1_or2; 
  assign metaAssert=TLB_1_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              sectored_entries_0_0_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                sectored_entries_0_0_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_0_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_0_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_0_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_7)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_0_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_0[0])
                                 begin 
                                   sectored_entries_0_0_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_0 <=_GEN_53;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=_GEN_53;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_0 <=_GEN_53;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_0 <=_GEN_53;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_0 <=_GEN_621;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_0 <=_GEN_473;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_1[0])
                                 begin 
                                   sectored_entries_0_0_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_1 <=_GEN_54;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=_GEN_54;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_1 <=_GEN_54;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_1 <=_GEN_54;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_1 <=_GEN_622;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_1 <=_GEN_474;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_2[0])
                                 begin 
                                   sectored_entries_0_0_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_2 <=_GEN_55;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=_GEN_55;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_2 <=_GEN_55;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_2 <=_GEN_55;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_2 <=_GEN_623;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_2 <=_GEN_475;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_0_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_0_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_59)
                            begin 
                              if (sectored_entries_0_0_data_3[0])
                                 begin 
                                   sectored_entries_0_0_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_5)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_0_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_7)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_0_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_0_valid_3 <=_GEN_56;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=_GEN_56;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_5)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_0_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_7)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_0_valid_3 <=_GEN_56;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_7)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_0_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_0_valid_3 <=_GEN_56;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_0_valid_3 <=_GEN_624;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_0_valid_3 <=_GEN_476;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                sectored_entries_0_1_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_1_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_1_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_1_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_9)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_1_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_0[0])
                                 begin 
                                   sectored_entries_0_1_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_0 <=_GEN_79;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=_GEN_79;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_0 <=_GEN_79;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_0 <=_GEN_79;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_0 <=_GEN_649;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_0 <=_GEN_483;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_1[0])
                                 begin 
                                   sectored_entries_0_1_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_1 <=_GEN_80;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=_GEN_80;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_1 <=_GEN_80;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_1 <=_GEN_80;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_1 <=_GEN_650;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_1 <=_GEN_484;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_2[0])
                                 begin 
                                   sectored_entries_0_1_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_2 <=_GEN_81;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=_GEN_81;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_2 <=_GEN_81;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_2 <=_GEN_81;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_2 <=_GEN_651;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_2 <=_GEN_485;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_1_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_1_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_198)
                            begin 
                              if (sectored_entries_0_1_data_3[0])
                                 begin 
                                   sectored_entries_0_1_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_11)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_1_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_9)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_1_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_1_valid_3 <=_GEN_82;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=_GEN_82;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_11)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_1_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_9)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_1_valid_3 <=_GEN_82;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_9)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_1_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_1_valid_3 <=_GEN_82;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_1_valid_3 <=_GEN_652;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_1_valid_3 <=_GEN_486;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                sectored_entries_0_2_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_2_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_2_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_2_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_11)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_2_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_0[0])
                                 begin 
                                   sectored_entries_0_2_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_0 <=_GEN_105;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=_GEN_105;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_0 <=_GEN_105;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_0 <=_GEN_105;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_0 <=_GEN_677;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_0 <=_GEN_493;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_1[0])
                                 begin 
                                   sectored_entries_0_2_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_1 <=_GEN_106;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=_GEN_106;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_1 <=_GEN_106;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_1 <=_GEN_106;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_1 <=_GEN_678;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_1 <=_GEN_494;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_2[0])
                                 begin 
                                   sectored_entries_0_2_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_2 <=_GEN_107;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=_GEN_107;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_2 <=_GEN_107;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_2 <=_GEN_107;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_2 <=_GEN_679;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_2 <=_GEN_495;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_2_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_2_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_337)
                            begin 
                              if (sectored_entries_0_2_data_3[0])
                                 begin 
                                   sectored_entries_0_2_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_17)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_2_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_11)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_2_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_2_valid_3 <=_GEN_108;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=_GEN_108;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_17)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_2_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_11)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_2_valid_3 <=_GEN_108;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_11)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_2_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_2_valid_3 <=_GEN_108;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_2_valid_3 <=_GEN_680;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_2_valid_3 <=_GEN_496;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                sectored_entries_0_3_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_3_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_3_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_3_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_13)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_3_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_0[0])
                                 begin 
                                   sectored_entries_0_3_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_0 <=_GEN_131;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=_GEN_131;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_0 <=_GEN_131;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_0 <=_GEN_131;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_0 <=_GEN_705;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_0 <=_GEN_503;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_1[0])
                                 begin 
                                   sectored_entries_0_3_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_1 <=_GEN_132;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=_GEN_132;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_1 <=_GEN_132;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_1 <=_GEN_132;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_1 <=_GEN_706;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_1 <=_GEN_504;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_2[0])
                                 begin 
                                   sectored_entries_0_3_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_2 <=_GEN_133;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=_GEN_133;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_2 <=_GEN_133;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_2 <=_GEN_133;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_2 <=_GEN_707;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_2 <=_GEN_505;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_3_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_3_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_476)
                            begin 
                              if (sectored_entries_0_3_data_3[0])
                                 begin 
                                   sectored_entries_0_3_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_23)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_3_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_13)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_3_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_3_valid_3 <=_GEN_134;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=_GEN_134;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_23)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_3_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_13)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_3_valid_3 <=_GEN_134;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_13)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_3_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_3_valid_3 <=_GEN_134;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_3_valid_3 <=_GEN_708;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_3_valid_3 <=_GEN_506;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                sectored_entries_0_4_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_4_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_4_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_4_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_15)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_4_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_0[0])
                                 begin 
                                   sectored_entries_0_4_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_0 <=_GEN_157;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=_GEN_157;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_0 <=_GEN_157;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_0 <=_GEN_157;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_0 <=_GEN_733;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_0 <=_GEN_513;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_1[0])
                                 begin 
                                   sectored_entries_0_4_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_1 <=_GEN_158;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=_GEN_158;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_1 <=_GEN_158;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_1 <=_GEN_158;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_1 <=_GEN_734;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_1 <=_GEN_514;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_2[0])
                                 begin 
                                   sectored_entries_0_4_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_2 <=_GEN_159;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=_GEN_159;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_2 <=_GEN_159;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_2 <=_GEN_159;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_2 <=_GEN_735;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_2 <=_GEN_515;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_4_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_4_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_615)
                            begin 
                              if (sectored_entries_0_4_data_3[0])
                                 begin 
                                   sectored_entries_0_4_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_29)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_4_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_15)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_4_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_4_valid_3 <=_GEN_160;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=_GEN_160;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_29)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_4_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_15)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_4_valid_3 <=_GEN_160;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_15)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_4_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_4_valid_3 <=_GEN_160;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_4_valid_3 <=_GEN_736;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_4_valid_3 <=_GEN_516;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                sectored_entries_0_5_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_5_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_5_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_5_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_17)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_5_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_0[0])
                                 begin 
                                   sectored_entries_0_5_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_0 <=_GEN_183;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=_GEN_183;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_0 <=_GEN_183;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_0 <=_GEN_183;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_0 <=_GEN_761;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_0 <=_GEN_523;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_1[0])
                                 begin 
                                   sectored_entries_0_5_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_1 <=_GEN_184;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=_GEN_184;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_1 <=_GEN_184;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_1 <=_GEN_184;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_1 <=_GEN_762;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_1 <=_GEN_524;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_2[0])
                                 begin 
                                   sectored_entries_0_5_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_2 <=_GEN_185;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=_GEN_185;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_2 <=_GEN_185;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_2 <=_GEN_185;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_2 <=_GEN_763;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_2 <=_GEN_525;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_5_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_5_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_754)
                            begin 
                              if (sectored_entries_0_5_data_3[0])
                                 begin 
                                   sectored_entries_0_5_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_35)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_5_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_17)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_5_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_5_valid_3 <=_GEN_186;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=_GEN_186;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_35)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_5_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_17)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_5_valid_3 <=_GEN_186;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_17)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_5_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_5_valid_3 <=_GEN_186;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_5_valid_3 <=_GEN_764;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_5_valid_3 <=_GEN_526;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                sectored_entries_0_6_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_6_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_6_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_6_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_19)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_6_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_0[0])
                                 begin 
                                   sectored_entries_0_6_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_0 <=_GEN_209;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=_GEN_209;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_0 <=_GEN_209;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_0 <=_GEN_209;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_0 <=_GEN_789;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_0 <=_GEN_533;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_1[0])
                                 begin 
                                   sectored_entries_0_6_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_1 <=_GEN_210;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=_GEN_210;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_1 <=_GEN_210;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_1 <=_GEN_210;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_1 <=_GEN_790;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_1 <=_GEN_534;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_2[0])
                                 begin 
                                   sectored_entries_0_6_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_2 <=_GEN_211;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=_GEN_211;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_2 <=_GEN_211;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_2 <=_GEN_211;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_2 <=_GEN_791;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_2 <=_GEN_535;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_6_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_6_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_893)
                            begin 
                              if (sectored_entries_0_6_data_3[0])
                                 begin 
                                   sectored_entries_0_6_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_41)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_6_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_19)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_6_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_6_valid_3 <=_GEN_212;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=_GEN_212;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_41)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_6_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_19)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_6_valid_3 <=_GEN_212;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_19)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_6_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_6_valid_3 <=_GEN_212;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_6_valid_3 <=_GEN_792;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_6_valid_3 <=_GEN_536;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                sectored_entries_0_7_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h0==idx)
                                   begin 
                                     sectored_entries_0_7_data_0 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_1 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h1==idx)
                                   begin 
                                     sectored_entries_0_7_data_1 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_2 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h2==idx)
                                   begin 
                                     sectored_entries_0_7_data_2 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_data_3 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (!(_T_2))
                         begin 
                           if (_T_21)
                              begin 
                                if (2'h3==idx)
                                   begin 
                                     sectored_entries_0_7_data_3 <=_special_entry_data_0_T;
                                   end 
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_0[0])
                                 begin 
                                   sectored_entries_0_7_valid_0 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h0==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_0 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_0 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_0 <=_GEN_235;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=_GEN_235;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h0==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_0 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_0 <=_GEN_235;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_0 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_0 <=_GEN_235;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_0 <=_GEN_817;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_0 <=_GEN_543;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_1 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_1 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_1[0])
                                 begin 
                                   sectored_entries_0_7_valid_1 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h1==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_1 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_1 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_1 <=_GEN_236;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=_GEN_236;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h1==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_1 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_1 <=_GEN_236;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_1 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_1 <=_GEN_236;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_1 <=_GEN_818;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_1 <=_GEN_544;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_2 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_2 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_2[0])
                                 begin 
                                   sectored_entries_0_7_valid_2 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h2==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_2 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_2 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_2 <=_GEN_237;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=_GEN_237;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h2==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_2 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_2 <=_GEN_237;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_2 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_2 <=_GEN_237;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_2 <=_GEN_819;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_2 <=_GEN_545;
                  end 
         if (metaReset)
            begin 
              sectored_entries_0_7_valid_3 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 sectored_entries_0_7_valid_3 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_T_1032)
                            begin 
                              if (sectored_entries_0_7_data_3[0])
                                 begin 
                                   sectored_entries_0_7_valid_3 <=1'h0;
                                 end 
                               else 
                                 if (_sector_hits_T_47)
                                    begin 
                                      if (2'h3==hitsVec_idx)
                                         begin 
                                           sectored_entries_0_7_valid_3 <=1'h0;
                                         end 
                                       else 
                                         if (io_ptw_resp_valid)
                                            begin 
                                              if (!(~io_ptw_resp_bits_homogeneous))
                                                 begin 
                                                   if (!(_T_2))
                                                      begin 
                                                        if (_T_21)
                                                           begin 
                                                             if (invalidate_refill)
                                                                begin 
                                                                  sectored_entries_0_7_valid_3 <=1'h0;
                                                                end 
                                                              else 
                                                                begin 
                                                                  sectored_entries_0_7_valid_3 <=_GEN_238;
                                                                end 
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=_GEN_238;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                            end 
                          else 
                            if (_sector_hits_T_47)
                               begin 
                                 if (2'h3==hitsVec_idx)
                                    begin 
                                      sectored_entries_0_7_valid_3 <=1'h0;
                                    end 
                                  else 
                                    if (io_ptw_resp_valid)
                                       begin 
                                         if (!(~io_ptw_resp_bits_homogeneous))
                                            begin 
                                              if (!(_T_2))
                                                 begin 
                                                   if (_T_21)
                                                      begin 
                                                        if (invalidate_refill)
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=1'h0;
                                                           end 
                                                         else 
                                                           begin 
                                                             sectored_entries_0_7_valid_3 <=_GEN_238;
                                                           end 
                                                      end 
                                                 end 
                                            end 
                                       end 
                               end 
                             else 
                               if (io_ptw_resp_valid)
                                  begin 
                                    if (!(~io_ptw_resp_bits_homogeneous))
                                       begin 
                                         if (!(_T_2))
                                            begin 
                                              if (_T_21)
                                                 begin 
                                                   if (invalidate_refill)
                                                      begin 
                                                        sectored_entries_0_7_valid_3 <=1'h0;
                                                      end 
                                                    else 
                                                      begin 
                                                        sectored_entries_0_7_valid_3 <=_GEN_238;
                                                      end 
                                                 end 
                                            end 
                                       end 
                                  end 
                       end 
                     else 
                       begin 
                         sectored_entries_0_7_valid_3 <=_GEN_820;
                       end 
                  end 
                else 
                  begin 
                    sectored_entries_0_7_valid_3 <=_GEN_546;
                  end 
         if (metaReset)
            begin 
              superpage_entries_0_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_3)
                              begin 
                                superpage_entries_0_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_0_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_3)
                              begin 
                                superpage_entries_0_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_0_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_3)
                              begin 
                                superpage_entries_0_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_0_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_0_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_0)
                            begin 
                              superpage_entries_0_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_3)
                                              begin 
                                                if (invalidate_refill)
                                                   begin 
                                                     superpage_entries_0_valid_0 <=1'h0;
                                                   end 
                                                 else 
                                                   begin 
                                                     superpage_entries_0_valid_0 <=1'h1;
                                                   end 
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_0_valid_0 <=_GEN_827;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_3)
                                    begin 
                                      if (invalidate_refill)
                                         begin 
                                           superpage_entries_0_valid_0 <=1'h0;
                                         end 
                                       else 
                                         begin 
                                           superpage_entries_0_valid_0 <=1'h1;
                                         end 
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              superpage_entries_1_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_4)
                              begin 
                                superpage_entries_1_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_1_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_4)
                              begin 
                                superpage_entries_1_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_1_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_4)
                              begin 
                                superpage_entries_1_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_1_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_1_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_1)
                            begin 
                              superpage_entries_1_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_4)
                                              begin 
                                                if (invalidate_refill)
                                                   begin 
                                                     superpage_entries_1_valid_0 <=1'h0;
                                                   end 
                                                 else 
                                                   begin 
                                                     superpage_entries_1_valid_0 <=1'h1;
                                                   end 
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_1_valid_0 <=_GEN_831;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_4)
                                    begin 
                                      if (invalidate_refill)
                                         begin 
                                           superpage_entries_1_valid_0 <=1'h0;
                                         end 
                                       else 
                                         begin 
                                           superpage_entries_1_valid_0 <=1'h1;
                                         end 
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              superpage_entries_2_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_5)
                              begin 
                                superpage_entries_2_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_2_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_5)
                              begin 
                                superpage_entries_2_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_2_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_5)
                              begin 
                                superpage_entries_2_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_2_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_2_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_2)
                            begin 
                              superpage_entries_2_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_5)
                                              begin 
                                                superpage_entries_2_valid_0 <=_GEN_32;
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_2_valid_0 <=_GEN_835;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_5)
                                    begin 
                                      superpage_entries_2_valid_0 <=_GEN_32;
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              superpage_entries_3_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_6)
                              begin 
                                superpage_entries_3_level <={1'b0,io_ptw_resp_bits_level[0]};
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_3_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_6)
                              begin 
                                superpage_entries_3_tag <=r_refill_tag;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_3_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (!(~io_ptw_resp_bits_homogeneous))
                    begin 
                      if (_T_2)
                         begin 
                           if (_T_6)
                              begin 
                                superpage_entries_3_data_0 <=_special_entry_data_0_T;
                              end 
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              superpage_entries_3_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 superpage_entries_3_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (superpage_hits_3)
                            begin 
                              superpage_entries_3_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (!(~io_ptw_resp_bits_homogeneous))
                                    begin 
                                      if (_T_2)
                                         begin 
                                           if (_T_6)
                                              begin 
                                                superpage_entries_3_valid_0 <=_GEN_32;
                                              end 
                                         end 
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         superpage_entries_3_valid_0 <=_GEN_839;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (!(~io_ptw_resp_bits_homogeneous))
                          begin 
                            if (_T_2)
                               begin 
                                 if (_T_6)
                                    begin 
                                      superpage_entries_3_valid_0 <=_GEN_32;
                                    end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              special_entry_level <=2'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (~io_ptw_resp_bits_homogeneous)
                    begin 
                      special_entry_level <=io_ptw_resp_bits_level;
                    end 
               end 
         if (metaReset)
            begin 
              special_entry_tag <=27'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (~io_ptw_resp_bits_homogeneous)
                    begin 
                      special_entry_tag <=r_refill_tag;
                    end 
               end 
         if (metaReset)
            begin 
              special_entry_data_0 <=35'h0;
            end 
          else 
            if (io_ptw_resp_valid)
               begin 
                 if (~io_ptw_resp_bits_homogeneous)
                    begin 
                      special_entry_data_0 <=_special_entry_data_0_T;
                    end 
               end 
         if (metaReset)
            begin 
              special_entry_valid_0 <=1'h0;
            end 
          else 
            if (_T_1326)
               begin 
                 special_entry_valid_0 <=1'h0;
               end 
             else 
               if (io_sfence_valid)
                  begin 
                    if (io_sfence_bits_rs1)
                       begin 
                         if (_hitsVec_T_106)
                            begin 
                              special_entry_valid_0 <=1'h0;
                            end 
                          else 
                            if (io_ptw_resp_valid)
                               begin 
                                 if (~io_ptw_resp_bits_homogeneous)
                                    begin 
                                      special_entry_valid_0 <=_GEN_32;
                                    end 
                               end 
                       end 
                     else 
                       begin 
                         special_entry_valid_0 <=_GEN_843;
                       end 
                  end 
                else 
                  if (io_ptw_resp_valid)
                     begin 
                       if (~io_ptw_resp_bits_homogeneous)
                          begin 
                            special_entry_valid_0 <=_GEN_32;
                          end 
                     end 
         if (metaReset)
            begin 
              state <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 state <=2'h0;
               end 
             else 
               if (io_ptw_resp_valid)
                  begin 
                    state <=2'h0;
                  end 
                else 
                  if (_T_45)
                     begin 
                       state <=2'h3;
                     end 
                   else 
                     if (_invalidate_refill_T)
                        begin 
                          if (io_kill)
                             begin 
                               state <=2'h0;
                             end 
                           else 
                             if (io_ptw_req_ready)
                                begin 
                                  if (io_sfence_valid)
                                     begin 
                                       state <=2'h3;
                                     end 
                                   else 
                                     begin 
                                       state <=2'h2;
                                     end 
                                end 
                              else 
                                if (io_sfence_valid)
                                   begin 
                                     state <=2'h0;
                                   end 
                                 else 
                                   if (_T_42)
                                      begin 
                                        state <=2'h1;
                                      end 
                        end 
                      else 
                        if (_T_42)
                           begin 
                             state <=2'h1;
                           end 
         if (metaReset)
            begin 
              r_refill_tag <=27'h0;
            end 
          else 
            if (_T_42)
               begin 
                 r_refill_tag <=vpn;
               end 
         if (metaReset)
            begin 
              r_superpage_repl_addr <=2'h0;
            end 
          else 
            if (_T_42)
               begin 
                 if (_r_superpage_repl_addr_T_3)
                    begin 
                      r_superpage_repl_addr <=_r_superpage_repl_addr_T_2;
                    end 
                  else 
                    if (_r_superpage_repl_addr_T_5)
                       begin 
                         r_superpage_repl_addr <=2'h0;
                       end 
                     else 
                       if (_r_superpage_repl_addr_T_6)
                          begin 
                            r_superpage_repl_addr <=2'h1;
                          end 
                        else 
                          if (_r_superpage_repl_addr_T_7)
                             begin 
                               r_superpage_repl_addr <=2'h2;
                             end 
                           else 
                             begin 
                               r_superpage_repl_addr <=2'h3;
                             end 
               end 
         if (metaReset)
            begin 
              r_sectored_repl_addr <=3'h0;
            end 
          else 
            if (_T_42)
               begin 
                 if (_r_sectored_repl_addr_T_7)
                    begin 
                      r_sectored_repl_addr <=_r_sectored_repl_addr_T_6;
                    end 
                  else 
                    if (_r_sectored_repl_addr_T_9)
                       begin 
                         r_sectored_repl_addr <=3'h0;
                       end 
                     else 
                       if (_r_sectored_repl_addr_T_10)
                          begin 
                            r_sectored_repl_addr <=3'h1;
                          end 
                        else 
                          if (_r_sectored_repl_addr_T_11)
                             begin 
                               r_sectored_repl_addr <=3'h2;
                             end 
                           else 
                             if (_r_sectored_repl_addr_T_12)
                                begin 
                                  r_sectored_repl_addr <=3'h3;
                                end 
                              else 
                                if (_r_sectored_repl_addr_T_13)
                                   begin 
                                     r_sectored_repl_addr <=3'h4;
                                   end 
                                 else 
                                   if (_r_sectored_repl_addr_T_14)
                                      begin 
                                        r_sectored_repl_addr <=3'h5;
                                      end 
                                    else 
                                      if (_r_sectored_repl_addr_T_15)
                                         begin 
                                           r_sectored_repl_addr <=3'h6;
                                         end 
                                       else 
                                         begin 
                                           r_sectored_repl_addr <=3'h7;
                                         end 
               end 
         if (metaReset)
            begin 
              r_sectored_hit_addr <=3'h0;
            end 
          else 
            if (_T_42)
               begin 
                 r_sectored_hit_addr <=state_vec_0_touch_way_sized;
               end 
         if (metaReset)
            begin 
              r_sectored_hit <=1'h0;
            end 
          else 
            if (_T_42)
               begin 
                 r_sectored_hit <=_T_30;
               end 
         if (metaReset)
            begin 
              state_vec_0 <=7'h0;
            end 
          else 
            if (reset)
               begin 
                 state_vec_0 <=7'h0;
               end 
             else 
               if (_T_23)
                  begin 
                    if (_T_30)
                       begin 
                         state_vec_0 <=_state_vec_0_T_16;
                       end 
                  end 
         if (metaReset)
            begin 
              state_reg_1 <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 state_reg_1 <=3'h0;
               end 
             else 
               if (_T_23)
                  begin 
                    if (_T_37)
                       begin 
                         state_reg_1 <=_state_reg_T_6;
                       end 
                  end 
         if (io_sfence_valid&~_T_51)
            begin $display("Assertion failed\n    at TLB.scala:385 assert(!io.sfence.bits.rs1 || (io.sfence.bits.addr >> pgIdxBits) === vpn)\n");
            end 
         if (io_sfence_valid&~_T_51)
            begin $display("fatal");
            end 
         TLB_1_state <=TLB_1_xor0;
         if (!(TLB_1_cov_read_data))
            begin 
              TLB_1_covSum <=TLB_1_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              TLB_1_metaAssert <=1'h0;
            end 
          else 
            begin 
              TLB_1_metaAssert <=TLB_1_metaAssert|TLB_1_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (TLB_1_cov_write_en&TLB_1_cov_write_mask)
            begin 
              TLB_1_cov [TLB_1_cov_write_addr]<=TLB_1_cov_write_data;
            end 
       end
  
endmodule
 
module BTB (
  input clock,
  input reset,
  input [38:0] io_req_bits_addr,
  output io_resp_valid,
  output io_resp_bits_taken,
  output io_resp_bits_bridx,
  output [38:0] io_resp_bits_target,
  output [4:0] io_resp_bits_entry,
  output [7:0] io_resp_bits_bht_history,
  output io_resp_bits_bht_value,
  input io_btb_update_valid,
  input [4:0] io_btb_update_bits_prediction_entry,
  input [38:0] io_btb_update_bits_pc,
  input io_btb_update_bits_isValid,
  input [38:0] io_btb_update_bits_br_pc,
  input [1:0] io_btb_update_bits_cfiType,
  input io_bht_update_valid,
  input [7:0] io_bht_update_bits_prediction_history,
  input [38:0] io_bht_update_bits_pc,
  input io_bht_update_bits_branch,
  input io_bht_update_bits_taken,
  input io_bht_update_bits_mispredict,
  input io_bht_advance_valid,
  input io_bht_advance_bits_bht_value,
  input io_ras_update_valid,
  input [1:0] io_ras_update_bits_cfiType,
  input [38:0] io_ras_update_bits_returnAddr,
  output io_ras_head_valid,
  output [38:0] io_ras_head_bits,
  input io_flush,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg table_[0:511] ;  
   reg [31:0] _RAND_0 ;  
   wire table__res_res_value_MPORT_data ;  
   wire [8:0] table__res_res_value_MPORT_addr ;  
   wire table__MPORT_data ;  
   wire [8:0] table__MPORT_addr ;  
   wire table__MPORT_mask ;  
   wire table__MPORT_en ;  
   reg [12:0] idxs_0 ;  
   reg [31:0] _RAND_1 ;  
   reg [12:0] idxs_1 ;  
   reg [31:0] _RAND_2 ;  
   reg [12:0] idxs_2 ;  
   reg [31:0] _RAND_3 ;  
   reg [12:0] idxs_3 ;  
   reg [31:0] _RAND_4 ;  
   reg [12:0] idxs_4 ;  
   reg [31:0] _RAND_5 ;  
   reg [12:0] idxs_5 ;  
   reg [31:0] _RAND_6 ;  
   reg [12:0] idxs_6 ;  
   reg [31:0] _RAND_7 ;  
   reg [12:0] idxs_7 ;  
   reg [31:0] _RAND_8 ;  
   reg [12:0] idxs_8 ;  
   reg [31:0] _RAND_9 ;  
   reg [12:0] idxs_9 ;  
   reg [31:0] _RAND_10 ;  
   reg [12:0] idxs_10 ;  
   reg [31:0] _RAND_11 ;  
   reg [12:0] idxs_11 ;  
   reg [31:0] _RAND_12 ;  
   reg [12:0] idxs_12 ;  
   reg [31:0] _RAND_13 ;  
   reg [12:0] idxs_13 ;  
   reg [31:0] _RAND_14 ;  
   reg [12:0] idxs_14 ;  
   reg [31:0] _RAND_15 ;  
   reg [12:0] idxs_15 ;  
   reg [31:0] _RAND_16 ;  
   reg [12:0] idxs_16 ;  
   reg [31:0] _RAND_17 ;  
   reg [12:0] idxs_17 ;  
   reg [31:0] _RAND_18 ;  
   reg [12:0] idxs_18 ;  
   reg [31:0] _RAND_19 ;  
   reg [12:0] idxs_19 ;  
   reg [31:0] _RAND_20 ;  
   reg [12:0] idxs_20 ;  
   reg [31:0] _RAND_21 ;  
   reg [12:0] idxs_21 ;  
   reg [31:0] _RAND_22 ;  
   reg [12:0] idxs_22 ;  
   reg [31:0] _RAND_23 ;  
   reg [12:0] idxs_23 ;  
   reg [31:0] _RAND_24 ;  
   reg [12:0] idxs_24 ;  
   reg [31:0] _RAND_25 ;  
   reg [12:0] idxs_25 ;  
   reg [31:0] _RAND_26 ;  
   reg [12:0] idxs_26 ;  
   reg [31:0] _RAND_27 ;  
   reg [12:0] idxs_27 ;  
   reg [31:0] _RAND_28 ;  
   reg [2:0] idxPages_0 ;  
   reg [31:0] _RAND_29 ;  
   reg [2:0] idxPages_1 ;  
   reg [31:0] _RAND_30 ;  
   reg [2:0] idxPages_2 ;  
   reg [31:0] _RAND_31 ;  
   reg [2:0] idxPages_3 ;  
   reg [31:0] _RAND_32 ;  
   reg [2:0] idxPages_4 ;  
   reg [31:0] _RAND_33 ;  
   reg [2:0] idxPages_5 ;  
   reg [31:0] _RAND_34 ;  
   reg [2:0] idxPages_6 ;  
   reg [31:0] _RAND_35 ;  
   reg [2:0] idxPages_7 ;  
   reg [31:0] _RAND_36 ;  
   reg [2:0] idxPages_8 ;  
   reg [31:0] _RAND_37 ;  
   reg [2:0] idxPages_9 ;  
   reg [31:0] _RAND_38 ;  
   reg [2:0] idxPages_10 ;  
   reg [31:0] _RAND_39 ;  
   reg [2:0] idxPages_11 ;  
   reg [31:0] _RAND_40 ;  
   reg [2:0] idxPages_12 ;  
   reg [31:0] _RAND_41 ;  
   reg [2:0] idxPages_13 ;  
   reg [31:0] _RAND_42 ;  
   reg [2:0] idxPages_14 ;  
   reg [31:0] _RAND_43 ;  
   reg [2:0] idxPages_15 ;  
   reg [31:0] _RAND_44 ;  
   reg [2:0] idxPages_16 ;  
   reg [31:0] _RAND_45 ;  
   reg [2:0] idxPages_17 ;  
   reg [31:0] _RAND_46 ;  
   reg [2:0] idxPages_18 ;  
   reg [31:0] _RAND_47 ;  
   reg [2:0] idxPages_19 ;  
   reg [31:0] _RAND_48 ;  
   reg [2:0] idxPages_20 ;  
   reg [31:0] _RAND_49 ;  
   reg [2:0] idxPages_21 ;  
   reg [31:0] _RAND_50 ;  
   reg [2:0] idxPages_22 ;  
   reg [31:0] _RAND_51 ;  
   reg [2:0] idxPages_23 ;  
   reg [31:0] _RAND_52 ;  
   reg [2:0] idxPages_24 ;  
   reg [31:0] _RAND_53 ;  
   reg [2:0] idxPages_25 ;  
   reg [31:0] _RAND_54 ;  
   reg [2:0] idxPages_26 ;  
   reg [31:0] _RAND_55 ;  
   reg [2:0] idxPages_27 ;  
   reg [31:0] _RAND_56 ;  
   reg [12:0] tgts_0 ;  
   reg [31:0] _RAND_57 ;  
   reg [12:0] tgts_1 ;  
   reg [31:0] _RAND_58 ;  
   reg [12:0] tgts_2 ;  
   reg [31:0] _RAND_59 ;  
   reg [12:0] tgts_3 ;  
   reg [31:0] _RAND_60 ;  
   reg [12:0] tgts_4 ;  
   reg [31:0] _RAND_61 ;  
   reg [12:0] tgts_5 ;  
   reg [31:0] _RAND_62 ;  
   reg [12:0] tgts_6 ;  
   reg [31:0] _RAND_63 ;  
   reg [12:0] tgts_7 ;  
   reg [31:0] _RAND_64 ;  
   reg [12:0] tgts_8 ;  
   reg [31:0] _RAND_65 ;  
   reg [12:0] tgts_9 ;  
   reg [31:0] _RAND_66 ;  
   reg [12:0] tgts_10 ;  
   reg [31:0] _RAND_67 ;  
   reg [12:0] tgts_11 ;  
   reg [31:0] _RAND_68 ;  
   reg [12:0] tgts_12 ;  
   reg [31:0] _RAND_69 ;  
   reg [12:0] tgts_13 ;  
   reg [31:0] _RAND_70 ;  
   reg [12:0] tgts_14 ;  
   reg [31:0] _RAND_71 ;  
   reg [12:0] tgts_15 ;  
   reg [31:0] _RAND_72 ;  
   reg [12:0] tgts_16 ;  
   reg [31:0] _RAND_73 ;  
   reg [12:0] tgts_17 ;  
   reg [31:0] _RAND_74 ;  
   reg [12:0] tgts_18 ;  
   reg [31:0] _RAND_75 ;  
   reg [12:0] tgts_19 ;  
   reg [31:0] _RAND_76 ;  
   reg [12:0] tgts_20 ;  
   reg [31:0] _RAND_77 ;  
   reg [12:0] tgts_21 ;  
   reg [31:0] _RAND_78 ;  
   reg [12:0] tgts_22 ;  
   reg [31:0] _RAND_79 ;  
   reg [12:0] tgts_23 ;  
   reg [31:0] _RAND_80 ;  
   reg [12:0] tgts_24 ;  
   reg [31:0] _RAND_81 ;  
   reg [12:0] tgts_25 ;  
   reg [31:0] _RAND_82 ;  
   reg [12:0] tgts_26 ;  
   reg [31:0] _RAND_83 ;  
   reg [12:0] tgts_27 ;  
   reg [31:0] _RAND_84 ;  
   reg [2:0] tgtPages_0 ;  
   reg [31:0] _RAND_85 ;  
   reg [2:0] tgtPages_1 ;  
   reg [31:0] _RAND_86 ;  
   reg [2:0] tgtPages_2 ;  
   reg [31:0] _RAND_87 ;  
   reg [2:0] tgtPages_3 ;  
   reg [31:0] _RAND_88 ;  
   reg [2:0] tgtPages_4 ;  
   reg [31:0] _RAND_89 ;  
   reg [2:0] tgtPages_5 ;  
   reg [31:0] _RAND_90 ;  
   reg [2:0] tgtPages_6 ;  
   reg [31:0] _RAND_91 ;  
   reg [2:0] tgtPages_7 ;  
   reg [31:0] _RAND_92 ;  
   reg [2:0] tgtPages_8 ;  
   reg [31:0] _RAND_93 ;  
   reg [2:0] tgtPages_9 ;  
   reg [31:0] _RAND_94 ;  
   reg [2:0] tgtPages_10 ;  
   reg [31:0] _RAND_95 ;  
   reg [2:0] tgtPages_11 ;  
   reg [31:0] _RAND_96 ;  
   reg [2:0] tgtPages_12 ;  
   reg [31:0] _RAND_97 ;  
   reg [2:0] tgtPages_13 ;  
   reg [31:0] _RAND_98 ;  
   reg [2:0] tgtPages_14 ;  
   reg [31:0] _RAND_99 ;  
   reg [2:0] tgtPages_15 ;  
   reg [31:0] _RAND_100 ;  
   reg [2:0] tgtPages_16 ;  
   reg [31:0] _RAND_101 ;  
   reg [2:0] tgtPages_17 ;  
   reg [31:0] _RAND_102 ;  
   reg [2:0] tgtPages_18 ;  
   reg [31:0] _RAND_103 ;  
   reg [2:0] tgtPages_19 ;  
   reg [31:0] _RAND_104 ;  
   reg [2:0] tgtPages_20 ;  
   reg [31:0] _RAND_105 ;  
   reg [2:0] tgtPages_21 ;  
   reg [31:0] _RAND_106 ;  
   reg [2:0] tgtPages_22 ;  
   reg [31:0] _RAND_107 ;  
   reg [2:0] tgtPages_23 ;  
   reg [31:0] _RAND_108 ;  
   reg [2:0] tgtPages_24 ;  
   reg [31:0] _RAND_109 ;  
   reg [2:0] tgtPages_25 ;  
   reg [31:0] _RAND_110 ;  
   reg [2:0] tgtPages_26 ;  
   reg [31:0] _RAND_111 ;  
   reg [2:0] tgtPages_27 ;  
   reg [31:0] _RAND_112 ;  
   reg [24:0] pages_0 ;  
   reg [31:0] _RAND_113 ;  
   reg [24:0] pages_1 ;  
   reg [31:0] _RAND_114 ;  
   reg [24:0] pages_2 ;  
   reg [31:0] _RAND_115 ;  
   reg [24:0] pages_3 ;  
   reg [31:0] _RAND_116 ;  
   reg [24:0] pages_4 ;  
   reg [31:0] _RAND_117 ;  
   reg [24:0] pages_5 ;  
   reg [31:0] _RAND_118 ;  
   reg [5:0] pageValid ;  
   reg [31:0] _RAND_119 ;  
   wire [24:0] pagesMasked_0 ;  
   wire [24:0] pagesMasked_1 ;  
   wire [24:0] pagesMasked_2 ;  
   wire [24:0] pagesMasked_3 ;  
   wire [24:0] pagesMasked_4 ;  
   wire [24:0] pagesMasked_5 ;  
   reg [27:0] isValid ;  
   reg [31:0] _RAND_120 ;  
   reg [1:0] cfiType_0 ;  
   reg [31:0] _RAND_121 ;  
   reg [1:0] cfiType_1 ;  
   reg [31:0] _RAND_122 ;  
   reg [1:0] cfiType_2 ;  
   reg [31:0] _RAND_123 ;  
   reg [1:0] cfiType_3 ;  
   reg [31:0] _RAND_124 ;  
   reg [1:0] cfiType_4 ;  
   reg [31:0] _RAND_125 ;  
   reg [1:0] cfiType_5 ;  
   reg [31:0] _RAND_126 ;  
   reg [1:0] cfiType_6 ;  
   reg [31:0] _RAND_127 ;  
   reg [1:0] cfiType_7 ;  
   reg [31:0] _RAND_128 ;  
   reg [1:0] cfiType_8 ;  
   reg [31:0] _RAND_129 ;  
   reg [1:0] cfiType_9 ;  
   reg [31:0] _RAND_130 ;  
   reg [1:0] cfiType_10 ;  
   reg [31:0] _RAND_131 ;  
   reg [1:0] cfiType_11 ;  
   reg [31:0] _RAND_132 ;  
   reg [1:0] cfiType_12 ;  
   reg [31:0] _RAND_133 ;  
   reg [1:0] cfiType_13 ;  
   reg [31:0] _RAND_134 ;  
   reg [1:0] cfiType_14 ;  
   reg [31:0] _RAND_135 ;  
   reg [1:0] cfiType_15 ;  
   reg [31:0] _RAND_136 ;  
   reg [1:0] cfiType_16 ;  
   reg [31:0] _RAND_137 ;  
   reg [1:0] cfiType_17 ;  
   reg [31:0] _RAND_138 ;  
   reg [1:0] cfiType_18 ;  
   reg [31:0] _RAND_139 ;  
   reg [1:0] cfiType_19 ;  
   reg [31:0] _RAND_140 ;  
   reg [1:0] cfiType_20 ;  
   reg [31:0] _RAND_141 ;  
   reg [1:0] cfiType_21 ;  
   reg [31:0] _RAND_142 ;  
   reg [1:0] cfiType_22 ;  
   reg [31:0] _RAND_143 ;  
   reg [1:0] cfiType_23 ;  
   reg [31:0] _RAND_144 ;  
   reg [1:0] cfiType_24 ;  
   reg [31:0] _RAND_145 ;  
   reg [1:0] cfiType_25 ;  
   reg [31:0] _RAND_146 ;  
   reg [1:0] cfiType_26 ;  
   reg [31:0] _RAND_147 ;  
   reg [1:0] cfiType_27 ;  
   reg [31:0] _RAND_148 ;  
   reg brIdx_0 ;  
   reg [31:0] _RAND_149 ;  
   reg brIdx_1 ;  
   reg [31:0] _RAND_150 ;  
   reg brIdx_2 ;  
   reg [31:0] _RAND_151 ;  
   reg brIdx_3 ;  
   reg [31:0] _RAND_152 ;  
   reg brIdx_4 ;  
   reg [31:0] _RAND_153 ;  
   reg brIdx_5 ;  
   reg [31:0] _RAND_154 ;  
   reg brIdx_6 ;  
   reg [31:0] _RAND_155 ;  
   reg brIdx_7 ;  
   reg [31:0] _RAND_156 ;  
   reg brIdx_8 ;  
   reg [31:0] _RAND_157 ;  
   reg brIdx_9 ;  
   reg [31:0] _RAND_158 ;  
   reg brIdx_10 ;  
   reg [31:0] _RAND_159 ;  
   reg brIdx_11 ;  
   reg [31:0] _RAND_160 ;  
   reg brIdx_12 ;  
   reg [31:0] _RAND_161 ;  
   reg brIdx_13 ;  
   reg [31:0] _RAND_162 ;  
   reg brIdx_14 ;  
   reg [31:0] _RAND_163 ;  
   reg brIdx_15 ;  
   reg [31:0] _RAND_164 ;  
   reg brIdx_16 ;  
   reg [31:0] _RAND_165 ;  
   reg brIdx_17 ;  
   reg [31:0] _RAND_166 ;  
   reg brIdx_18 ;  
   reg [31:0] _RAND_167 ;  
   reg brIdx_19 ;  
   reg [31:0] _RAND_168 ;  
   reg brIdx_20 ;  
   reg [31:0] _RAND_169 ;  
   reg brIdx_21 ;  
   reg [31:0] _RAND_170 ;  
   reg brIdx_22 ;  
   reg [31:0] _RAND_171 ;  
   reg brIdx_23 ;  
   reg [31:0] _RAND_172 ;  
   reg brIdx_24 ;  
   reg [31:0] _RAND_173 ;  
   reg brIdx_25 ;  
   reg [31:0] _RAND_174 ;  
   reg brIdx_26 ;  
   reg [31:0] _RAND_175 ;  
   reg brIdx_27 ;  
   reg [31:0] _RAND_176 ;  
   reg r_btb_updatePipe_valid ;  
   reg [31:0] _RAND_177 ;  
   reg [4:0] r_btb_updatePipe_bits_prediction_entry ;  
   reg [31:0] _RAND_178 ;  
   reg [38:0] r_btb_updatePipe_bits_pc ;  
   reg [63:0] _RAND_179 ;  
   reg r_btb_updatePipe_bits_isValid ;  
   reg [31:0] _RAND_180 ;  
   reg [38:0] r_btb_updatePipe_bits_br_pc ;  
   reg [63:0] _RAND_181 ;  
   reg [1:0] r_btb_updatePipe_bits_cfiType ;  
   reg [31:0] _RAND_182 ;  
   wire [24:0] pageHit_p ;  
   wire pageHit_lo_lo ;  
   wire pageHit_lo_hi_lo ;  
   wire pageHit_lo_hi_hi ;  
   wire pageHit_hi_lo ;  
   wire pageHit_hi_hi_lo ;  
   wire pageHit_hi_hi_hi ;  
   wire [5:0] _pageHit_T ;  
   wire [5:0] pageHit ;  
   wire [12:0] idxHit_idx ;  
   wire idxHit_lo_lo_lo_lo ;  
   wire idxHit_lo_lo_lo_hi_lo ;  
   wire idxHit_lo_lo_lo_hi_hi ;  
   wire idxHit_lo_lo_hi_lo_lo ;  
   wire idxHit_lo_lo_hi_lo_hi ;  
   wire idxHit_lo_lo_hi_hi_lo ;  
   wire idxHit_lo_lo_hi_hi_hi ;  
   wire idxHit_lo_hi_lo_lo ;  
   wire idxHit_lo_hi_lo_hi_lo ;  
   wire idxHit_lo_hi_lo_hi_hi ;  
   wire idxHit_lo_hi_hi_lo_lo ;  
   wire idxHit_lo_hi_hi_lo_hi ;  
   wire idxHit_lo_hi_hi_hi_lo ;  
   wire idxHit_lo_hi_hi_hi_hi ;  
   wire idxHit_hi_lo_lo_lo ;  
   wire idxHit_hi_lo_lo_hi_lo ;  
   wire idxHit_hi_lo_lo_hi_hi ;  
   wire idxHit_hi_lo_hi_lo_lo ;  
   wire idxHit_hi_lo_hi_lo_hi ;  
   wire idxHit_hi_lo_hi_hi_lo ;  
   wire idxHit_hi_lo_hi_hi_hi ;  
   wire idxHit_hi_hi_lo_lo ;  
   wire idxHit_hi_hi_lo_hi_lo ;  
   wire idxHit_hi_hi_lo_hi_hi ;  
   wire idxHit_hi_hi_hi_lo_lo ;  
   wire idxHit_hi_hi_hi_lo_hi ;  
   wire idxHit_hi_hi_hi_hi_lo ;  
   wire idxHit_hi_hi_hi_hi_hi ;  
   wire [6:0] idxHit_lo_lo ;  
   wire [13:0] idxHit_lo ;  
   wire [6:0] idxHit_hi_lo ;  
   wire [27:0] _idxHit_T ;  
   wire [27:0] idxHit ;  
   wire [24:0] updatePageHit_p ;  
   wire updatePageHit_lo_lo ;  
   wire updatePageHit_lo_hi_lo ;  
   wire updatePageHit_lo_hi_hi ;  
   wire updatePageHit_hi_lo ;  
   wire updatePageHit_hi_hi_lo ;  
   wire updatePageHit_hi_hi_hi ;  
   wire [5:0] _updatePageHit_T ;  
   wire [5:0] updatePageHit ;  
   wire updateHit ;  
   wire useUpdatePageHit ;  
   wire usePageHit ;  
   wire doIdxPageRepl ;  
   reg [2:0] nextPageRepl ;  
   reg [31:0] _RAND_183 ;  
   wire [4:0] idxPageRepl_hi ;  
   wire idxPageRepl_lo ;  
   wire [5:0] _idxPageRepl_T ;  
   wire [7:0] _idxPageRepl_T_1 ;  
   wire [7:0] _idxPageRepl_T_2 ;  
   wire [7:0] _GEN_430 ;  
   wire [7:0] idxPageRepl ;  
   wire [7:0] idxPageUpdateOH ;  
   wire [3:0] idxPageUpdate_hi ;  
   wire [3:0] idxPageUpdate_lo ;  
   wire idxPageUpdate_hi_1 ;  
   wire [3:0] _idxPageUpdate_T ;  
   wire [1:0] idxPageUpdate_hi_2 ;  
   wire [1:0] idxPageUpdate_lo_1 ;  
   wire idxPageUpdate_hi_3 ;  
   wire [1:0] _idxPageUpdate_T_1 ;  
   wire idxPageUpdate_lo_2 ;  
   wire [2:0] idxPageUpdate ;  
   wire [7:0] idxPageReplEn ;  
   wire samePage ;  
   wire doTgtPageRepl ;  
   wire [4:0] tgtPageRepl_hi ;  
   wire tgtPageRepl_lo ;  
   wire [5:0] _tgtPageRepl_T ;  
   wire [7:0] tgtPageRepl ;  
   wire [7:0] _tgtPageUpdate_T ;  
   wire [7:0] _GEN_431 ;  
   wire [7:0] _tgtPageUpdate_T_1 ;  
   wire [3:0] tgtPageUpdate_hi ;  
   wire [3:0] tgtPageUpdate_lo ;  
   wire tgtPageUpdate_hi_1 ;  
   wire [3:0] _tgtPageUpdate_T_2 ;  
   wire [1:0] tgtPageUpdate_hi_2 ;  
   wire [1:0] tgtPageUpdate_lo_1 ;  
   wire tgtPageUpdate_hi_3 ;  
   wire [1:0] _tgtPageUpdate_T_3 ;  
   wire tgtPageUpdate_lo_2 ;  
   wire [2:0] tgtPageUpdate ;  
   wire [7:0] tgtPageReplEn ;  
   wire _T ;  
   wire _T_1 ;  
   wire both ;  
   wire [1:0] _next_T ;  
   wire [2:0] _GEN_432 ;  
   wire [2:0] next ;  
   wire _nextPageRepl_T ;  
   reg [26:0] state_reg ;  
   reg [31:0] _RAND_184 ;  
   wire waddr_hi ;  
   wire [10:0] waddr_left_subtree_state ;  
   wire [14:0] waddr_right_subtree_state ;  
   wire waddr_hi_1 ;  
   wire [2:0] waddr_left_subtree_state_1 ;  
   wire [6:0] waddr_right_subtree_state_1 ;  
   wire waddr_hi_2 ;  
   wire waddr_left_subtree_state_2 ;  
   wire waddr_right_subtree_state_2 ;  
   wire waddr_lo ;  
   wire [1:0] _waddr_T_2 ;  
   wire waddr_hi_3 ;  
   wire [2:0] waddr_left_subtree_state_3 ;  
   wire [2:0] waddr_right_subtree_state_3 ;  
   wire waddr_hi_4 ;  
   wire waddr_left_subtree_state_4 ;  
   wire waddr_right_subtree_state_4 ;  
   wire waddr_lo_1 ;  
   wire [1:0] _waddr_T_5 ;  
   wire waddr_hi_5 ;  
   wire waddr_left_subtree_state_5 ;  
   wire waddr_right_subtree_state_5 ;  
   wire waddr_lo_2 ;  
   wire [1:0] _waddr_T_8 ;  
   wire [1:0] waddr_lo_3 ;  
   wire [2:0] _waddr_T_9 ;  
   wire [2:0] waddr_lo_4 ;  
   wire [3:0] _waddr_T_10 ;  
   wire waddr_hi_6 ;  
   wire [6:0] waddr_left_subtree_state_6 ;  
   wire [6:0] waddr_right_subtree_state_6 ;  
   wire waddr_hi_7 ;  
   wire [2:0] waddr_left_subtree_state_7 ;  
   wire [2:0] waddr_right_subtree_state_7 ;  
   wire waddr_hi_8 ;  
   wire waddr_left_subtree_state_8 ;  
   wire waddr_right_subtree_state_8 ;  
   wire waddr_lo_5 ;  
   wire [1:0] _waddr_T_13 ;  
   wire waddr_hi_9 ;  
   wire waddr_left_subtree_state_9 ;  
   wire waddr_right_subtree_state_9 ;  
   wire waddr_lo_6 ;  
   wire [1:0] _waddr_T_16 ;  
   wire [1:0] waddr_lo_7 ;  
   wire [2:0] _waddr_T_17 ;  
   wire waddr_hi_10 ;  
   wire [2:0] waddr_left_subtree_state_10 ;  
   wire [2:0] waddr_right_subtree_state_10 ;  
   wire waddr_hi_11 ;  
   wire waddr_left_subtree_state_11 ;  
   wire waddr_right_subtree_state_11 ;  
   wire waddr_lo_8 ;  
   wire [1:0] _waddr_T_20 ;  
   wire waddr_hi_12 ;  
   wire waddr_left_subtree_state_12 ;  
   wire waddr_right_subtree_state_12 ;  
   wire waddr_lo_9 ;  
   wire [1:0] _waddr_T_23 ;  
   wire [1:0] waddr_lo_10 ;  
   wire [2:0] _waddr_T_24 ;  
   wire [2:0] waddr_lo_11 ;  
   wire [3:0] _waddr_T_25 ;  
   wire [3:0] waddr_lo_12 ;  
   wire [4:0] _waddr_T_26 ;  
   wire [4:0] waddr ;  
   reg r_respPipe_valid ;  
   reg [31:0] _RAND_185 ;  
   reg r_respPipe_bits_taken ;  
   reg [31:0] _RAND_186 ;  
   reg [4:0] r_respPipe_bits_entry ;  
   reg [31:0] _RAND_187 ;  
   wire _T_2 ;  
   wire _T_3 ;  
   wire [4:0] state_reg_touch_way_sized ;  
   wire state_reg_hi_hi ;  
   wire state_reg_hi_hi_1 ;  
   wire state_reg_hi_hi_2 ;  
   wire state_reg_hi_lo ;  
   wire state_reg_lo ;  
   wire [2:0] _state_reg_T_8 ;  
   wire [2:0] state_reg_hi_lo_1 ;  
   wire state_reg_hi_hi_3 ;  
   wire state_reg_hi_hi_4 ;  
   wire state_reg_hi_lo_2 ;  
   wire state_reg_lo_1 ;  
   wire [2:0] _state_reg_T_17 ;  
   wire [2:0] state_reg_hi_lo_3 ;  
   wire state_reg_hi_lo_4 ;  
   wire state_reg_lo_2 ;  
   wire [2:0] _state_reg_T_25 ;  
   wire [2:0] state_reg_lo_3 ;  
   wire [6:0] _state_reg_T_26 ;  
   wire [6:0] state_reg_lo_4 ;  
   wire [10:0] _state_reg_T_27 ;  
   wire [10:0] state_reg_hi_lo_5 ;  
   wire state_reg_hi_lo_6 ;  
   wire state_reg_lo_5 ;  
   wire [2:0] _state_reg_T_37 ;  
   wire [2:0] state_reg_hi_lo_7 ;  
   wire state_reg_hi_lo_8 ;  
   wire state_reg_lo_6 ;  
   wire [2:0] _state_reg_T_45 ;  
   wire [2:0] state_reg_lo_7 ;  
   wire [6:0] _state_reg_T_46 ;  
   wire [6:0] state_reg_hi_lo_9 ;  
   wire state_reg_hi_lo_10 ;  
   wire state_reg_lo_8 ;  
   wire [2:0] _state_reg_T_55 ;  
   wire [2:0] state_reg_hi_lo_11 ;  
   wire state_reg_hi_lo_12 ;  
   wire state_reg_lo_9 ;  
   wire [2:0] _state_reg_T_63 ;  
   wire [2:0] state_reg_lo_10 ;  
   wire [6:0] _state_reg_T_64 ;  
   wire [6:0] state_reg_lo_11 ;  
   wire [14:0] _state_reg_T_65 ;  
   wire [14:0] state_reg_lo_12 ;  
   wire [26:0] _state_reg_T_66 ;  
   wire [31:0] mask ;  
   wire [3:0] _idxPages_T ;  
   wire [31:0] _GEN_433 ;  
   wire [31:0] _isValid_T ;  
   wire [31:0] _isValid_T_2 ;  
   wire [31:0] _isValid_T_3 ;  
   wire idxWritesEven ;  
   wire [7:0] _T_5 ;  
   wire [7:0] _T_12 ;  
   wire [7:0] _GEN_435 ;  
   wire [7:0] _pageValid_T ;  
   wire [7:0] _pageValid_T_1 ;  
   wire [31:0] _GEN_338 ;  
   wire [7:0] _GEN_373 ;  
   wire [6:0] _io_resp_valid_T ;  
   wire [2:0] _io_resp_valid_T_29 ;  
   wire [2:0] _io_resp_valid_T_30 ;  
   wire [2:0] _io_resp_valid_T_31 ;  
   wire [2:0] _io_resp_valid_T_32 ;  
   wire [2:0] _io_resp_valid_T_33 ;  
   wire [2:0] _io_resp_valid_T_34 ;  
   wire [2:0] _io_resp_valid_T_35 ;  
   wire [2:0] _io_resp_valid_T_36 ;  
   wire [2:0] _io_resp_valid_T_37 ;  
   wire [2:0] _io_resp_valid_T_38 ;  
   wire [2:0] _io_resp_valid_T_39 ;  
   wire [2:0] _io_resp_valid_T_40 ;  
   wire [2:0] _io_resp_valid_T_41 ;  
   wire [2:0] _io_resp_valid_T_42 ;  
   wire [2:0] _io_resp_valid_T_43 ;  
   wire [2:0] _io_resp_valid_T_44 ;  
   wire [2:0] _io_resp_valid_T_45 ;  
   wire [2:0] _io_resp_valid_T_46 ;  
   wire [2:0] _io_resp_valid_T_47 ;  
   wire [2:0] _io_resp_valid_T_48 ;  
   wire [2:0] _io_resp_valid_T_49 ;  
   wire [2:0] _io_resp_valid_T_50 ;  
   wire [2:0] _io_resp_valid_T_51 ;  
   wire [2:0] _io_resp_valid_T_52 ;  
   wire [2:0] _io_resp_valid_T_53 ;  
   wire [2:0] _io_resp_valid_T_54 ;  
   wire [2:0] _io_resp_valid_T_55 ;  
   wire [2:0] _io_resp_valid_T_56 ;  
   wire [2:0] _io_resp_valid_T_57 ;  
   wire [2:0] _io_resp_valid_T_58 ;  
   wire [2:0] _io_resp_valid_T_59 ;  
   wire [2:0] _io_resp_valid_T_60 ;  
   wire [2:0] _io_resp_valid_T_61 ;  
   wire [2:0] _io_resp_valid_T_62 ;  
   wire [2:0] _io_resp_valid_T_63 ;  
   wire [2:0] _io_resp_valid_T_64 ;  
   wire [2:0] _io_resp_valid_T_65 ;  
   wire [2:0] _io_resp_valid_T_66 ;  
   wire [2:0] _io_resp_valid_T_67 ;  
   wire [2:0] _io_resp_valid_T_68 ;  
   wire [2:0] _io_resp_valid_T_69 ;  
   wire [2:0] _io_resp_valid_T_70 ;  
   wire [2:0] _io_resp_valid_T_71 ;  
   wire [2:0] _io_resp_valid_T_72 ;  
   wire [2:0] _io_resp_valid_T_73 ;  
   wire [2:0] _io_resp_valid_T_74 ;  
   wire [2:0] _io_resp_valid_T_75 ;  
   wire [2:0] _io_resp_valid_T_76 ;  
   wire [2:0] _io_resp_valid_T_77 ;  
   wire [2:0] _io_resp_valid_T_78 ;  
   wire [2:0] _io_resp_valid_T_79 ;  
   wire [2:0] _io_resp_valid_T_80 ;  
   wire [2:0] _io_resp_valid_T_81 ;  
   wire [2:0] _io_resp_valid_T_82 ;  
   wire [2:0] _io_resp_valid_T_83 ;  
   wire [6:0] _io_resp_valid_T_84 ;  
   wire [2:0] _io_resp_bits_target_T_28 ;  
   wire [2:0] _io_resp_bits_target_T_29 ;  
   wire [2:0] _io_resp_bits_target_T_30 ;  
   wire [2:0] _io_resp_bits_target_T_31 ;  
   wire [2:0] _io_resp_bits_target_T_32 ;  
   wire [2:0] _io_resp_bits_target_T_33 ;  
   wire [2:0] _io_resp_bits_target_T_34 ;  
   wire [2:0] _io_resp_bits_target_T_35 ;  
   wire [2:0] _io_resp_bits_target_T_36 ;  
   wire [2:0] _io_resp_bits_target_T_37 ;  
   wire [2:0] _io_resp_bits_target_T_38 ;  
   wire [2:0] _io_resp_bits_target_T_39 ;  
   wire [2:0] _io_resp_bits_target_T_40 ;  
   wire [2:0] _io_resp_bits_target_T_41 ;  
   wire [2:0] _io_resp_bits_target_T_42 ;  
   wire [2:0] _io_resp_bits_target_T_43 ;  
   wire [2:0] _io_resp_bits_target_T_44 ;  
   wire [2:0] _io_resp_bits_target_T_45 ;  
   wire [2:0] _io_resp_bits_target_T_46 ;  
   wire [2:0] _io_resp_bits_target_T_47 ;  
   wire [2:0] _io_resp_bits_target_T_48 ;  
   wire [2:0] _io_resp_bits_target_T_49 ;  
   wire [2:0] _io_resp_bits_target_T_50 ;  
   wire [2:0] _io_resp_bits_target_T_51 ;  
   wire [2:0] _io_resp_bits_target_T_52 ;  
   wire [2:0] _io_resp_bits_target_T_53 ;  
   wire [2:0] _io_resp_bits_target_T_54 ;  
   wire [2:0] _io_resp_bits_target_T_55 ;  
   wire [2:0] _io_resp_bits_target_T_56 ;  
   wire [2:0] _io_resp_bits_target_T_57 ;  
   wire [2:0] _io_resp_bits_target_T_58 ;  
   wire [2:0] _io_resp_bits_target_T_59 ;  
   wire [2:0] _io_resp_bits_target_T_60 ;  
   wire [2:0] _io_resp_bits_target_T_61 ;  
   wire [2:0] _io_resp_bits_target_T_62 ;  
   wire [2:0] _io_resp_bits_target_T_63 ;  
   wire [2:0] _io_resp_bits_target_T_64 ;  
   wire [2:0] _io_resp_bits_target_T_65 ;  
   wire [2:0] _io_resp_bits_target_T_66 ;  
   wire [2:0] _io_resp_bits_target_T_67 ;  
   wire [2:0] _io_resp_bits_target_T_68 ;  
   wire [2:0] _io_resp_bits_target_T_69 ;  
   wire [2:0] _io_resp_bits_target_T_70 ;  
   wire [2:0] _io_resp_bits_target_T_71 ;  
   wire [2:0] _io_resp_bits_target_T_72 ;  
   wire [2:0] _io_resp_bits_target_T_73 ;  
   wire [2:0] _io_resp_bits_target_T_74 ;  
   wire [2:0] _io_resp_bits_target_T_75 ;  
   wire [2:0] _io_resp_bits_target_T_76 ;  
   wire [2:0] _io_resp_bits_target_T_77 ;  
   wire [2:0] _io_resp_bits_target_T_78 ;  
   wire [2:0] _io_resp_bits_target_T_79 ;  
   wire [2:0] _io_resp_bits_target_T_80 ;  
   wire [2:0] _io_resp_bits_target_T_81 ;  
   wire [2:0] _io_resp_bits_target_T_82 ;  
   wire _io_resp_bits_target_T_83 ;  
   wire [24:0] _io_resp_bits_target_T_84 ;  
   wire _io_resp_bits_target_T_85 ;  
   wire [24:0] _io_resp_bits_target_T_86 ;  
   wire _io_resp_bits_target_T_87 ;  
   wire [24:0] _io_resp_bits_target_T_88 ;  
   wire _io_resp_bits_target_T_89 ;  
   wire [24:0] _io_resp_bits_target_T_90 ;  
   wire _io_resp_bits_target_T_91 ;  
   wire [24:0] _io_resp_bits_target_T_92 ;  
   wire _io_resp_bits_target_T_93 ;  
   wire [24:0] _io_resp_bits_target_T_94 ;  
   wire _io_resp_bits_target_T_95 ;  
   wire [24:0] io_resp_bits_target_hi ;  
   wire [12:0] _io_resp_bits_target_T_124 ;  
   wire [12:0] _io_resp_bits_target_T_125 ;  
   wire [12:0] _io_resp_bits_target_T_126 ;  
   wire [12:0] _io_resp_bits_target_T_127 ;  
   wire [12:0] _io_resp_bits_target_T_128 ;  
   wire [12:0] _io_resp_bits_target_T_129 ;  
   wire [12:0] _io_resp_bits_target_T_130 ;  
   wire [12:0] _io_resp_bits_target_T_131 ;  
   wire [12:0] _io_resp_bits_target_T_132 ;  
   wire [12:0] _io_resp_bits_target_T_133 ;  
   wire [12:0] _io_resp_bits_target_T_134 ;  
   wire [12:0] _io_resp_bits_target_T_135 ;  
   wire [12:0] _io_resp_bits_target_T_136 ;  
   wire [12:0] _io_resp_bits_target_T_137 ;  
   wire [12:0] _io_resp_bits_target_T_138 ;  
   wire [12:0] _io_resp_bits_target_T_139 ;  
   wire [12:0] _io_resp_bits_target_T_140 ;  
   wire [12:0] _io_resp_bits_target_T_141 ;  
   wire [12:0] _io_resp_bits_target_T_142 ;  
   wire [12:0] _io_resp_bits_target_T_143 ;  
   wire [12:0] _io_resp_bits_target_T_144 ;  
   wire [12:0] _io_resp_bits_target_T_145 ;  
   wire [12:0] _io_resp_bits_target_T_146 ;  
   wire [12:0] _io_resp_bits_target_T_147 ;  
   wire [12:0] _io_resp_bits_target_T_148 ;  
   wire [12:0] _io_resp_bits_target_T_149 ;  
   wire [12:0] _io_resp_bits_target_T_150 ;  
   wire [12:0] _io_resp_bits_target_T_151 ;  
   wire [12:0] _io_resp_bits_target_T_152 ;  
   wire [12:0] _io_resp_bits_target_T_153 ;  
   wire [12:0] _io_resp_bits_target_T_154 ;  
   wire [12:0] _io_resp_bits_target_T_155 ;  
   wire [12:0] _io_resp_bits_target_T_156 ;  
   wire [12:0] _io_resp_bits_target_T_157 ;  
   wire [12:0] _io_resp_bits_target_T_158 ;  
   wire [12:0] _io_resp_bits_target_T_159 ;  
   wire [12:0] _io_resp_bits_target_T_160 ;  
   wire [12:0] _io_resp_bits_target_T_161 ;  
   wire [12:0] _io_resp_bits_target_T_162 ;  
   wire [12:0] _io_resp_bits_target_T_163 ;  
   wire [12:0] _io_resp_bits_target_T_164 ;  
   wire [12:0] _io_resp_bits_target_T_165 ;  
   wire [12:0] _io_resp_bits_target_T_166 ;  
   wire [12:0] _io_resp_bits_target_T_167 ;  
   wire [12:0] _io_resp_bits_target_T_168 ;  
   wire [12:0] _io_resp_bits_target_T_169 ;  
   wire [12:0] _io_resp_bits_target_T_170 ;  
   wire [12:0] _io_resp_bits_target_T_171 ;  
   wire [12:0] _io_resp_bits_target_T_172 ;  
   wire [12:0] _io_resp_bits_target_T_173 ;  
   wire [12:0] _io_resp_bits_target_T_174 ;  
   wire [12:0] _io_resp_bits_target_T_175 ;  
   wire [12:0] _io_resp_bits_target_T_176 ;  
   wire [12:0] _io_resp_bits_target_T_177 ;  
   wire [12:0] _io_resp_bits_target_T_178 ;  
   wire [13:0] io_resp_bits_target_lo ;  
   wire [38:0] _io_resp_bits_target_T_179 ;  
   wire [11:0] io_resp_bits_entry_hi ;  
   wire [15:0] io_resp_bits_entry_lo ;  
   wire io_resp_bits_entry_hi_1 ;  
   wire [15:0] _GEN_436 ;  
   wire [15:0] _io_resp_bits_entry_T ;  
   wire [7:0] io_resp_bits_entry_hi_2 ;  
   wire [7:0] io_resp_bits_entry_lo_1 ;  
   wire io_resp_bits_entry_hi_3 ;  
   wire [7:0] _io_resp_bits_entry_T_1 ;  
   wire [3:0] io_resp_bits_entry_hi_4 ;  
   wire [3:0] io_resp_bits_entry_lo_2 ;  
   wire io_resp_bits_entry_hi_5 ;  
   wire [3:0] _io_resp_bits_entry_T_2 ;  
   wire [1:0] io_resp_bits_entry_hi_6 ;  
   wire [1:0] io_resp_bits_entry_lo_3 ;  
   wire io_resp_bits_entry_hi_7 ;  
   wire [1:0] _io_resp_bits_entry_T_3 ;  
   wire io_resp_bits_entry_lo_4 ;  
   wire [3:0] io_resp_bits_entry_lo_7 ;  
   wire _io_resp_bits_bridx_T_28 ;  
   wire _io_resp_bits_bridx_T_29 ;  
   wire _io_resp_bits_bridx_T_30 ;  
   wire _io_resp_bits_bridx_T_31 ;  
   wire _io_resp_bits_bridx_T_32 ;  
   wire _io_resp_bits_bridx_T_33 ;  
   wire _io_resp_bits_bridx_T_34 ;  
   wire _io_resp_bits_bridx_T_35 ;  
   wire _io_resp_bits_bridx_T_36 ;  
   wire _io_resp_bits_bridx_T_37 ;  
   wire _io_resp_bits_bridx_T_38 ;  
   wire _io_resp_bits_bridx_T_39 ;  
   wire _io_resp_bits_bridx_T_40 ;  
   wire _io_resp_bits_bridx_T_41 ;  
   wire _io_resp_bits_bridx_T_42 ;  
   wire _io_resp_bits_bridx_T_43 ;  
   wire _io_resp_bits_bridx_T_44 ;  
   wire _io_resp_bits_bridx_T_45 ;  
   wire _io_resp_bits_bridx_T_46 ;  
   wire _io_resp_bits_bridx_T_47 ;  
   wire _io_resp_bits_bridx_T_48 ;  
   wire _io_resp_bits_bridx_T_49 ;  
   wire _io_resp_bits_bridx_T_50 ;  
   wire _io_resp_bits_bridx_T_51 ;  
   wire _io_resp_bits_bridx_T_52 ;  
   wire _io_resp_bits_bridx_T_53 ;  
   wire _io_resp_bits_bridx_T_54 ;  
   wire _io_resp_bits_bridx_T_55 ;  
   wire _io_resp_bits_bridx_T_56 ;  
   wire _io_resp_bits_bridx_T_57 ;  
   wire _io_resp_bits_bridx_T_58 ;  
   wire _io_resp_bits_bridx_T_59 ;  
   wire _io_resp_bits_bridx_T_60 ;  
   wire _io_resp_bits_bridx_T_61 ;  
   wire _io_resp_bits_bridx_T_62 ;  
   wire _io_resp_bits_bridx_T_63 ;  
   wire _io_resp_bits_bridx_T_64 ;  
   wire _io_resp_bits_bridx_T_65 ;  
   wire _io_resp_bits_bridx_T_66 ;  
   wire _io_resp_bits_bridx_T_67 ;  
   wire _io_resp_bits_bridx_T_68 ;  
   wire _io_resp_bits_bridx_T_69 ;  
   wire _io_resp_bits_bridx_T_70 ;  
   wire _io_resp_bits_bridx_T_71 ;  
   wire _io_resp_bits_bridx_T_72 ;  
   wire _io_resp_bits_bridx_T_73 ;  
   wire _io_resp_bits_bridx_T_74 ;  
   wire _io_resp_bits_bridx_T_75 ;  
   wire _io_resp_bits_bridx_T_76 ;  
   wire _io_resp_bits_bridx_T_77 ;  
   wire _io_resp_bits_bridx_T_78 ;  
   wire _io_resp_bits_bridx_T_79 ;  
   wire _io_resp_bits_bridx_T_80 ;  
   wire _io_resp_bits_bridx_T_81 ;  
   wire leftOne ;  
   wire leftOne_1 ;  
   wire rightOne ;  
   wire rightOne_1 ;  
   wire rightTwo ;  
   wire leftOne_2 ;  
   wire _T_29 ;  
   wire leftTwo ;  
   wire leftOne_3 ;  
   wire rightOne_2 ;  
   wire leftOne_4 ;  
   wire leftTwo_1 ;  
   wire leftOne_5 ;  
   wire rightOne_3 ;  
   wire rightOne_4 ;  
   wire rightTwo_1 ;  
   wire rightOne_5 ;  
   wire _T_41 ;  
   wire _T_42 ;  
   wire rightTwo_2 ;  
   wire leftOne_6 ;  
   wire _T_43 ;  
   wire _T_44 ;  
   wire leftTwo_2 ;  
   wire leftOne_7 ;  
   wire leftOne_8 ;  
   wire rightOne_6 ;  
   wire rightOne_7 ;  
   wire rightTwo_3 ;  
   wire leftOne_9 ;  
   wire _T_54 ;  
   wire leftTwo_3 ;  
   wire leftOne_10 ;  
   wire rightOne_8 ;  
   wire leftOne_11 ;  
   wire leftTwo_4 ;  
   wire leftOne_12 ;  
   wire rightOne_9 ;  
   wire rightOne_10 ;  
   wire rightTwo_4 ;  
   wire rightOne_11 ;  
   wire _T_66 ;  
   wire _T_67 ;  
   wire rightTwo_5 ;  
   wire rightOne_12 ;  
   wire _T_68 ;  
   wire _T_69 ;  
   wire rightTwo_6 ;  
   wire leftOne_13 ;  
   wire _T_70 ;  
   wire _T_71 ;  
   wire leftTwo_5 ;  
   wire leftOne_14 ;  
   wire leftOne_15 ;  
   wire rightOne_13 ;  
   wire rightOne_14 ;  
   wire rightTwo_7 ;  
   wire leftOne_16 ;  
   wire _T_82 ;  
   wire leftTwo_6 ;  
   wire leftOne_17 ;  
   wire rightOne_15 ;  
   wire leftOne_18 ;  
   wire leftTwo_7 ;  
   wire leftOne_19 ;  
   wire rightOne_16 ;  
   wire rightOne_17 ;  
   wire rightTwo_8 ;  
   wire rightOne_18 ;  
   wire _T_94 ;  
   wire _T_95 ;  
   wire rightTwo_9 ;  
   wire leftOne_20 ;  
   wire _T_96 ;  
   wire _T_97 ;  
   wire leftTwo_8 ;  
   wire leftOne_21 ;  
   wire leftOne_22 ;  
   wire rightOne_19 ;  
   wire rightOne_20 ;  
   wire rightTwo_10 ;  
   wire leftOne_23 ;  
   wire _T_107 ;  
   wire leftTwo_9 ;  
   wire leftOne_24 ;  
   wire rightOne_21 ;  
   wire leftOne_25 ;  
   wire leftTwo_10 ;  
   wire leftOne_26 ;  
   wire rightOne_22 ;  
   wire rightOne_23 ;  
   wire rightTwo_11 ;  
   wire rightOne_24 ;  
   wire _T_119 ;  
   wire _T_120 ;  
   wire rightTwo_12 ;  
   wire rightOne_25 ;  
   wire _T_121 ;  
   wire _T_122 ;  
   wire rightTwo_13 ;  
   wire rightOne_26 ;  
   wire _T_123 ;  
   wire _T_124 ;  
   wire rightTwo_14 ;  
   wire _T_126 ;  
   wire _T_127 ;  
   wire _T_128 ;  
   wire [27:0] _isValid_T_5 ;  
   wire [31:0] _GEN_374 ;  
   wire [31:0] _GEN_375 ;  
   reg [7:0] history ;  
   reg [31:0] _RAND_188 ;  
   reg [9:0] reset_waddr ;  
   reg [31:0] _RAND_189 ;  
   wire resetting ;  
   wire [9:0] _reset_waddr_T_1 ;  
   wire [36:0] waddr_hi_13 ;  
   wire [8:0] _GEN_437 ;  
   wire [8:0] _waddr_T_30 ;  
   wire [15:0] _waddr_T_31 ;  
   wire [8:0] _waddr_T_33 ;  
   wire [8:0] _waddr_T_34 ;  
   wire [9:0] _GEN_383 ;  
   wire [9:0] _GEN_388 ;  
   wire [9:0] waddr_1 ;  
   wire _GEN_387 ;  
   wire _GEN_384 ;  
   wire _GEN_389 ;  
   wire isBranch_lo_lo_lo_lo ;  
   wire isBranch_lo_lo_lo_hi_lo ;  
   wire isBranch_lo_lo_lo_hi_hi ;  
   wire isBranch_lo_lo_hi_lo_lo ;  
   wire isBranch_lo_lo_hi_lo_hi ;  
   wire isBranch_lo_lo_hi_hi_lo ;  
   wire isBranch_lo_lo_hi_hi_hi ;  
   wire isBranch_lo_hi_lo_lo ;  
   wire isBranch_lo_hi_lo_hi_lo ;  
   wire isBranch_lo_hi_lo_hi_hi ;  
   wire isBranch_lo_hi_hi_lo_lo ;  
   wire isBranch_lo_hi_hi_lo_hi ;  
   wire isBranch_lo_hi_hi_hi_lo ;  
   wire isBranch_lo_hi_hi_hi_hi ;  
   wire isBranch_hi_lo_lo_lo ;  
   wire isBranch_hi_lo_lo_hi_lo ;  
   wire isBranch_hi_lo_lo_hi_hi ;  
   wire isBranch_hi_lo_hi_lo_lo ;  
   wire isBranch_hi_lo_hi_lo_hi ;  
   wire isBranch_hi_lo_hi_hi_lo ;  
   wire isBranch_hi_lo_hi_hi_hi ;  
   wire isBranch_hi_hi_lo_lo ;  
   wire isBranch_hi_hi_lo_hi_lo ;  
   wire isBranch_hi_hi_lo_hi_hi ;  
   wire isBranch_hi_hi_hi_lo_lo ;  
   wire isBranch_hi_hi_hi_lo_hi ;  
   wire isBranch_hi_hi_hi_hi_lo ;  
   wire isBranch_hi_hi_hi_hi_hi ;  
   wire [6:0] isBranch_lo_lo ;  
   wire [13:0] isBranch_lo ;  
   wire [6:0] isBranch_hi_lo ;  
   wire [27:0] _isBranch_T ;  
   wire [27:0] _isBranch_T_1 ;  
   wire isBranch ;  
   wire [36:0] res_res_value_hi ;  
   wire [8:0] _GEN_438 ;  
   wire [8:0] _res_res_value_T_3 ;  
   wire [15:0] _res_res_value_T_4 ;  
   wire [8:0] _res_res_value_T_6 ;  
   wire res_value ;  
   wire [6:0] history_lo ;  
   wire [7:0] _history_T ;  
   wire [6:0] history_lo_1 ;  
   wire [7:0] _history_T_1 ;  
   wire _T_134 ;  
   reg [2:0] count ;  
   reg [31:0] _RAND_190 ;  
   reg [2:0] pos ;  
   reg [31:0] _RAND_191 ;  
   reg [38:0] stack_0 ;  
   reg [63:0] _RAND_192 ;  
   reg [38:0] stack_1 ;  
   reg [63:0] _RAND_193 ;  
   reg [38:0] stack_2 ;  
   reg [63:0] _RAND_194 ;  
   reg [38:0] stack_3 ;  
   reg [63:0] _RAND_195 ;  
   reg [38:0] stack_4 ;  
   reg [63:0] _RAND_196 ;  
   reg [38:0] stack_5 ;  
   reg [63:0] _RAND_197 ;  
   wire doPeek_lo_lo_lo_lo ;  
   wire doPeek_lo_lo_lo_hi_lo ;  
   wire doPeek_lo_lo_lo_hi_hi ;  
   wire doPeek_lo_lo_hi_lo_lo ;  
   wire doPeek_lo_lo_hi_lo_hi ;  
   wire doPeek_lo_lo_hi_hi_lo ;  
   wire doPeek_lo_lo_hi_hi_hi ;  
   wire doPeek_lo_hi_lo_lo ;  
   wire doPeek_lo_hi_lo_hi_lo ;  
   wire doPeek_lo_hi_lo_hi_hi ;  
   wire doPeek_lo_hi_hi_lo_lo ;  
   wire doPeek_lo_hi_hi_lo_hi ;  
   wire doPeek_lo_hi_hi_hi_lo ;  
   wire doPeek_lo_hi_hi_hi_hi ;  
   wire doPeek_hi_lo_lo_lo ;  
   wire doPeek_hi_lo_lo_hi_lo ;  
   wire doPeek_hi_lo_lo_hi_hi ;  
   wire doPeek_hi_lo_hi_lo_lo ;  
   wire doPeek_hi_lo_hi_lo_hi ;  
   wire doPeek_hi_lo_hi_hi_lo ;  
   wire doPeek_hi_lo_hi_hi_hi ;  
   wire doPeek_hi_hi_lo_lo ;  
   wire doPeek_hi_hi_lo_hi_lo ;  
   wire doPeek_hi_hi_lo_hi_hi ;  
   wire doPeek_hi_hi_hi_lo_lo ;  
   wire doPeek_hi_hi_hi_lo_hi ;  
   wire doPeek_hi_hi_hi_hi_lo ;  
   wire doPeek_hi_hi_hi_hi_hi ;  
   wire [6:0] doPeek_lo_lo ;  
   wire [13:0] doPeek_lo ;  
   wire [6:0] doPeek_hi_lo ;  
   wire [27:0] _doPeek_T ;  
   wire [27:0] _doPeek_T_1 ;  
   wire doPeek ;  
   wire _io_ras_head_valid_T ;  
   wire [38:0] _GEN_397 ;  
   wire [38:0] _GEN_398 ;  
   wire [38:0] _GEN_399 ;  
   wire [38:0] _GEN_400 ;  
   wire [38:0] _GEN_401 ;  
   wire _T_137 ;  
   wire _T_138 ;  
   wire _T_139 ;  
   wire [2:0] _count_T_1 ;  
   wire _nextPos_T ;  
   wire [2:0] _nextPos_T_3 ;  
   wire [2:0] nextPos ;  
   wire _T_140 ;  
   wire [2:0] _count_T_3 ;  
   wire _pos_T ;  
   wire [2:0] _pos_T_3 ;  
   reg [19:0] BTB_state ;  
   reg [31:0] _RAND_198 ;  
   reg BTB_cov[0:1048575] ;  
   reg [31:0] _RAND_199 ;  
   wire BTB_cov_read_data ;  
   wire [19:0] BTB_cov_read_addr ;  
   wire BTB_cov_write_data ;  
   wire [19:0] BTB_cov_write_addr ;  
   wire BTB_cov_write_mask ;  
   wire BTB_cov_write_en ;  
   reg [29:0] BTB_covSum ;  
   reg [31:0] _RAND_200 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire mux_cond_4 ;  
   wire mux_cond_5 ;  
   wire mux_cond_6 ;  
   wire mux_cond_7 ;  
   wire mux_cond_8 ;  
   wire mux_cond_9 ;  
   wire mux_cond_10 ;  
   wire mux_cond_11 ;  
   wire mux_cond_12 ;  
   wire mux_cond_13 ;  
   wire mux_cond_14 ;  
   wire mux_cond_15 ;  
   wire mux_cond_16 ;  
   wire mux_cond_17 ;  
   wire mux_cond_18 ;  
   wire mux_cond_19 ;  
   wire mux_cond_20 ;  
   wire mux_cond_21 ;  
   wire mux_cond_22 ;  
   wire mux_cond_23 ;  
   wire mux_cond_24 ;  
   wire mux_cond_25 ;  
   wire mux_cond_26 ;  
   wire mux_cond_27 ;  
   wire mux_cond_28 ;  
   wire [9:0] nextPageRepl_shl ;  
   wire [19:0] nextPageRepl_pad ;  
   wire [3:0] r_respPipe_bits_taken_shl ;  
   wire [19:0] r_respPipe_bits_taken_pad ;  
   wire [16:0] r_btb_updatePipe_valid_shl ;  
   wire [19:0] r_btb_updatePipe_valid_pad ;  
   wire [14:0] count_shl ;  
   wire [19:0] count_pad ;  
   wire [13:0] r_respPipe_valid_shl ;  
   wire [19:0] r_respPipe_valid_pad ;  
   wire [3:0] pos_shl ;  
   wire [19:0] pos_pad ;  
   wire [13:0] pageValid_shl ;  
   wire [19:0] pageValid_pad ;  
   wire [17:0] r_btb_updatePipe_bits_isValid_shl ;  
   wire [19:0] r_btb_updatePipe_bits_isValid_pad ;  
   wire [14:0] mux_cond_0_shl ;  
   wire [19:0] mux_cond_0_pad ;  
   wire [17:0] mux_cond_1_shl ;  
   wire [19:0] mux_cond_1_pad ;  
   wire [3:0] mux_cond_2_shl ;  
   wire [19:0] mux_cond_2_pad ;  
   wire [17:0] mux_cond_3_shl ;  
   wire [19:0] mux_cond_3_pad ;  
   wire [13:0] mux_cond_4_shl ;  
   wire [19:0] mux_cond_4_pad ;  
   wire [3:0] mux_cond_5_shl ;  
   wire [19:0] mux_cond_5_pad ;  
   wire [1:0] mux_cond_6_shl ;  
   wire [19:0] mux_cond_6_pad ;  
   wire [13:0] mux_cond_7_shl ;  
   wire [19:0] mux_cond_7_pad ;  
   wire [16:0] mux_cond_8_shl ;  
   wire [19:0] mux_cond_8_pad ;  
   wire [3:0] mux_cond_9_shl ;  
   wire [19:0] mux_cond_9_pad ;  
   wire [9:0] mux_cond_10_shl ;  
   wire [19:0] mux_cond_10_pad ;  
   wire [3:0] mux_cond_11_shl ;  
   wire [19:0] mux_cond_11_pad ;  
   wire [17:0] mux_cond_12_shl ;  
   wire [19:0] mux_cond_12_pad ;  
   wire [8:0] mux_cond_13_shl ;  
   wire [19:0] mux_cond_13_pad ;  
   wire [4:0] mux_cond_14_shl ;  
   wire [19:0] mux_cond_14_pad ;  
   wire [11:0] mux_cond_15_shl ;  
   wire [19:0] mux_cond_15_pad ;  
   wire [12:0] mux_cond_16_shl ;  
   wire [19:0] mux_cond_16_pad ;  
   wire [5:0] mux_cond_17_shl ;  
   wire [19:0] mux_cond_17_pad ;  
   wire mux_cond_18_shl ;  
   wire [19:0] mux_cond_18_pad ;  
   wire [1:0] mux_cond_19_shl ;  
   wire [19:0] mux_cond_19_pad ;  
   wire [2:0] mux_cond_20_shl ;  
   wire [19:0] mux_cond_20_pad ;  
   wire [5:0] mux_cond_21_shl ;  
   wire [19:0] mux_cond_21_pad ;  
   wire [16:0] mux_cond_22_shl ;  
   wire [19:0] mux_cond_22_pad ;  
   wire [13:0] mux_cond_23_shl ;  
   wire [19:0] mux_cond_23_pad ;  
   wire [19:0] mux_cond_24_shl ;  
   wire [19:0] mux_cond_24_pad ;  
   wire [14:0] mux_cond_25_shl ;  
   wire [19:0] mux_cond_25_pad ;  
   wire [8:0] mux_cond_26_shl ;  
   wire [19:0] mux_cond_26_pad ;  
   wire [18:0] mux_cond_27_shl ;  
   wire [19:0] mux_cond_27_pad ;  
   wire [5:0] mux_cond_28_shl ;  
   wire [19:0] mux_cond_28_pad ;  
   wire [12:0] cfiType_17_shl ;  
   wire [19:0] cfiType_17_pad ;  
   wire [12:0] cfiType_22_shl ;  
   wire [19:0] cfiType_22_pad ;  
   wire [12:0] cfiType_21_shl ;  
   wire [19:0] cfiType_21_pad ;  
   wire [17:0] tgtPages_4_shl ;  
   wire [19:0] tgtPages_4_pad ;  
   wire [17:0] tgtPages_6_shl ;  
   wire [19:0] tgtPages_6_pad ;  
   wire [17:0] tgtPages_11_shl ;  
   wire [19:0] tgtPages_11_pad ;  
   wire [17:0] tgtPages_7_shl ;  
   wire [19:0] tgtPages_7_pad ;  
   wire [17:0] tgtPages_20_shl ;  
   wire [19:0] tgtPages_20_pad ;  
   wire [12:0] cfiType_3_shl ;  
   wire [19:0] cfiType_3_pad ;  
   wire [17:0] tgtPages_16_shl ;  
   wire [19:0] tgtPages_16_pad ;  
   wire [12:0] cfiType_24_shl ;  
   wire [19:0] cfiType_24_pad ;  
   wire [17:0] tgtPages_17_shl ;  
   wire [19:0] tgtPages_17_pad ;  
   wire [12:0] cfiType_6_shl ;  
   wire [19:0] cfiType_6_pad ;  
   wire [17:0] tgtPages_9_shl ;  
   wire [19:0] tgtPages_9_pad ;  
   wire [17:0] tgtPages_2_shl ;  
   wire [19:0] tgtPages_2_pad ;  
   wire [12:0] cfiType_10_shl ;  
   wire [19:0] cfiType_10_pad ;  
   wire [17:0] tgtPages_18_shl ;  
   wire [19:0] tgtPages_18_pad ;  
   wire [17:0] tgtPages_0_shl ;  
   wire [19:0] tgtPages_0_pad ;  
   wire [17:0] tgtPages_25_shl ;  
   wire [19:0] tgtPages_25_pad ;  
   wire [17:0] tgtPages_22_shl ;  
   wire [19:0] tgtPages_22_pad ;  
   wire [12:0] cfiType_5_shl ;  
   wire [19:0] cfiType_5_pad ;  
   wire [12:0] cfiType_12_shl ;  
   wire [19:0] cfiType_12_pad ;  
   wire [12:0] cfiType_18_shl ;  
   wire [19:0] cfiType_18_pad ;  
   wire [17:0] tgtPages_24_shl ;  
   wire [19:0] tgtPages_24_pad ;  
   wire [17:0] tgtPages_26_shl ;  
   wire [19:0] tgtPages_26_pad ;  
   wire [17:0] tgtPages_1_shl ;  
   wire [19:0] tgtPages_1_pad ;  
   wire [17:0] tgtPages_10_shl ;  
   wire [19:0] tgtPages_10_pad ;  
   wire [12:0] cfiType_25_shl ;  
   wire [19:0] cfiType_25_pad ;  
   wire [12:0] cfiType_16_shl ;  
   wire [19:0] cfiType_16_pad ;  
   wire [17:0] tgtPages_13_shl ;  
   wire [19:0] tgtPages_13_pad ;  
   wire [12:0] cfiType_19_shl ;  
   wire [19:0] cfiType_19_pad ;  
   wire [12:0] cfiType_2_shl ;  
   wire [19:0] cfiType_2_pad ;  
   wire [12:0] cfiType_20_shl ;  
   wire [19:0] cfiType_20_pad ;  
   wire [17:0] tgtPages_15_shl ;  
   wire [19:0] tgtPages_15_pad ;  
   wire [17:0] tgtPages_8_shl ;  
   wire [19:0] tgtPages_8_pad ;  
   wire [17:0] tgtPages_5_shl ;  
   wire [19:0] tgtPages_5_pad ;  
   wire [12:0] cfiType_0_shl ;  
   wire [19:0] cfiType_0_pad ;  
   wire [17:0] tgtPages_3_shl ;  
   wire [19:0] tgtPages_3_pad ;  
   wire [17:0] tgtPages_27_shl ;  
   wire [19:0] tgtPages_27_pad ;  
   wire [12:0] cfiType_27_shl ;  
   wire [19:0] cfiType_27_pad ;  
   wire [17:0] tgtPages_14_shl ;  
   wire [19:0] tgtPages_14_pad ;  
   wire [12:0] cfiType_13_shl ;  
   wire [19:0] cfiType_13_pad ;  
   wire [12:0] cfiType_23_shl ;  
   wire [19:0] cfiType_23_pad ;  
   wire [12:0] cfiType_4_shl ;  
   wire [19:0] cfiType_4_pad ;  
   wire [12:0] cfiType_1_shl ;  
   wire [19:0] cfiType_1_pad ;  
   wire [17:0] tgtPages_21_shl ;  
   wire [19:0] tgtPages_21_pad ;  
   wire [12:0] cfiType_8_shl ;  
   wire [19:0] cfiType_8_pad ;  
   wire [17:0] tgtPages_23_shl ;  
   wire [19:0] tgtPages_23_pad ;  
   wire [17:0] tgtPages_19_shl ;  
   wire [19:0] tgtPages_19_pad ;  
   wire [12:0] cfiType_11_shl ;  
   wire [19:0] cfiType_11_pad ;  
   wire [17:0] tgtPages_12_shl ;  
   wire [19:0] tgtPages_12_pad ;  
   wire [12:0] cfiType_9_shl ;  
   wire [19:0] cfiType_9_pad ;  
   wire [12:0] cfiType_14_shl ;  
   wire [19:0] cfiType_14_pad ;  
   wire [12:0] cfiType_7_shl ;  
   wire [19:0] cfiType_7_pad ;  
   wire [12:0] cfiType_26_shl ;  
   wire [19:0] cfiType_26_pad ;  
   wire [12:0] cfiType_15_shl ;  
   wire [19:0] cfiType_15_pad ;  
   wire [19:0] BTB_xor31 ;  
   wire [19:0] BTB_xor66 ;  
   wire [19:0] BTB_xor32 ;  
   wire [19:0] BTB_xor15 ;  
   wire [19:0] BTB_xor68 ;  
   wire [19:0] BTB_xor33 ;  
   wire [19:0] BTB_xor70 ;  
   wire [19:0] BTB_xor34 ;  
   wire [19:0] BTB_xor16 ;  
   wire [19:0] BTB_xor7 ;  
   wire [19:0] BTB_xor72 ;  
   wire [19:0] BTB_xor35 ;  
   wire [19:0] BTB_xor74 ;  
   wire [19:0] BTB_xor36 ;  
   wire [19:0] BTB_xor17 ;  
   wire [19:0] BTB_xor76 ;  
   wire [19:0] BTB_xor37 ;  
   wire [19:0] BTB_xor78 ;  
   wire [19:0] BTB_xor38 ;  
   wire [19:0] BTB_xor18 ;  
   wire [19:0] BTB_xor8 ;  
   wire [19:0] BTB_xor3 ;  
   wire [19:0] BTB_xor39 ;  
   wire [19:0] BTB_xor82 ;  
   wire [19:0] BTB_xor40 ;  
   wire [19:0] BTB_xor19 ;  
   wire [19:0] BTB_xor84 ;  
   wire [19:0] BTB_xor41 ;  
   wire [19:0] BTB_xor86 ;  
   wire [19:0] BTB_xor42 ;  
   wire [19:0] BTB_xor20 ;  
   wire [19:0] BTB_xor9 ;  
   wire [19:0] BTB_xor88 ;  
   wire [19:0] BTB_xor43 ;  
   wire [19:0] BTB_xor90 ;  
   wire [19:0] BTB_xor44 ;  
   wire [19:0] BTB_xor21 ;  
   wire [19:0] BTB_xor92 ;  
   wire [19:0] BTB_xor45 ;  
   wire [19:0] BTB_xor94 ;  
   wire [19:0] BTB_xor46 ;  
   wire [19:0] BTB_xor22 ;  
   wire [19:0] BTB_xor10 ;  
   wire [19:0] BTB_xor4 ;  
   wire [19:0] BTB_xor1 ;  
   wire [19:0] BTB_xor47 ;  
   wire [19:0] BTB_xor98 ;  
   wire [19:0] BTB_xor48 ;  
   wire [19:0] BTB_xor23 ;  
   wire [19:0] BTB_xor100 ;  
   wire [19:0] BTB_xor49 ;  
   wire [19:0] BTB_xor102 ;  
   wire [19:0] BTB_xor50 ;  
   wire [19:0] BTB_xor24 ;  
   wire [19:0] BTB_xor11 ;  
   wire [19:0] BTB_xor104 ;  
   wire [19:0] BTB_xor51 ;  
   wire [19:0] BTB_xor106 ;  
   wire [19:0] BTB_xor52 ;  
   wire [19:0] BTB_xor25 ;  
   wire [19:0] BTB_xor108 ;  
   wire [19:0] BTB_xor53 ;  
   wire [19:0] BTB_xor110 ;  
   wire [19:0] BTB_xor54 ;  
   wire [19:0] BTB_xor26 ;  
   wire [19:0] BTB_xor12 ;  
   wire [19:0] BTB_xor5 ;  
   wire [19:0] BTB_xor112 ;  
   wire [19:0] BTB_xor55 ;  
   wire [19:0] BTB_xor114 ;  
   wire [19:0] BTB_xor56 ;  
   wire [19:0] BTB_xor27 ;  
   wire [19:0] BTB_xor116 ;  
   wire [19:0] BTB_xor57 ;  
   wire [19:0] BTB_xor118 ;  
   wire [19:0] BTB_xor58 ;  
   wire [19:0] BTB_xor28 ;  
   wire [19:0] BTB_xor13 ;  
   wire [19:0] BTB_xor120 ;  
   wire [19:0] BTB_xor59 ;  
   wire [19:0] BTB_xor122 ;  
   wire [19:0] BTB_xor60 ;  
   wire [19:0] BTB_xor29 ;  
   wire [19:0] BTB_xor124 ;  
   wire [19:0] BTB_xor61 ;  
   wire [19:0] BTB_xor126 ;  
   wire [19:0] BTB_xor62 ;  
   wire [19:0] BTB_xor30 ;  
   wire [19:0] BTB_xor14 ;  
   wire [19:0] BTB_xor6 ;  
   wire [19:0] BTB_xor2 ;  
   wire [19:0] BTB_xor0 ;  
  assign table__res_res_value_MPORT_addr=_res_res_value_T_3^_res_res_value_T_6; 
  assign table__res_res_value_MPORT_data=table_[table__res_res_value_MPORT_addr]; 
  assign table__MPORT_data=io_bht_update_valid&_GEN_389; 
  assign table__MPORT_addr=waddr_1[8:0]; 
  assign table__MPORT_mask=1'h1; 
  assign table__MPORT_en=io_bht_update_valid ? _GEN_387:resetting; 
  assign pagesMasked_0=pageValid[0] ? pages_0:25'h0; 
  assign pagesMasked_1=pageValid[1] ? pages_1:25'h0; 
  assign pagesMasked_2=pageValid[2] ? pages_2:25'h0; 
  assign pagesMasked_3=pageValid[3] ? pages_3:25'h0; 
  assign pagesMasked_4=pageValid[4] ? pages_4:25'h0; 
  assign pagesMasked_5=pageValid[5] ? pages_5:25'h0; 
  assign pageHit_p=io_req_bits_addr[38:14]; 
  assign pageHit_lo_lo=pages_0==pageHit_p; 
  assign pageHit_lo_hi_lo=pages_1==pageHit_p; 
  assign pageHit_lo_hi_hi=pages_2==pageHit_p; 
  assign pageHit_hi_lo=pages_3==pageHit_p; 
  assign pageHit_hi_hi_lo=pages_4==pageHit_p; 
  assign pageHit_hi_hi_hi=pages_5==pageHit_p; 
  assign _pageHit_T={pageHit_hi_hi_hi,pageHit_hi_hi_lo,pageHit_hi_lo,pageHit_lo_hi_hi,pageHit_lo_hi_lo,pageHit_lo_lo}; 
  assign pageHit=pageValid&_pageHit_T; 
  assign idxHit_idx=io_req_bits_addr[13:1]; 
  assign idxHit_lo_lo_lo_lo=idxs_0==idxHit_idx; 
  assign idxHit_lo_lo_lo_hi_lo=idxs_1==idxHit_idx; 
  assign idxHit_lo_lo_lo_hi_hi=idxs_2==idxHit_idx; 
  assign idxHit_lo_lo_hi_lo_lo=idxs_3==idxHit_idx; 
  assign idxHit_lo_lo_hi_lo_hi=idxs_4==idxHit_idx; 
  assign idxHit_lo_lo_hi_hi_lo=idxs_5==idxHit_idx; 
  assign idxHit_lo_lo_hi_hi_hi=idxs_6==idxHit_idx; 
  assign idxHit_lo_hi_lo_lo=idxs_7==idxHit_idx; 
  assign idxHit_lo_hi_lo_hi_lo=idxs_8==idxHit_idx; 
  assign idxHit_lo_hi_lo_hi_hi=idxs_9==idxHit_idx; 
  assign idxHit_lo_hi_hi_lo_lo=idxs_10==idxHit_idx; 
  assign idxHit_lo_hi_hi_lo_hi=idxs_11==idxHit_idx; 
  assign idxHit_lo_hi_hi_hi_lo=idxs_12==idxHit_idx; 
  assign idxHit_lo_hi_hi_hi_hi=idxs_13==idxHit_idx; 
  assign idxHit_hi_lo_lo_lo=idxs_14==idxHit_idx; 
  assign idxHit_hi_lo_lo_hi_lo=idxs_15==idxHit_idx; 
  assign idxHit_hi_lo_lo_hi_hi=idxs_16==idxHit_idx; 
  assign idxHit_hi_lo_hi_lo_lo=idxs_17==idxHit_idx; 
  assign idxHit_hi_lo_hi_lo_hi=idxs_18==idxHit_idx; 
  assign idxHit_hi_lo_hi_hi_lo=idxs_19==idxHit_idx; 
  assign idxHit_hi_lo_hi_hi_hi=idxs_20==idxHit_idx; 
  assign idxHit_hi_hi_lo_lo=idxs_21==idxHit_idx; 
  assign idxHit_hi_hi_lo_hi_lo=idxs_22==idxHit_idx; 
  assign idxHit_hi_hi_lo_hi_hi=idxs_23==idxHit_idx; 
  assign idxHit_hi_hi_hi_lo_lo=idxs_24==idxHit_idx; 
  assign idxHit_hi_hi_hi_lo_hi=idxs_25==idxHit_idx; 
  assign idxHit_hi_hi_hi_hi_lo=idxs_26==idxHit_idx; 
  assign idxHit_hi_hi_hi_hi_hi=idxs_27==idxHit_idx; 
  assign idxHit_lo_lo={idxHit_lo_lo_hi_hi_hi,idxHit_lo_lo_hi_hi_lo,idxHit_lo_lo_hi_lo_hi,idxHit_lo_lo_hi_lo_lo,idxHit_lo_lo_lo_hi_hi,idxHit_lo_lo_lo_hi_lo,idxHit_lo_lo_lo_lo}; 
  assign idxHit_lo={idxHit_lo_hi_hi_hi_hi,idxHit_lo_hi_hi_hi_lo,idxHit_lo_hi_hi_lo_hi,idxHit_lo_hi_hi_lo_lo,idxHit_lo_hi_lo_hi_hi,idxHit_lo_hi_lo_hi_lo,idxHit_lo_hi_lo_lo,idxHit_lo_lo}; 
  assign idxHit_hi_lo={idxHit_hi_lo_hi_hi_hi,idxHit_hi_lo_hi_hi_lo,idxHit_hi_lo_hi_lo_hi,idxHit_hi_lo_hi_lo_lo,idxHit_hi_lo_lo_hi_hi,idxHit_hi_lo_lo_hi_lo,idxHit_hi_lo_lo_lo}; 
  assign _idxHit_T={idxHit_hi_hi_hi_hi_hi,idxHit_hi_hi_hi_hi_lo,idxHit_hi_hi_hi_lo_hi,idxHit_hi_hi_hi_lo_lo,idxHit_hi_hi_lo_hi_hi,idxHit_hi_hi_lo_hi_lo,idxHit_hi_hi_lo_lo,idxHit_hi_lo,idxHit_lo}; 
  assign idxHit=_idxHit_T&isValid; 
  assign updatePageHit_p=r_btb_updatePipe_bits_pc[38:14]; 
  assign updatePageHit_lo_lo=pages_0==updatePageHit_p; 
  assign updatePageHit_lo_hi_lo=pages_1==updatePageHit_p; 
  assign updatePageHit_lo_hi_hi=pages_2==updatePageHit_p; 
  assign updatePageHit_hi_lo=pages_3==updatePageHit_p; 
  assign updatePageHit_hi_hi_lo=pages_4==updatePageHit_p; 
  assign updatePageHit_hi_hi_hi=pages_5==updatePageHit_p; 
  assign _updatePageHit_T={updatePageHit_hi_hi_hi,updatePageHit_hi_hi_lo,updatePageHit_hi_lo,updatePageHit_lo_hi_hi,updatePageHit_lo_hi_lo,updatePageHit_lo_lo}; 
  assign updatePageHit=pageValid&_updatePageHit_T; 
  assign updateHit=r_btb_updatePipe_bits_prediction_entry<5'h1c; 
  assign useUpdatePageHit=|updatePageHit; 
  assign usePageHit=|pageHit; 
  assign doIdxPageRepl=~useUpdatePageHit; 
  assign idxPageRepl_hi=pageHit[4:0]; 
  assign idxPageRepl_lo=pageHit[5]; 
  assign _idxPageRepl_T={idxPageRepl_hi,idxPageRepl_lo}; 
  assign _idxPageRepl_T_1=8'h1<<nextPageRepl; 
  assign _idxPageRepl_T_2=usePageHit ? 8'h0:_idxPageRepl_T_1; 
  assign _GEN_430={2'b0,_idxPageRepl_T}; 
  assign idxPageRepl=_GEN_430|_idxPageRepl_T_2; 
  assign idxPageUpdateOH=useUpdatePageHit ? {2'b0,updatePageHit}:idxPageRepl; 
  assign idxPageUpdate_hi=idxPageUpdateOH[7:4]; 
  assign idxPageUpdate_lo=idxPageUpdateOH[3:0]; 
  assign idxPageUpdate_hi_1=|idxPageUpdate_hi; 
  assign _idxPageUpdate_T=idxPageUpdate_hi|idxPageUpdate_lo; 
  assign idxPageUpdate_hi_2=_idxPageUpdate_T[3:2]; 
  assign idxPageUpdate_lo_1=_idxPageUpdate_T[1:0]; 
  assign idxPageUpdate_hi_3=|idxPageUpdate_hi_2; 
  assign _idxPageUpdate_T_1=idxPageUpdate_hi_2|idxPageUpdate_lo_1; 
  assign idxPageUpdate_lo_2=_idxPageUpdate_T_1[1]; 
  assign idxPageUpdate={idxPageUpdate_hi_1,idxPageUpdate_hi_3,idxPageUpdate_lo_2}; 
  assign idxPageReplEn=doIdxPageRepl ? idxPageRepl:8'h0; 
  assign samePage=updatePageHit_p==pageHit_p; 
  assign doTgtPageRepl=~samePage&~usePageHit; 
  assign tgtPageRepl_hi=idxPageUpdateOH[4:0]; 
  assign tgtPageRepl_lo=idxPageUpdateOH[5]; 
  assign _tgtPageRepl_T={tgtPageRepl_hi,tgtPageRepl_lo}; 
  assign tgtPageRepl=samePage ? idxPageUpdateOH:{2'b0,_tgtPageRepl_T}; 
  assign _tgtPageUpdate_T=usePageHit ? 8'h0:tgtPageRepl; 
  assign _GEN_431={2'b0,pageHit}; 
  assign _tgtPageUpdate_T_1=_GEN_431|_tgtPageUpdate_T; 
  assign tgtPageUpdate_hi=_tgtPageUpdate_T_1[7:4]; 
  assign tgtPageUpdate_lo=_tgtPageUpdate_T_1[3:0]; 
  assign tgtPageUpdate_hi_1=|tgtPageUpdate_hi; 
  assign _tgtPageUpdate_T_2=tgtPageUpdate_hi|tgtPageUpdate_lo; 
  assign tgtPageUpdate_hi_2=_tgtPageUpdate_T_2[3:2]; 
  assign tgtPageUpdate_lo_1=_tgtPageUpdate_T_2[1:0]; 
  assign tgtPageUpdate_hi_3=|tgtPageUpdate_hi_2; 
  assign _tgtPageUpdate_T_3=tgtPageUpdate_hi_2|tgtPageUpdate_lo_1; 
  assign tgtPageUpdate_lo_2=_tgtPageUpdate_T_3[1]; 
  assign tgtPageUpdate={tgtPageUpdate_hi_1,tgtPageUpdate_hi_3,tgtPageUpdate_lo_2}; 
  assign tgtPageReplEn=doTgtPageRepl ? tgtPageRepl:8'h0; 
  assign _T=doIdxPageRepl|doTgtPageRepl; 
  assign _T_1=r_btb_updatePipe_valid&_T; 
  assign both=doIdxPageRepl&doTgtPageRepl; 
  assign _next_T=both ? 2'h2:2'h1; 
  assign _GEN_432={1'b0,_next_T}; 
  assign next=nextPageRepl+_GEN_432; 
  assign _nextPageRepl_T=next>=3'h6; 
  assign waddr_hi=state_reg[26]; 
  assign waddr_left_subtree_state=state_reg[25:15]; 
  assign waddr_right_subtree_state=state_reg[14:0]; 
  assign waddr_hi_1=waddr_left_subtree_state[10]; 
  assign waddr_left_subtree_state_1=waddr_left_subtree_state[9:7]; 
  assign waddr_right_subtree_state_1=waddr_left_subtree_state[6:0]; 
  assign waddr_hi_2=waddr_left_subtree_state_1[2]; 
  assign waddr_left_subtree_state_2=waddr_left_subtree_state_1[1]; 
  assign waddr_right_subtree_state_2=waddr_left_subtree_state_1[0]; 
  assign waddr_lo=waddr_hi_2 ? waddr_left_subtree_state_2:waddr_right_subtree_state_2; 
  assign _waddr_T_2={waddr_hi_2,waddr_lo}; 
  assign waddr_hi_3=waddr_right_subtree_state_1[6]; 
  assign waddr_left_subtree_state_3=waddr_right_subtree_state_1[5:3]; 
  assign waddr_right_subtree_state_3=waddr_right_subtree_state_1[2:0]; 
  assign waddr_hi_4=waddr_left_subtree_state_3[2]; 
  assign waddr_left_subtree_state_4=waddr_left_subtree_state_3[1]; 
  assign waddr_right_subtree_state_4=waddr_left_subtree_state_3[0]; 
  assign waddr_lo_1=waddr_hi_4 ? waddr_left_subtree_state_4:waddr_right_subtree_state_4; 
  assign _waddr_T_5={waddr_hi_4,waddr_lo_1}; 
  assign waddr_hi_5=waddr_right_subtree_state_3[2]; 
  assign waddr_left_subtree_state_5=waddr_right_subtree_state_3[1]; 
  assign waddr_right_subtree_state_5=waddr_right_subtree_state_3[0]; 
  assign waddr_lo_2=waddr_hi_5 ? waddr_left_subtree_state_5:waddr_right_subtree_state_5; 
  assign _waddr_T_8={waddr_hi_5,waddr_lo_2}; 
  assign waddr_lo_3=waddr_hi_3 ? _waddr_T_5:_waddr_T_8; 
  assign _waddr_T_9={waddr_hi_3,waddr_lo_3}; 
  assign waddr_lo_4=waddr_hi_1 ? {1'b0,_waddr_T_2}:_waddr_T_9; 
  assign _waddr_T_10={waddr_hi_1,waddr_lo_4}; 
  assign waddr_hi_6=waddr_right_subtree_state[14]; 
  assign waddr_left_subtree_state_6=waddr_right_subtree_state[13:7]; 
  assign waddr_right_subtree_state_6=waddr_right_subtree_state[6:0]; 
  assign waddr_hi_7=waddr_left_subtree_state_6[6]; 
  assign waddr_left_subtree_state_7=waddr_left_subtree_state_6[5:3]; 
  assign waddr_right_subtree_state_7=waddr_left_subtree_state_6[2:0]; 
  assign waddr_hi_8=waddr_left_subtree_state_7[2]; 
  assign waddr_left_subtree_state_8=waddr_left_subtree_state_7[1]; 
  assign waddr_right_subtree_state_8=waddr_left_subtree_state_7[0]; 
  assign waddr_lo_5=waddr_hi_8 ? waddr_left_subtree_state_8:waddr_right_subtree_state_8; 
  assign _waddr_T_13={waddr_hi_8,waddr_lo_5}; 
  assign waddr_hi_9=waddr_right_subtree_state_7[2]; 
  assign waddr_left_subtree_state_9=waddr_right_subtree_state_7[1]; 
  assign waddr_right_subtree_state_9=waddr_right_subtree_state_7[0]; 
  assign waddr_lo_6=waddr_hi_9 ? waddr_left_subtree_state_9:waddr_right_subtree_state_9; 
  assign _waddr_T_16={waddr_hi_9,waddr_lo_6}; 
  assign waddr_lo_7=waddr_hi_7 ? _waddr_T_13:_waddr_T_16; 
  assign _waddr_T_17={waddr_hi_7,waddr_lo_7}; 
  assign waddr_hi_10=waddr_right_subtree_state_6[6]; 
  assign waddr_left_subtree_state_10=waddr_right_subtree_state_6[5:3]; 
  assign waddr_right_subtree_state_10=waddr_right_subtree_state_6[2:0]; 
  assign waddr_hi_11=waddr_left_subtree_state_10[2]; 
  assign waddr_left_subtree_state_11=waddr_left_subtree_state_10[1]; 
  assign waddr_right_subtree_state_11=waddr_left_subtree_state_10[0]; 
  assign waddr_lo_8=waddr_hi_11 ? waddr_left_subtree_state_11:waddr_right_subtree_state_11; 
  assign _waddr_T_20={waddr_hi_11,waddr_lo_8}; 
  assign waddr_hi_12=waddr_right_subtree_state_10[2]; 
  assign waddr_left_subtree_state_12=waddr_right_subtree_state_10[1]; 
  assign waddr_right_subtree_state_12=waddr_right_subtree_state_10[0]; 
  assign waddr_lo_9=waddr_hi_12 ? waddr_left_subtree_state_12:waddr_right_subtree_state_12; 
  assign _waddr_T_23={waddr_hi_12,waddr_lo_9}; 
  assign waddr_lo_10=waddr_hi_10 ? _waddr_T_20:_waddr_T_23; 
  assign _waddr_T_24={waddr_hi_10,waddr_lo_10}; 
  assign waddr_lo_11=waddr_hi_6 ? _waddr_T_17:_waddr_T_24; 
  assign _waddr_T_25={waddr_hi_6,waddr_lo_11}; 
  assign waddr_lo_12=waddr_hi ? _waddr_T_10:_waddr_T_25; 
  assign _waddr_T_26={waddr_hi,waddr_lo_12}; 
  assign waddr=updateHit ? r_btb_updatePipe_bits_prediction_entry:_waddr_T_26; 
  assign _T_2=r_respPipe_valid&r_respPipe_bits_taken; 
  assign _T_3=_T_2|r_btb_updatePipe_valid; 
  assign state_reg_touch_way_sized=r_btb_updatePipe_valid ? waddr:r_respPipe_bits_entry; 
  assign state_reg_hi_hi=~state_reg_touch_way_sized[4]; 
  assign state_reg_hi_hi_1=~state_reg_touch_way_sized[3]; 
  assign state_reg_hi_hi_2=~state_reg_touch_way_sized[1]; 
  assign state_reg_hi_lo=state_reg_hi_hi_2 ? waddr_left_subtree_state_2:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo=state_reg_hi_hi_2 ? ~state_reg_touch_way_sized[0]:waddr_right_subtree_state_2; 
  assign _state_reg_T_8={state_reg_hi_hi_2,state_reg_hi_lo,state_reg_lo}; 
  assign state_reg_hi_lo_1=state_reg_hi_hi_1 ? waddr_left_subtree_state_1:_state_reg_T_8; 
  assign state_reg_hi_hi_3=~state_reg_touch_way_sized[2]; 
  assign state_reg_hi_hi_4=~state_reg_touch_way_sized[1]; 
  assign state_reg_hi_lo_2=state_reg_hi_hi_4 ? waddr_left_subtree_state_4:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo_1=state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0]:waddr_right_subtree_state_4; 
  assign _state_reg_T_17={state_reg_hi_hi_4,state_reg_hi_lo_2,state_reg_lo_1}; 
  assign state_reg_hi_lo_3=state_reg_hi_hi_3 ? waddr_left_subtree_state_3:_state_reg_T_17; 
  assign state_reg_hi_lo_4=state_reg_hi_hi_4 ? waddr_left_subtree_state_5:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo_2=state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0]:waddr_right_subtree_state_5; 
  assign _state_reg_T_25={state_reg_hi_hi_4,state_reg_hi_lo_4,state_reg_lo_2}; 
  assign state_reg_lo_3=state_reg_hi_hi_3 ? _state_reg_T_25:waddr_right_subtree_state_3; 
  assign _state_reg_T_26={state_reg_hi_hi_3,state_reg_hi_lo_3,state_reg_lo_3}; 
  assign state_reg_lo_4=state_reg_hi_hi_1 ? _state_reg_T_26:waddr_right_subtree_state_1; 
  assign _state_reg_T_27={state_reg_hi_hi_1,state_reg_hi_lo_1,state_reg_lo_4}; 
  assign state_reg_hi_lo_5=state_reg_hi_hi ? waddr_left_subtree_state:_state_reg_T_27; 
  assign state_reg_hi_lo_6=state_reg_hi_hi_4 ? waddr_left_subtree_state_8:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo_5=state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0]:waddr_right_subtree_state_8; 
  assign _state_reg_T_37={state_reg_hi_hi_4,state_reg_hi_lo_6,state_reg_lo_5}; 
  assign state_reg_hi_lo_7=state_reg_hi_hi_3 ? waddr_left_subtree_state_7:_state_reg_T_37; 
  assign state_reg_hi_lo_8=state_reg_hi_hi_4 ? waddr_left_subtree_state_9:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo_6=state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0]:waddr_right_subtree_state_9; 
  assign _state_reg_T_45={state_reg_hi_hi_4,state_reg_hi_lo_8,state_reg_lo_6}; 
  assign state_reg_lo_7=state_reg_hi_hi_3 ? _state_reg_T_45:waddr_right_subtree_state_7; 
  assign _state_reg_T_46={state_reg_hi_hi_3,state_reg_hi_lo_7,state_reg_lo_7}; 
  assign state_reg_hi_lo_9=state_reg_hi_hi_1 ? waddr_left_subtree_state_6:_state_reg_T_46; 
  assign state_reg_hi_lo_10=state_reg_hi_hi_4 ? waddr_left_subtree_state_11:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo_8=state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0]:waddr_right_subtree_state_11; 
  assign _state_reg_T_55={state_reg_hi_hi_4,state_reg_hi_lo_10,state_reg_lo_8}; 
  assign state_reg_hi_lo_11=state_reg_hi_hi_3 ? waddr_left_subtree_state_10:_state_reg_T_55; 
  assign state_reg_hi_lo_12=state_reg_hi_hi_4 ? waddr_left_subtree_state_12:~state_reg_touch_way_sized[0]; 
  assign state_reg_lo_9=state_reg_hi_hi_4 ? ~state_reg_touch_way_sized[0]:waddr_right_subtree_state_12; 
  assign _state_reg_T_63={state_reg_hi_hi_4,state_reg_hi_lo_12,state_reg_lo_9}; 
  assign state_reg_lo_10=state_reg_hi_hi_3 ? _state_reg_T_63:waddr_right_subtree_state_10; 
  assign _state_reg_T_64={state_reg_hi_hi_3,state_reg_hi_lo_11,state_reg_lo_10}; 
  assign state_reg_lo_11=state_reg_hi_hi_1 ? _state_reg_T_64:waddr_right_subtree_state_6; 
  assign _state_reg_T_65={state_reg_hi_hi_1,state_reg_hi_lo_9,state_reg_lo_11}; 
  assign state_reg_lo_12=state_reg_hi_hi ? _state_reg_T_65:waddr_right_subtree_state; 
  assign _state_reg_T_66={state_reg_hi_hi,state_reg_hi_lo_5,state_reg_lo_12}; 
  assign mask=32'h1<<waddr; 
  assign _idxPages_T=idxPageUpdate+3'h1; 
  assign _GEN_433={4'b0,isValid}; 
  assign _isValid_T=_GEN_433|mask; 
  assign _isValid_T_2=_GEN_433&~mask; 
  assign _isValid_T_3=r_btb_updatePipe_bits_isValid ? _isValid_T:_isValid_T_2; 
  assign idxWritesEven=~idxPageUpdate[0]; 
  assign _T_5=idxWritesEven ? idxPageReplEn:tgtPageReplEn; 
  assign _T_12=idxWritesEven ? tgtPageReplEn:idxPageReplEn; 
  assign _GEN_435={2'b0,pageValid}; 
  assign _pageValid_T=_GEN_435|tgtPageReplEn; 
  assign _pageValid_T_1=_pageValid_T|idxPageReplEn; 
  assign _GEN_338=r_btb_updatePipe_valid ? _isValid_T_3:{4'b0,isValid}; 
  assign _GEN_373=r_btb_updatePipe_valid ? _pageValid_T_1:{2'b0,pageValid}; 
  assign _io_resp_valid_T={pageHit,1'h0}; 
  assign _io_resp_valid_T_29=idxHit[0] ? idxPages_0:3'h0; 
  assign _io_resp_valid_T_30=idxHit[1] ? idxPages_1:3'h0; 
  assign _io_resp_valid_T_31=idxHit[2] ? idxPages_2:3'h0; 
  assign _io_resp_valid_T_32=idxHit[3] ? idxPages_3:3'h0; 
  assign _io_resp_valid_T_33=idxHit[4] ? idxPages_4:3'h0; 
  assign _io_resp_valid_T_34=idxHit[5] ? idxPages_5:3'h0; 
  assign _io_resp_valid_T_35=idxHit[6] ? idxPages_6:3'h0; 
  assign _io_resp_valid_T_36=idxHit[7] ? idxPages_7:3'h0; 
  assign _io_resp_valid_T_37=idxHit[8] ? idxPages_8:3'h0; 
  assign _io_resp_valid_T_38=idxHit[9] ? idxPages_9:3'h0; 
  assign _io_resp_valid_T_39=idxHit[10] ? idxPages_10:3'h0; 
  assign _io_resp_valid_T_40=idxHit[11] ? idxPages_11:3'h0; 
  assign _io_resp_valid_T_41=idxHit[12] ? idxPages_12:3'h0; 
  assign _io_resp_valid_T_42=idxHit[13] ? idxPages_13:3'h0; 
  assign _io_resp_valid_T_43=idxHit[14] ? idxPages_14:3'h0; 
  assign _io_resp_valid_T_44=idxHit[15] ? idxPages_15:3'h0; 
  assign _io_resp_valid_T_45=idxHit[16] ? idxPages_16:3'h0; 
  assign _io_resp_valid_T_46=idxHit[17] ? idxPages_17:3'h0; 
  assign _io_resp_valid_T_47=idxHit[18] ? idxPages_18:3'h0; 
  assign _io_resp_valid_T_48=idxHit[19] ? idxPages_19:3'h0; 
  assign _io_resp_valid_T_49=idxHit[20] ? idxPages_20:3'h0; 
  assign _io_resp_valid_T_50=idxHit[21] ? idxPages_21:3'h0; 
  assign _io_resp_valid_T_51=idxHit[22] ? idxPages_22:3'h0; 
  assign _io_resp_valid_T_52=idxHit[23] ? idxPages_23:3'h0; 
  assign _io_resp_valid_T_53=idxHit[24] ? idxPages_24:3'h0; 
  assign _io_resp_valid_T_54=idxHit[25] ? idxPages_25:3'h0; 
  assign _io_resp_valid_T_55=idxHit[26] ? idxPages_26:3'h0; 
  assign _io_resp_valid_T_56=idxHit[27] ? idxPages_27:3'h0; 
  assign _io_resp_valid_T_57=_io_resp_valid_T_29|_io_resp_valid_T_30; 
  assign _io_resp_valid_T_58=_io_resp_valid_T_57|_io_resp_valid_T_31; 
  assign _io_resp_valid_T_59=_io_resp_valid_T_58|_io_resp_valid_T_32; 
  assign _io_resp_valid_T_60=_io_resp_valid_T_59|_io_resp_valid_T_33; 
  assign _io_resp_valid_T_61=_io_resp_valid_T_60|_io_resp_valid_T_34; 
  assign _io_resp_valid_T_62=_io_resp_valid_T_61|_io_resp_valid_T_35; 
  assign _io_resp_valid_T_63=_io_resp_valid_T_62|_io_resp_valid_T_36; 
  assign _io_resp_valid_T_64=_io_resp_valid_T_63|_io_resp_valid_T_37; 
  assign _io_resp_valid_T_65=_io_resp_valid_T_64|_io_resp_valid_T_38; 
  assign _io_resp_valid_T_66=_io_resp_valid_T_65|_io_resp_valid_T_39; 
  assign _io_resp_valid_T_67=_io_resp_valid_T_66|_io_resp_valid_T_40; 
  assign _io_resp_valid_T_68=_io_resp_valid_T_67|_io_resp_valid_T_41; 
  assign _io_resp_valid_T_69=_io_resp_valid_T_68|_io_resp_valid_T_42; 
  assign _io_resp_valid_T_70=_io_resp_valid_T_69|_io_resp_valid_T_43; 
  assign _io_resp_valid_T_71=_io_resp_valid_T_70|_io_resp_valid_T_44; 
  assign _io_resp_valid_T_72=_io_resp_valid_T_71|_io_resp_valid_T_45; 
  assign _io_resp_valid_T_73=_io_resp_valid_T_72|_io_resp_valid_T_46; 
  assign _io_resp_valid_T_74=_io_resp_valid_T_73|_io_resp_valid_T_47; 
  assign _io_resp_valid_T_75=_io_resp_valid_T_74|_io_resp_valid_T_48; 
  assign _io_resp_valid_T_76=_io_resp_valid_T_75|_io_resp_valid_T_49; 
  assign _io_resp_valid_T_77=_io_resp_valid_T_76|_io_resp_valid_T_50; 
  assign _io_resp_valid_T_78=_io_resp_valid_T_77|_io_resp_valid_T_51; 
  assign _io_resp_valid_T_79=_io_resp_valid_T_78|_io_resp_valid_T_52; 
  assign _io_resp_valid_T_80=_io_resp_valid_T_79|_io_resp_valid_T_53; 
  assign _io_resp_valid_T_81=_io_resp_valid_T_80|_io_resp_valid_T_54; 
  assign _io_resp_valid_T_82=_io_resp_valid_T_81|_io_resp_valid_T_55; 
  assign _io_resp_valid_T_83=_io_resp_valid_T_82|_io_resp_valid_T_56; 
  assign _io_resp_valid_T_84=_io_resp_valid_T>>_io_resp_valid_T_83; 
  assign _io_resp_bits_target_T_28=idxHit[0] ? tgtPages_0:3'h0; 
  assign _io_resp_bits_target_T_29=idxHit[1] ? tgtPages_1:3'h0; 
  assign _io_resp_bits_target_T_30=idxHit[2] ? tgtPages_2:3'h0; 
  assign _io_resp_bits_target_T_31=idxHit[3] ? tgtPages_3:3'h0; 
  assign _io_resp_bits_target_T_32=idxHit[4] ? tgtPages_4:3'h0; 
  assign _io_resp_bits_target_T_33=idxHit[5] ? tgtPages_5:3'h0; 
  assign _io_resp_bits_target_T_34=idxHit[6] ? tgtPages_6:3'h0; 
  assign _io_resp_bits_target_T_35=idxHit[7] ? tgtPages_7:3'h0; 
  assign _io_resp_bits_target_T_36=idxHit[8] ? tgtPages_8:3'h0; 
  assign _io_resp_bits_target_T_37=idxHit[9] ? tgtPages_9:3'h0; 
  assign _io_resp_bits_target_T_38=idxHit[10] ? tgtPages_10:3'h0; 
  assign _io_resp_bits_target_T_39=idxHit[11] ? tgtPages_11:3'h0; 
  assign _io_resp_bits_target_T_40=idxHit[12] ? tgtPages_12:3'h0; 
  assign _io_resp_bits_target_T_41=idxHit[13] ? tgtPages_13:3'h0; 
  assign _io_resp_bits_target_T_42=idxHit[14] ? tgtPages_14:3'h0; 
  assign _io_resp_bits_target_T_43=idxHit[15] ? tgtPages_15:3'h0; 
  assign _io_resp_bits_target_T_44=idxHit[16] ? tgtPages_16:3'h0; 
  assign _io_resp_bits_target_T_45=idxHit[17] ? tgtPages_17:3'h0; 
  assign _io_resp_bits_target_T_46=idxHit[18] ? tgtPages_18:3'h0; 
  assign _io_resp_bits_target_T_47=idxHit[19] ? tgtPages_19:3'h0; 
  assign _io_resp_bits_target_T_48=idxHit[20] ? tgtPages_20:3'h0; 
  assign _io_resp_bits_target_T_49=idxHit[21] ? tgtPages_21:3'h0; 
  assign _io_resp_bits_target_T_50=idxHit[22] ? tgtPages_22:3'h0; 
  assign _io_resp_bits_target_T_51=idxHit[23] ? tgtPages_23:3'h0; 
  assign _io_resp_bits_target_T_52=idxHit[24] ? tgtPages_24:3'h0; 
  assign _io_resp_bits_target_T_53=idxHit[25] ? tgtPages_25:3'h0; 
  assign _io_resp_bits_target_T_54=idxHit[26] ? tgtPages_26:3'h0; 
  assign _io_resp_bits_target_T_55=idxHit[27] ? tgtPages_27:3'h0; 
  assign _io_resp_bits_target_T_56=_io_resp_bits_target_T_28|_io_resp_bits_target_T_29; 
  assign _io_resp_bits_target_T_57=_io_resp_bits_target_T_56|_io_resp_bits_target_T_30; 
  assign _io_resp_bits_target_T_58=_io_resp_bits_target_T_57|_io_resp_bits_target_T_31; 
  assign _io_resp_bits_target_T_59=_io_resp_bits_target_T_58|_io_resp_bits_target_T_32; 
  assign _io_resp_bits_target_T_60=_io_resp_bits_target_T_59|_io_resp_bits_target_T_33; 
  assign _io_resp_bits_target_T_61=_io_resp_bits_target_T_60|_io_resp_bits_target_T_34; 
  assign _io_resp_bits_target_T_62=_io_resp_bits_target_T_61|_io_resp_bits_target_T_35; 
  assign _io_resp_bits_target_T_63=_io_resp_bits_target_T_62|_io_resp_bits_target_T_36; 
  assign _io_resp_bits_target_T_64=_io_resp_bits_target_T_63|_io_resp_bits_target_T_37; 
  assign _io_resp_bits_target_T_65=_io_resp_bits_target_T_64|_io_resp_bits_target_T_38; 
  assign _io_resp_bits_target_T_66=_io_resp_bits_target_T_65|_io_resp_bits_target_T_39; 
  assign _io_resp_bits_target_T_67=_io_resp_bits_target_T_66|_io_resp_bits_target_T_40; 
  assign _io_resp_bits_target_T_68=_io_resp_bits_target_T_67|_io_resp_bits_target_T_41; 
  assign _io_resp_bits_target_T_69=_io_resp_bits_target_T_68|_io_resp_bits_target_T_42; 
  assign _io_resp_bits_target_T_70=_io_resp_bits_target_T_69|_io_resp_bits_target_T_43; 
  assign _io_resp_bits_target_T_71=_io_resp_bits_target_T_70|_io_resp_bits_target_T_44; 
  assign _io_resp_bits_target_T_72=_io_resp_bits_target_T_71|_io_resp_bits_target_T_45; 
  assign _io_resp_bits_target_T_73=_io_resp_bits_target_T_72|_io_resp_bits_target_T_46; 
  assign _io_resp_bits_target_T_74=_io_resp_bits_target_T_73|_io_resp_bits_target_T_47; 
  assign _io_resp_bits_target_T_75=_io_resp_bits_target_T_74|_io_resp_bits_target_T_48; 
  assign _io_resp_bits_target_T_76=_io_resp_bits_target_T_75|_io_resp_bits_target_T_49; 
  assign _io_resp_bits_target_T_77=_io_resp_bits_target_T_76|_io_resp_bits_target_T_50; 
  assign _io_resp_bits_target_T_78=_io_resp_bits_target_T_77|_io_resp_bits_target_T_51; 
  assign _io_resp_bits_target_T_79=_io_resp_bits_target_T_78|_io_resp_bits_target_T_52; 
  assign _io_resp_bits_target_T_80=_io_resp_bits_target_T_79|_io_resp_bits_target_T_53; 
  assign _io_resp_bits_target_T_81=_io_resp_bits_target_T_80|_io_resp_bits_target_T_54; 
  assign _io_resp_bits_target_T_82=_io_resp_bits_target_T_81|_io_resp_bits_target_T_55; 
  assign _io_resp_bits_target_T_83=_io_resp_bits_target_T_82==3'h1; 
  assign _io_resp_bits_target_T_84=_io_resp_bits_target_T_83 ? pagesMasked_1:pagesMasked_0; 
  assign _io_resp_bits_target_T_85=_io_resp_bits_target_T_82==3'h2; 
  assign _io_resp_bits_target_T_86=_io_resp_bits_target_T_85 ? pagesMasked_2:_io_resp_bits_target_T_84; 
  assign _io_resp_bits_target_T_87=_io_resp_bits_target_T_82==3'h3; 
  assign _io_resp_bits_target_T_88=_io_resp_bits_target_T_87 ? pagesMasked_3:_io_resp_bits_target_T_86; 
  assign _io_resp_bits_target_T_89=_io_resp_bits_target_T_82==3'h4; 
  assign _io_resp_bits_target_T_90=_io_resp_bits_target_T_89 ? pagesMasked_4:_io_resp_bits_target_T_88; 
  assign _io_resp_bits_target_T_91=_io_resp_bits_target_T_82==3'h5; 
  assign _io_resp_bits_target_T_92=_io_resp_bits_target_T_91 ? pagesMasked_5:_io_resp_bits_target_T_90; 
  assign _io_resp_bits_target_T_93=_io_resp_bits_target_T_82==3'h6; 
  assign _io_resp_bits_target_T_94=_io_resp_bits_target_T_93 ? pagesMasked_4:_io_resp_bits_target_T_92; 
  assign _io_resp_bits_target_T_95=_io_resp_bits_target_T_82==3'h7; 
  assign io_resp_bits_target_hi=_io_resp_bits_target_T_95 ? pagesMasked_5:_io_resp_bits_target_T_94; 
  assign _io_resp_bits_target_T_124=idxHit[0] ? tgts_0:13'h0; 
  assign _io_resp_bits_target_T_125=idxHit[1] ? tgts_1:13'h0; 
  assign _io_resp_bits_target_T_126=idxHit[2] ? tgts_2:13'h0; 
  assign _io_resp_bits_target_T_127=idxHit[3] ? tgts_3:13'h0; 
  assign _io_resp_bits_target_T_128=idxHit[4] ? tgts_4:13'h0; 
  assign _io_resp_bits_target_T_129=idxHit[5] ? tgts_5:13'h0; 
  assign _io_resp_bits_target_T_130=idxHit[6] ? tgts_6:13'h0; 
  assign _io_resp_bits_target_T_131=idxHit[7] ? tgts_7:13'h0; 
  assign _io_resp_bits_target_T_132=idxHit[8] ? tgts_8:13'h0; 
  assign _io_resp_bits_target_T_133=idxHit[9] ? tgts_9:13'h0; 
  assign _io_resp_bits_target_T_134=idxHit[10] ? tgts_10:13'h0; 
  assign _io_resp_bits_target_T_135=idxHit[11] ? tgts_11:13'h0; 
  assign _io_resp_bits_target_T_136=idxHit[12] ? tgts_12:13'h0; 
  assign _io_resp_bits_target_T_137=idxHit[13] ? tgts_13:13'h0; 
  assign _io_resp_bits_target_T_138=idxHit[14] ? tgts_14:13'h0; 
  assign _io_resp_bits_target_T_139=idxHit[15] ? tgts_15:13'h0; 
  assign _io_resp_bits_target_T_140=idxHit[16] ? tgts_16:13'h0; 
  assign _io_resp_bits_target_T_141=idxHit[17] ? tgts_17:13'h0; 
  assign _io_resp_bits_target_T_142=idxHit[18] ? tgts_18:13'h0; 
  assign _io_resp_bits_target_T_143=idxHit[19] ? tgts_19:13'h0; 
  assign _io_resp_bits_target_T_144=idxHit[20] ? tgts_20:13'h0; 
  assign _io_resp_bits_target_T_145=idxHit[21] ? tgts_21:13'h0; 
  assign _io_resp_bits_target_T_146=idxHit[22] ? tgts_22:13'h0; 
  assign _io_resp_bits_target_T_147=idxHit[23] ? tgts_23:13'h0; 
  assign _io_resp_bits_target_T_148=idxHit[24] ? tgts_24:13'h0; 
  assign _io_resp_bits_target_T_149=idxHit[25] ? tgts_25:13'h0; 
  assign _io_resp_bits_target_T_150=idxHit[26] ? tgts_26:13'h0; 
  assign _io_resp_bits_target_T_151=idxHit[27] ? tgts_27:13'h0; 
  assign _io_resp_bits_target_T_152=_io_resp_bits_target_T_124|_io_resp_bits_target_T_125; 
  assign _io_resp_bits_target_T_153=_io_resp_bits_target_T_152|_io_resp_bits_target_T_126; 
  assign _io_resp_bits_target_T_154=_io_resp_bits_target_T_153|_io_resp_bits_target_T_127; 
  assign _io_resp_bits_target_T_155=_io_resp_bits_target_T_154|_io_resp_bits_target_T_128; 
  assign _io_resp_bits_target_T_156=_io_resp_bits_target_T_155|_io_resp_bits_target_T_129; 
  assign _io_resp_bits_target_T_157=_io_resp_bits_target_T_156|_io_resp_bits_target_T_130; 
  assign _io_resp_bits_target_T_158=_io_resp_bits_target_T_157|_io_resp_bits_target_T_131; 
  assign _io_resp_bits_target_T_159=_io_resp_bits_target_T_158|_io_resp_bits_target_T_132; 
  assign _io_resp_bits_target_T_160=_io_resp_bits_target_T_159|_io_resp_bits_target_T_133; 
  assign _io_resp_bits_target_T_161=_io_resp_bits_target_T_160|_io_resp_bits_target_T_134; 
  assign _io_resp_bits_target_T_162=_io_resp_bits_target_T_161|_io_resp_bits_target_T_135; 
  assign _io_resp_bits_target_T_163=_io_resp_bits_target_T_162|_io_resp_bits_target_T_136; 
  assign _io_resp_bits_target_T_164=_io_resp_bits_target_T_163|_io_resp_bits_target_T_137; 
  assign _io_resp_bits_target_T_165=_io_resp_bits_target_T_164|_io_resp_bits_target_T_138; 
  assign _io_resp_bits_target_T_166=_io_resp_bits_target_T_165|_io_resp_bits_target_T_139; 
  assign _io_resp_bits_target_T_167=_io_resp_bits_target_T_166|_io_resp_bits_target_T_140; 
  assign _io_resp_bits_target_T_168=_io_resp_bits_target_T_167|_io_resp_bits_target_T_141; 
  assign _io_resp_bits_target_T_169=_io_resp_bits_target_T_168|_io_resp_bits_target_T_142; 
  assign _io_resp_bits_target_T_170=_io_resp_bits_target_T_169|_io_resp_bits_target_T_143; 
  assign _io_resp_bits_target_T_171=_io_resp_bits_target_T_170|_io_resp_bits_target_T_144; 
  assign _io_resp_bits_target_T_172=_io_resp_bits_target_T_171|_io_resp_bits_target_T_145; 
  assign _io_resp_bits_target_T_173=_io_resp_bits_target_T_172|_io_resp_bits_target_T_146; 
  assign _io_resp_bits_target_T_174=_io_resp_bits_target_T_173|_io_resp_bits_target_T_147; 
  assign _io_resp_bits_target_T_175=_io_resp_bits_target_T_174|_io_resp_bits_target_T_148; 
  assign _io_resp_bits_target_T_176=_io_resp_bits_target_T_175|_io_resp_bits_target_T_149; 
  assign _io_resp_bits_target_T_177=_io_resp_bits_target_T_176|_io_resp_bits_target_T_150; 
  assign _io_resp_bits_target_T_178=_io_resp_bits_target_T_177|_io_resp_bits_target_T_151; 
  assign io_resp_bits_target_lo={_io_resp_bits_target_T_178,1'h0}; 
  assign _io_resp_bits_target_T_179={io_resp_bits_target_hi,io_resp_bits_target_lo}; 
  assign io_resp_bits_entry_hi=idxHit[27:16]; 
  assign io_resp_bits_entry_lo=idxHit[15:0]; 
  assign io_resp_bits_entry_hi_1=|io_resp_bits_entry_hi; 
  assign _GEN_436={4'b0,io_resp_bits_entry_hi}; 
  assign _io_resp_bits_entry_T=_GEN_436|io_resp_bits_entry_lo; 
  assign io_resp_bits_entry_hi_2=_io_resp_bits_entry_T[15:8]; 
  assign io_resp_bits_entry_lo_1=_io_resp_bits_entry_T[7:0]; 
  assign io_resp_bits_entry_hi_3=|io_resp_bits_entry_hi_2; 
  assign _io_resp_bits_entry_T_1=io_resp_bits_entry_hi_2|io_resp_bits_entry_lo_1; 
  assign io_resp_bits_entry_hi_4=_io_resp_bits_entry_T_1[7:4]; 
  assign io_resp_bits_entry_lo_2=_io_resp_bits_entry_T_1[3:0]; 
  assign io_resp_bits_entry_hi_5=|io_resp_bits_entry_hi_4; 
  assign _io_resp_bits_entry_T_2=io_resp_bits_entry_hi_4|io_resp_bits_entry_lo_2; 
  assign io_resp_bits_entry_hi_6=_io_resp_bits_entry_T_2[3:2]; 
  assign io_resp_bits_entry_lo_3=_io_resp_bits_entry_T_2[1:0]; 
  assign io_resp_bits_entry_hi_7=|io_resp_bits_entry_hi_6; 
  assign _io_resp_bits_entry_T_3=io_resp_bits_entry_hi_6|io_resp_bits_entry_lo_3; 
  assign io_resp_bits_entry_lo_4=_io_resp_bits_entry_T_3[1]; 
  assign io_resp_bits_entry_lo_7={io_resp_bits_entry_hi_3,io_resp_bits_entry_hi_5,io_resp_bits_entry_hi_7,io_resp_bits_entry_lo_4}; 
  assign _io_resp_bits_bridx_T_28=idxHit[0]&brIdx_0; 
  assign _io_resp_bits_bridx_T_29=idxHit[1]&brIdx_1; 
  assign _io_resp_bits_bridx_T_30=idxHit[2]&brIdx_2; 
  assign _io_resp_bits_bridx_T_31=idxHit[3]&brIdx_3; 
  assign _io_resp_bits_bridx_T_32=idxHit[4]&brIdx_4; 
  assign _io_resp_bits_bridx_T_33=idxHit[5]&brIdx_5; 
  assign _io_resp_bits_bridx_T_34=idxHit[6]&brIdx_6; 
  assign _io_resp_bits_bridx_T_35=idxHit[7]&brIdx_7; 
  assign _io_resp_bits_bridx_T_36=idxHit[8]&brIdx_8; 
  assign _io_resp_bits_bridx_T_37=idxHit[9]&brIdx_9; 
  assign _io_resp_bits_bridx_T_38=idxHit[10]&brIdx_10; 
  assign _io_resp_bits_bridx_T_39=idxHit[11]&brIdx_11; 
  assign _io_resp_bits_bridx_T_40=idxHit[12]&brIdx_12; 
  assign _io_resp_bits_bridx_T_41=idxHit[13]&brIdx_13; 
  assign _io_resp_bits_bridx_T_42=idxHit[14]&brIdx_14; 
  assign _io_resp_bits_bridx_T_43=idxHit[15]&brIdx_15; 
  assign _io_resp_bits_bridx_T_44=idxHit[16]&brIdx_16; 
  assign _io_resp_bits_bridx_T_45=idxHit[17]&brIdx_17; 
  assign _io_resp_bits_bridx_T_46=idxHit[18]&brIdx_18; 
  assign _io_resp_bits_bridx_T_47=idxHit[19]&brIdx_19; 
  assign _io_resp_bits_bridx_T_48=idxHit[20]&brIdx_20; 
  assign _io_resp_bits_bridx_T_49=idxHit[21]&brIdx_21; 
  assign _io_resp_bits_bridx_T_50=idxHit[22]&brIdx_22; 
  assign _io_resp_bits_bridx_T_51=idxHit[23]&brIdx_23; 
  assign _io_resp_bits_bridx_T_52=idxHit[24]&brIdx_24; 
  assign _io_resp_bits_bridx_T_53=idxHit[25]&brIdx_25; 
  assign _io_resp_bits_bridx_T_54=idxHit[26]&brIdx_26; 
  assign _io_resp_bits_bridx_T_55=idxHit[27]&brIdx_27; 
  assign _io_resp_bits_bridx_T_56=_io_resp_bits_bridx_T_28|_io_resp_bits_bridx_T_29; 
  assign _io_resp_bits_bridx_T_57=_io_resp_bits_bridx_T_56|_io_resp_bits_bridx_T_30; 
  assign _io_resp_bits_bridx_T_58=_io_resp_bits_bridx_T_57|_io_resp_bits_bridx_T_31; 
  assign _io_resp_bits_bridx_T_59=_io_resp_bits_bridx_T_58|_io_resp_bits_bridx_T_32; 
  assign _io_resp_bits_bridx_T_60=_io_resp_bits_bridx_T_59|_io_resp_bits_bridx_T_33; 
  assign _io_resp_bits_bridx_T_61=_io_resp_bits_bridx_T_60|_io_resp_bits_bridx_T_34; 
  assign _io_resp_bits_bridx_T_62=_io_resp_bits_bridx_T_61|_io_resp_bits_bridx_T_35; 
  assign _io_resp_bits_bridx_T_63=_io_resp_bits_bridx_T_62|_io_resp_bits_bridx_T_36; 
  assign _io_resp_bits_bridx_T_64=_io_resp_bits_bridx_T_63|_io_resp_bits_bridx_T_37; 
  assign _io_resp_bits_bridx_T_65=_io_resp_bits_bridx_T_64|_io_resp_bits_bridx_T_38; 
  assign _io_resp_bits_bridx_T_66=_io_resp_bits_bridx_T_65|_io_resp_bits_bridx_T_39; 
  assign _io_resp_bits_bridx_T_67=_io_resp_bits_bridx_T_66|_io_resp_bits_bridx_T_40; 
  assign _io_resp_bits_bridx_T_68=_io_resp_bits_bridx_T_67|_io_resp_bits_bridx_T_41; 
  assign _io_resp_bits_bridx_T_69=_io_resp_bits_bridx_T_68|_io_resp_bits_bridx_T_42; 
  assign _io_resp_bits_bridx_T_70=_io_resp_bits_bridx_T_69|_io_resp_bits_bridx_T_43; 
  assign _io_resp_bits_bridx_T_71=_io_resp_bits_bridx_T_70|_io_resp_bits_bridx_T_44; 
  assign _io_resp_bits_bridx_T_72=_io_resp_bits_bridx_T_71|_io_resp_bits_bridx_T_45; 
  assign _io_resp_bits_bridx_T_73=_io_resp_bits_bridx_T_72|_io_resp_bits_bridx_T_46; 
  assign _io_resp_bits_bridx_T_74=_io_resp_bits_bridx_T_73|_io_resp_bits_bridx_T_47; 
  assign _io_resp_bits_bridx_T_75=_io_resp_bits_bridx_T_74|_io_resp_bits_bridx_T_48; 
  assign _io_resp_bits_bridx_T_76=_io_resp_bits_bridx_T_75|_io_resp_bits_bridx_T_49; 
  assign _io_resp_bits_bridx_T_77=_io_resp_bits_bridx_T_76|_io_resp_bits_bridx_T_50; 
  assign _io_resp_bits_bridx_T_78=_io_resp_bits_bridx_T_77|_io_resp_bits_bridx_T_51; 
  assign _io_resp_bits_bridx_T_79=_io_resp_bits_bridx_T_78|_io_resp_bits_bridx_T_52; 
  assign _io_resp_bits_bridx_T_80=_io_resp_bits_bridx_T_79|_io_resp_bits_bridx_T_53; 
  assign _io_resp_bits_bridx_T_81=_io_resp_bits_bridx_T_80|_io_resp_bits_bridx_T_54; 
  assign leftOne=idxHit[0]; 
  assign leftOne_1=idxHit[1]; 
  assign rightOne=idxHit[2]; 
  assign rightOne_1=leftOne_1|rightOne; 
  assign rightTwo=leftOne_1&rightOne; 
  assign leftOne_2=leftOne|rightOne_1; 
  assign _T_29=leftOne&rightOne_1; 
  assign leftTwo=rightTwo|_T_29; 
  assign leftOne_3=idxHit[3]; 
  assign rightOne_2=idxHit[4]; 
  assign leftOne_4=leftOne_3|rightOne_2; 
  assign leftTwo_1=leftOne_3&rightOne_2; 
  assign leftOne_5=idxHit[5]; 
  assign rightOne_3=idxHit[6]; 
  assign rightOne_4=leftOne_5|rightOne_3; 
  assign rightTwo_1=leftOne_5&rightOne_3; 
  assign rightOne_5=leftOne_4|rightOne_4; 
  assign _T_41=leftTwo_1|rightTwo_1; 
  assign _T_42=leftOne_4&rightOne_4; 
  assign rightTwo_2=_T_41|_T_42; 
  assign leftOne_6=leftOne_2|rightOne_5; 
  assign _T_43=leftTwo|rightTwo_2; 
  assign _T_44=leftOne_2&rightOne_5; 
  assign leftTwo_2=_T_43|_T_44; 
  assign leftOne_7=idxHit[7]; 
  assign leftOne_8=idxHit[8]; 
  assign rightOne_6=idxHit[9]; 
  assign rightOne_7=leftOne_8|rightOne_6; 
  assign rightTwo_3=leftOne_8&rightOne_6; 
  assign leftOne_9=leftOne_7|rightOne_7; 
  assign _T_54=leftOne_7&rightOne_7; 
  assign leftTwo_3=rightTwo_3|_T_54; 
  assign leftOne_10=idxHit[10]; 
  assign rightOne_8=idxHit[11]; 
  assign leftOne_11=leftOne_10|rightOne_8; 
  assign leftTwo_4=leftOne_10&rightOne_8; 
  assign leftOne_12=idxHit[12]; 
  assign rightOne_9=idxHit[13]; 
  assign rightOne_10=leftOne_12|rightOne_9; 
  assign rightTwo_4=leftOne_12&rightOne_9; 
  assign rightOne_11=leftOne_11|rightOne_10; 
  assign _T_66=leftTwo_4|rightTwo_4; 
  assign _T_67=leftOne_11&rightOne_10; 
  assign rightTwo_5=_T_66|_T_67; 
  assign rightOne_12=leftOne_9|rightOne_11; 
  assign _T_68=leftTwo_3|rightTwo_5; 
  assign _T_69=leftOne_9&rightOne_11; 
  assign rightTwo_6=_T_68|_T_69; 
  assign leftOne_13=leftOne_6|rightOne_12; 
  assign _T_70=leftTwo_2|rightTwo_6; 
  assign _T_71=leftOne_6&rightOne_12; 
  assign leftTwo_5=_T_70|_T_71; 
  assign leftOne_14=idxHit[14]; 
  assign leftOne_15=idxHit[15]; 
  assign rightOne_13=idxHit[16]; 
  assign rightOne_14=leftOne_15|rightOne_13; 
  assign rightTwo_7=leftOne_15&rightOne_13; 
  assign leftOne_16=leftOne_14|rightOne_14; 
  assign _T_82=leftOne_14&rightOne_14; 
  assign leftTwo_6=rightTwo_7|_T_82; 
  assign leftOne_17=idxHit[17]; 
  assign rightOne_15=idxHit[18]; 
  assign leftOne_18=leftOne_17|rightOne_15; 
  assign leftTwo_7=leftOne_17&rightOne_15; 
  assign leftOne_19=idxHit[19]; 
  assign rightOne_16=idxHit[20]; 
  assign rightOne_17=leftOne_19|rightOne_16; 
  assign rightTwo_8=leftOne_19&rightOne_16; 
  assign rightOne_18=leftOne_18|rightOne_17; 
  assign _T_94=leftTwo_7|rightTwo_8; 
  assign _T_95=leftOne_18&rightOne_17; 
  assign rightTwo_9=_T_94|_T_95; 
  assign leftOne_20=leftOne_16|rightOne_18; 
  assign _T_96=leftTwo_6|rightTwo_9; 
  assign _T_97=leftOne_16&rightOne_18; 
  assign leftTwo_8=_T_96|_T_97; 
  assign leftOne_21=idxHit[21]; 
  assign leftOne_22=idxHit[22]; 
  assign rightOne_19=idxHit[23]; 
  assign rightOne_20=leftOne_22|rightOne_19; 
  assign rightTwo_10=leftOne_22&rightOne_19; 
  assign leftOne_23=leftOne_21|rightOne_20; 
  assign _T_107=leftOne_21&rightOne_20; 
  assign leftTwo_9=rightTwo_10|_T_107; 
  assign leftOne_24=idxHit[24]; 
  assign rightOne_21=idxHit[25]; 
  assign leftOne_25=leftOne_24|rightOne_21; 
  assign leftTwo_10=leftOne_24&rightOne_21; 
  assign leftOne_26=idxHit[26]; 
  assign rightOne_22=idxHit[27]; 
  assign rightOne_23=leftOne_26|rightOne_22; 
  assign rightTwo_11=leftOne_26&rightOne_22; 
  assign rightOne_24=leftOne_25|rightOne_23; 
  assign _T_119=leftTwo_10|rightTwo_11; 
  assign _T_120=leftOne_25&rightOne_23; 
  assign rightTwo_12=_T_119|_T_120; 
  assign rightOne_25=leftOne_23|rightOne_24; 
  assign _T_121=leftTwo_9|rightTwo_12; 
  assign _T_122=leftOne_23&rightOne_24; 
  assign rightTwo_13=_T_121|_T_122; 
  assign rightOne_26=leftOne_20|rightOne_25; 
  assign _T_123=leftTwo_8|rightTwo_13; 
  assign _T_124=leftOne_20&rightOne_25; 
  assign rightTwo_14=_T_123|_T_124; 
  assign _T_126=leftTwo_5|rightTwo_14; 
  assign _T_127=leftOne_13&rightOne_26; 
  assign _T_128=_T_126|_T_127; 
  assign _isValid_T_5=isValid&~idxHit; 
  assign _GEN_374=_T_128 ? {4'b0,_isValid_T_5}:_GEN_338; 
  assign _GEN_375=io_flush ? 32'h0:_GEN_374; 
  assign resetting=~reset_waddr[9]; 
  assign _reset_waddr_T_1=reset_waddr+10'h1; 
  assign waddr_hi_13=io_bht_update_bits_pc[38:2]; 
  assign _GEN_437={7'b0,waddr_hi_13[10:9]}; 
  assign _waddr_T_30=waddr_hi_13[8:0]^_GEN_437; 
  assign _waddr_T_31=8'hdd*io_bht_update_bits_prediction_history; 
  assign _waddr_T_33={_waddr_T_31[7:5],6'h0}; 
  assign _waddr_T_34=_waddr_T_30^_waddr_T_33; 
  assign _GEN_383=resetting ? reset_waddr:{1'b0,_waddr_T_34}; 
  assign _GEN_388=io_bht_update_bits_branch ? _GEN_383:reset_waddr; 
  assign waddr_1=io_bht_update_valid ? _GEN_388:reset_waddr; 
  assign _GEN_387=io_bht_update_bits_branch|resetting; 
  assign _GEN_384=~resetting&io_bht_update_bits_taken; 
  assign _GEN_389=io_bht_update_bits_branch&_GEN_384; 
  assign isBranch_lo_lo_lo_lo=cfiType_0==2'h0; 
  assign isBranch_lo_lo_lo_hi_lo=cfiType_1==2'h0; 
  assign isBranch_lo_lo_lo_hi_hi=cfiType_2==2'h0; 
  assign isBranch_lo_lo_hi_lo_lo=cfiType_3==2'h0; 
  assign isBranch_lo_lo_hi_lo_hi=cfiType_4==2'h0; 
  assign isBranch_lo_lo_hi_hi_lo=cfiType_5==2'h0; 
  assign isBranch_lo_lo_hi_hi_hi=cfiType_6==2'h0; 
  assign isBranch_lo_hi_lo_lo=cfiType_7==2'h0; 
  assign isBranch_lo_hi_lo_hi_lo=cfiType_8==2'h0; 
  assign isBranch_lo_hi_lo_hi_hi=cfiType_9==2'h0; 
  assign isBranch_lo_hi_hi_lo_lo=cfiType_10==2'h0; 
  assign isBranch_lo_hi_hi_lo_hi=cfiType_11==2'h0; 
  assign isBranch_lo_hi_hi_hi_lo=cfiType_12==2'h0; 
  assign isBranch_lo_hi_hi_hi_hi=cfiType_13==2'h0; 
  assign isBranch_hi_lo_lo_lo=cfiType_14==2'h0; 
  assign isBranch_hi_lo_lo_hi_lo=cfiType_15==2'h0; 
  assign isBranch_hi_lo_lo_hi_hi=cfiType_16==2'h0; 
  assign isBranch_hi_lo_hi_lo_lo=cfiType_17==2'h0; 
  assign isBranch_hi_lo_hi_lo_hi=cfiType_18==2'h0; 
  assign isBranch_hi_lo_hi_hi_lo=cfiType_19==2'h0; 
  assign isBranch_hi_lo_hi_hi_hi=cfiType_20==2'h0; 
  assign isBranch_hi_hi_lo_lo=cfiType_21==2'h0; 
  assign isBranch_hi_hi_lo_hi_lo=cfiType_22==2'h0; 
  assign isBranch_hi_hi_lo_hi_hi=cfiType_23==2'h0; 
  assign isBranch_hi_hi_hi_lo_lo=cfiType_24==2'h0; 
  assign isBranch_hi_hi_hi_lo_hi=cfiType_25==2'h0; 
  assign isBranch_hi_hi_hi_hi_lo=cfiType_26==2'h0; 
  assign isBranch_hi_hi_hi_hi_hi=cfiType_27==2'h0; 
  assign isBranch_lo_lo={isBranch_lo_lo_hi_hi_hi,isBranch_lo_lo_hi_hi_lo,isBranch_lo_lo_hi_lo_hi,isBranch_lo_lo_hi_lo_lo,isBranch_lo_lo_lo_hi_hi,isBranch_lo_lo_lo_hi_lo,isBranch_lo_lo_lo_lo}; 
  assign isBranch_lo={isBranch_lo_hi_hi_hi_hi,isBranch_lo_hi_hi_hi_lo,isBranch_lo_hi_hi_lo_hi,isBranch_lo_hi_hi_lo_lo,isBranch_lo_hi_lo_hi_hi,isBranch_lo_hi_lo_hi_lo,isBranch_lo_hi_lo_lo,isBranch_lo_lo}; 
  assign isBranch_hi_lo={isBranch_hi_lo_hi_hi_hi,isBranch_hi_lo_hi_hi_lo,isBranch_hi_lo_hi_lo_hi,isBranch_hi_lo_hi_lo_lo,isBranch_hi_lo_lo_hi_hi,isBranch_hi_lo_lo_hi_lo,isBranch_hi_lo_lo_lo}; 
  assign _isBranch_T={isBranch_hi_hi_hi_hi_hi,isBranch_hi_hi_hi_hi_lo,isBranch_hi_hi_hi_lo_hi,isBranch_hi_hi_hi_lo_lo,isBranch_hi_hi_lo_hi_hi,isBranch_hi_hi_lo_hi_lo,isBranch_hi_hi_lo_lo,isBranch_hi_lo,isBranch_lo}; 
  assign _isBranch_T_1=idxHit&_isBranch_T; 
  assign isBranch=|_isBranch_T_1; 
  assign res_res_value_hi=io_req_bits_addr[38:2]; 
  assign _GEN_438={7'b0,res_res_value_hi[10:9]}; 
  assign _res_res_value_T_3=res_res_value_hi[8:0]^_GEN_438; 
  assign _res_res_value_T_4=8'hdd*history; 
  assign _res_res_value_T_6={_res_res_value_T_4[7:5],6'h0}; 
  assign res_value=resetting ? 1'h0:table__res_res_value_MPORT_data; 
  assign history_lo=history[7:1]; 
  assign _history_T={io_bht_advance_bits_bht_value,history_lo}; 
  assign history_lo_1=io_bht_update_bits_prediction_history[7:1]; 
  assign _history_T_1={io_bht_update_bits_taken,history_lo_1}; 
  assign _T_134=~res_value&isBranch; 
  assign doPeek_lo_lo_lo_lo=cfiType_0==2'h3; 
  assign doPeek_lo_lo_lo_hi_lo=cfiType_1==2'h3; 
  assign doPeek_lo_lo_lo_hi_hi=cfiType_2==2'h3; 
  assign doPeek_lo_lo_hi_lo_lo=cfiType_3==2'h3; 
  assign doPeek_lo_lo_hi_lo_hi=cfiType_4==2'h3; 
  assign doPeek_lo_lo_hi_hi_lo=cfiType_5==2'h3; 
  assign doPeek_lo_lo_hi_hi_hi=cfiType_6==2'h3; 
  assign doPeek_lo_hi_lo_lo=cfiType_7==2'h3; 
  assign doPeek_lo_hi_lo_hi_lo=cfiType_8==2'h3; 
  assign doPeek_lo_hi_lo_hi_hi=cfiType_9==2'h3; 
  assign doPeek_lo_hi_hi_lo_lo=cfiType_10==2'h3; 
  assign doPeek_lo_hi_hi_lo_hi=cfiType_11==2'h3; 
  assign doPeek_lo_hi_hi_hi_lo=cfiType_12==2'h3; 
  assign doPeek_lo_hi_hi_hi_hi=cfiType_13==2'h3; 
  assign doPeek_hi_lo_lo_lo=cfiType_14==2'h3; 
  assign doPeek_hi_lo_lo_hi_lo=cfiType_15==2'h3; 
  assign doPeek_hi_lo_lo_hi_hi=cfiType_16==2'h3; 
  assign doPeek_hi_lo_hi_lo_lo=cfiType_17==2'h3; 
  assign doPeek_hi_lo_hi_lo_hi=cfiType_18==2'h3; 
  assign doPeek_hi_lo_hi_hi_lo=cfiType_19==2'h3; 
  assign doPeek_hi_lo_hi_hi_hi=cfiType_20==2'h3; 
  assign doPeek_hi_hi_lo_lo=cfiType_21==2'h3; 
  assign doPeek_hi_hi_lo_hi_lo=cfiType_22==2'h3; 
  assign doPeek_hi_hi_lo_hi_hi=cfiType_23==2'h3; 
  assign doPeek_hi_hi_hi_lo_lo=cfiType_24==2'h3; 
  assign doPeek_hi_hi_hi_lo_hi=cfiType_25==2'h3; 
  assign doPeek_hi_hi_hi_hi_lo=cfiType_26==2'h3; 
  assign doPeek_hi_hi_hi_hi_hi=cfiType_27==2'h3; 
  assign doPeek_lo_lo={doPeek_lo_lo_hi_hi_hi,doPeek_lo_lo_hi_hi_lo,doPeek_lo_lo_hi_lo_hi,doPeek_lo_lo_hi_lo_lo,doPeek_lo_lo_lo_hi_hi,doPeek_lo_lo_lo_hi_lo,doPeek_lo_lo_lo_lo}; 
  assign doPeek_lo={doPeek_lo_hi_hi_hi_hi,doPeek_lo_hi_hi_hi_lo,doPeek_lo_hi_hi_lo_hi,doPeek_lo_hi_hi_lo_lo,doPeek_lo_hi_lo_hi_hi,doPeek_lo_hi_lo_hi_lo,doPeek_lo_hi_lo_lo,doPeek_lo_lo}; 
  assign doPeek_hi_lo={doPeek_hi_lo_hi_hi_hi,doPeek_hi_lo_hi_hi_lo,doPeek_hi_lo_hi_lo_hi,doPeek_hi_lo_hi_lo_lo,doPeek_hi_lo_lo_hi_hi,doPeek_hi_lo_lo_hi_lo,doPeek_hi_lo_lo_lo}; 
  assign _doPeek_T={doPeek_hi_hi_hi_hi_hi,doPeek_hi_hi_hi_hi_lo,doPeek_hi_hi_hi_lo_hi,doPeek_hi_hi_hi_lo_lo,doPeek_hi_hi_lo_hi_hi,doPeek_hi_hi_lo_hi_lo,doPeek_hi_hi_lo_lo,doPeek_hi_lo,doPeek_lo}; 
  assign _doPeek_T_1=idxHit&_doPeek_T; 
  assign doPeek=|_doPeek_T_1; 
  assign _io_ras_head_valid_T=count==3'h0; 
  assign _GEN_397=3'h1==pos ? stack_1:stack_0; 
  assign _GEN_398=3'h2==pos ? stack_2:_GEN_397; 
  assign _GEN_399=3'h3==pos ? stack_3:_GEN_398; 
  assign _GEN_400=3'h4==pos ? stack_4:_GEN_399; 
  assign _GEN_401=3'h5==pos ? stack_5:_GEN_400; 
  assign _T_137=~_io_ras_head_valid_T&doPeek; 
  assign _T_138=io_ras_update_bits_cfiType==2'h2; 
  assign _T_139=count<3'h6; 
  assign _count_T_1=count+3'h1; 
  assign _nextPos_T=pos<3'h5; 
  assign _nextPos_T_3=pos+3'h1; 
  assign nextPos=_nextPos_T ? _nextPos_T_3:3'h0; 
  assign _T_140=io_ras_update_bits_cfiType==2'h3; 
  assign _count_T_3=count-3'h1; 
  assign _pos_T=pos>3'h0; 
  assign _pos_T_3=pos-3'h1; 
  assign io_resp_valid=_io_resp_valid_T_84[0]; 
  assign io_resp_bits_taken=_T_134 ? 1'h0:1'h1; 
  assign io_resp_bits_bridx=_io_resp_bits_bridx_T_81|_io_resp_bits_bridx_T_55; 
  assign io_resp_bits_target=_T_137 ? _GEN_401:_io_resp_bits_target_T_179; 
  assign io_resp_bits_entry={io_resp_bits_entry_hi_1,io_resp_bits_entry_lo_7}; 
  assign io_resp_bits_bht_history=history; 
  assign io_resp_bits_bht_value=resetting ? 1'h0:table__res_res_value_MPORT_data; 
  assign io_ras_head_valid=~_io_ras_head_valid_T; 
  assign io_ras_head_bits=3'h5==pos ? stack_5:_GEN_400; 
  assign BTB_cov_read_addr=BTB_state; 
  assign BTB_cov_read_data=BTB_cov[BTB_cov_read_addr]; 
  assign BTB_cov_write_data=1'h1; 
  assign BTB_cov_write_addr=BTB_state; 
  assign BTB_cov_write_mask=1'h1; 
  assign BTB_cov_write_en=1'h1; 
  assign mux_cond_0=idxHit[19]; 
  assign mux_cond_1=idxHit[20]; 
  assign mux_cond_2=idxHit[27]; 
  assign mux_cond_3=idxHit[5]; 
  assign mux_cond_4=idxHit[6]; 
  assign mux_cond_5=idxHit[15]; 
  assign mux_cond_6=idxHit[23]; 
  assign mux_cond_7=idxHit[1]; 
  assign mux_cond_8=idxHit[10]; 
  assign mux_cond_9=idxHit[26]; 
  assign mux_cond_10=idxHit[13]; 
  assign mux_cond_11=idxHit[24]; 
  assign mux_cond_12=idxHit[2]; 
  assign mux_cond_13=idxHit[12]; 
  assign mux_cond_14=idxHit[17]; 
  assign mux_cond_15=idxHit[0]; 
  assign mux_cond_16=idxHit[4]; 
  assign mux_cond_17=idxHit[22]; 
  assign mux_cond_18=idxHit[3]; 
  assign mux_cond_19=idxHit[18]; 
  assign mux_cond_20=idxHit[11]; 
  assign mux_cond_21=idxHit[8]; 
  assign mux_cond_22=idxHit[21]; 
  assign mux_cond_23=idxHit[25]; 
  assign mux_cond_24=_T_128; 
  assign mux_cond_25=idxHit[7]; 
  assign mux_cond_26=idxHit[14]; 
  assign mux_cond_27=idxHit[16]; 
  assign mux_cond_28=idxHit[9]; 
  assign nextPageRepl_shl={nextPageRepl,7'h0}; 
  assign nextPageRepl_pad={10'h0,nextPageRepl_shl}; 
  assign r_respPipe_bits_taken_shl={r_respPipe_bits_taken,3'h0}; 
  assign r_respPipe_bits_taken_pad={16'h0,r_respPipe_bits_taken_shl}; 
  assign r_btb_updatePipe_valid_shl={r_btb_updatePipe_valid,16'h0}; 
  assign r_btb_updatePipe_valid_pad={3'h0,r_btb_updatePipe_valid_shl}; 
  assign count_shl={count,12'h0}; 
  assign count_pad={5'h0,count_shl}; 
  assign r_respPipe_valid_shl={r_respPipe_valid,13'h0}; 
  assign r_respPipe_valid_pad={6'h0,r_respPipe_valid_shl}; 
  assign pos_shl={pos,1'h0}; 
  assign pos_pad={16'h0,pos_shl}; 
  assign pageValid_shl={pageValid,8'h0}; 
  assign pageValid_pad={6'h0,pageValid_shl}; 
  assign r_btb_updatePipe_bits_isValid_shl={r_btb_updatePipe_bits_isValid,17'h0}; 
  assign r_btb_updatePipe_bits_isValid_pad={2'h0,r_btb_updatePipe_bits_isValid_shl}; 
  assign mux_cond_0_shl={mux_cond_0,14'h0}; 
  assign mux_cond_0_pad={5'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,17'h0}; 
  assign mux_cond_1_pad={2'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl={mux_cond_2,3'h0}; 
  assign mux_cond_2_pad={16'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,17'h0}; 
  assign mux_cond_3_pad={2'h0,mux_cond_3_shl}; 
  assign mux_cond_4_shl={mux_cond_4,13'h0}; 
  assign mux_cond_4_pad={6'h0,mux_cond_4_shl}; 
  assign mux_cond_5_shl={mux_cond_5,3'h0}; 
  assign mux_cond_5_pad={16'h0,mux_cond_5_shl}; 
  assign mux_cond_6_shl={mux_cond_6,1'h0}; 
  assign mux_cond_6_pad={18'h0,mux_cond_6_shl}; 
  assign mux_cond_7_shl={mux_cond_7,13'h0}; 
  assign mux_cond_7_pad={6'h0,mux_cond_7_shl}; 
  assign mux_cond_8_shl={mux_cond_8,16'h0}; 
  assign mux_cond_8_pad={3'h0,mux_cond_8_shl}; 
  assign mux_cond_9_shl={mux_cond_9,3'h0}; 
  assign mux_cond_9_pad={16'h0,mux_cond_9_shl}; 
  assign mux_cond_10_shl={mux_cond_10,9'h0}; 
  assign mux_cond_10_pad={10'h0,mux_cond_10_shl}; 
  assign mux_cond_11_shl={mux_cond_11,3'h0}; 
  assign mux_cond_11_pad={16'h0,mux_cond_11_shl}; 
  assign mux_cond_12_shl={mux_cond_12,17'h0}; 
  assign mux_cond_12_pad={2'h0,mux_cond_12_shl}; 
  assign mux_cond_13_shl={mux_cond_13,8'h0}; 
  assign mux_cond_13_pad={11'h0,mux_cond_13_shl}; 
  assign mux_cond_14_shl={mux_cond_14,4'h0}; 
  assign mux_cond_14_pad={15'h0,mux_cond_14_shl}; 
  assign mux_cond_15_shl={mux_cond_15,11'h0}; 
  assign mux_cond_15_pad={8'h0,mux_cond_15_shl}; 
  assign mux_cond_16_shl={mux_cond_16,12'h0}; 
  assign mux_cond_16_pad={7'h0,mux_cond_16_shl}; 
  assign mux_cond_17_shl={mux_cond_17,5'h0}; 
  assign mux_cond_17_pad={14'h0,mux_cond_17_shl}; 
  assign mux_cond_18_shl=mux_cond_18; 
  assign mux_cond_18_pad={19'h0,mux_cond_18_shl}; 
  assign mux_cond_19_shl={mux_cond_19,1'h0}; 
  assign mux_cond_19_pad={18'h0,mux_cond_19_shl}; 
  assign mux_cond_20_shl={mux_cond_20,2'h0}; 
  assign mux_cond_20_pad={17'h0,mux_cond_20_shl}; 
  assign mux_cond_21_shl={mux_cond_21,5'h0}; 
  assign mux_cond_21_pad={14'h0,mux_cond_21_shl}; 
  assign mux_cond_22_shl={mux_cond_22,16'h0}; 
  assign mux_cond_22_pad={3'h0,mux_cond_22_shl}; 
  assign mux_cond_23_shl={mux_cond_23,13'h0}; 
  assign mux_cond_23_pad={6'h0,mux_cond_23_shl}; 
  assign mux_cond_24_shl={mux_cond_24,19'h0}; 
  assign mux_cond_24_pad=mux_cond_24_shl; 
  assign mux_cond_25_shl={mux_cond_25,14'h0}; 
  assign mux_cond_25_pad={5'h0,mux_cond_25_shl}; 
  assign mux_cond_26_shl={mux_cond_26,8'h0}; 
  assign mux_cond_26_pad={11'h0,mux_cond_26_shl}; 
  assign mux_cond_27_shl={mux_cond_27,18'h0}; 
  assign mux_cond_27_pad={1'h0,mux_cond_27_shl}; 
  assign mux_cond_28_shl={mux_cond_28,5'h0}; 
  assign mux_cond_28_pad={14'h0,mux_cond_28_shl}; 
  assign cfiType_17_shl={cfiType_17,11'h0}; 
  assign cfiType_17_pad={7'h0,cfiType_17_shl}; 
  assign cfiType_22_shl={cfiType_22,11'h0}; 
  assign cfiType_22_pad={7'h0,cfiType_22_shl}; 
  assign cfiType_21_shl={cfiType_21,11'h0}; 
  assign cfiType_21_pad={7'h0,cfiType_21_shl}; 
  assign tgtPages_4_shl={tgtPages_4,15'h0}; 
  assign tgtPages_4_pad={2'h0,tgtPages_4_shl}; 
  assign tgtPages_6_shl={tgtPages_6,15'h0}; 
  assign tgtPages_6_pad={2'h0,tgtPages_6_shl}; 
  assign tgtPages_11_shl={tgtPages_11,15'h0}; 
  assign tgtPages_11_pad={2'h0,tgtPages_11_shl}; 
  assign tgtPages_7_shl={tgtPages_7,15'h0}; 
  assign tgtPages_7_pad={2'h0,tgtPages_7_shl}; 
  assign tgtPages_20_shl={tgtPages_20,15'h0}; 
  assign tgtPages_20_pad={2'h0,tgtPages_20_shl}; 
  assign cfiType_3_shl={cfiType_3,11'h0}; 
  assign cfiType_3_pad={7'h0,cfiType_3_shl}; 
  assign tgtPages_16_shl={tgtPages_16,15'h0}; 
  assign tgtPages_16_pad={2'h0,tgtPages_16_shl}; 
  assign cfiType_24_shl={cfiType_24,11'h0}; 
  assign cfiType_24_pad={7'h0,cfiType_24_shl}; 
  assign tgtPages_17_shl={tgtPages_17,15'h0}; 
  assign tgtPages_17_pad={2'h0,tgtPages_17_shl}; 
  assign cfiType_6_shl={cfiType_6,11'h0}; 
  assign cfiType_6_pad={7'h0,cfiType_6_shl}; 
  assign tgtPages_9_shl={tgtPages_9,15'h0}; 
  assign tgtPages_9_pad={2'h0,tgtPages_9_shl}; 
  assign tgtPages_2_shl={tgtPages_2,15'h0}; 
  assign tgtPages_2_pad={2'h0,tgtPages_2_shl}; 
  assign cfiType_10_shl={cfiType_10,11'h0}; 
  assign cfiType_10_pad={7'h0,cfiType_10_shl}; 
  assign tgtPages_18_shl={tgtPages_18,15'h0}; 
  assign tgtPages_18_pad={2'h0,tgtPages_18_shl}; 
  assign tgtPages_0_shl={tgtPages_0,15'h0}; 
  assign tgtPages_0_pad={2'h0,tgtPages_0_shl}; 
  assign tgtPages_25_shl={tgtPages_25,15'h0}; 
  assign tgtPages_25_pad={2'h0,tgtPages_25_shl}; 
  assign tgtPages_22_shl={tgtPages_22,15'h0}; 
  assign tgtPages_22_pad={2'h0,tgtPages_22_shl}; 
  assign cfiType_5_shl={cfiType_5,11'h0}; 
  assign cfiType_5_pad={7'h0,cfiType_5_shl}; 
  assign cfiType_12_shl={cfiType_12,11'h0}; 
  assign cfiType_12_pad={7'h0,cfiType_12_shl}; 
  assign cfiType_18_shl={cfiType_18,11'h0}; 
  assign cfiType_18_pad={7'h0,cfiType_18_shl}; 
  assign tgtPages_24_shl={tgtPages_24,15'h0}; 
  assign tgtPages_24_pad={2'h0,tgtPages_24_shl}; 
  assign tgtPages_26_shl={tgtPages_26,15'h0}; 
  assign tgtPages_26_pad={2'h0,tgtPages_26_shl}; 
  assign tgtPages_1_shl={tgtPages_1,15'h0}; 
  assign tgtPages_1_pad={2'h0,tgtPages_1_shl}; 
  assign tgtPages_10_shl={tgtPages_10,15'h0}; 
  assign tgtPages_10_pad={2'h0,tgtPages_10_shl}; 
  assign cfiType_25_shl={cfiType_25,11'h0}; 
  assign cfiType_25_pad={7'h0,cfiType_25_shl}; 
  assign cfiType_16_shl={cfiType_16,11'h0}; 
  assign cfiType_16_pad={7'h0,cfiType_16_shl}; 
  assign tgtPages_13_shl={tgtPages_13,15'h0}; 
  assign tgtPages_13_pad={2'h0,tgtPages_13_shl}; 
  assign cfiType_19_shl={cfiType_19,11'h0}; 
  assign cfiType_19_pad={7'h0,cfiType_19_shl}; 
  assign cfiType_2_shl={cfiType_2,11'h0}; 
  assign cfiType_2_pad={7'h0,cfiType_2_shl}; 
  assign cfiType_20_shl={cfiType_20,11'h0}; 
  assign cfiType_20_pad={7'h0,cfiType_20_shl}; 
  assign tgtPages_15_shl={tgtPages_15,15'h0}; 
  assign tgtPages_15_pad={2'h0,tgtPages_15_shl}; 
  assign tgtPages_8_shl={tgtPages_8,15'h0}; 
  assign tgtPages_8_pad={2'h0,tgtPages_8_shl}; 
  assign tgtPages_5_shl={tgtPages_5,15'h0}; 
  assign tgtPages_5_pad={2'h0,tgtPages_5_shl}; 
  assign cfiType_0_shl={cfiType_0,11'h0}; 
  assign cfiType_0_pad={7'h0,cfiType_0_shl}; 
  assign tgtPages_3_shl={tgtPages_3,15'h0}; 
  assign tgtPages_3_pad={2'h0,tgtPages_3_shl}; 
  assign tgtPages_27_shl={tgtPages_27,15'h0}; 
  assign tgtPages_27_pad={2'h0,tgtPages_27_shl}; 
  assign cfiType_27_shl={cfiType_27,11'h0}; 
  assign cfiType_27_pad={7'h0,cfiType_27_shl}; 
  assign tgtPages_14_shl={tgtPages_14,15'h0}; 
  assign tgtPages_14_pad={2'h0,tgtPages_14_shl}; 
  assign cfiType_13_shl={cfiType_13,11'h0}; 
  assign cfiType_13_pad={7'h0,cfiType_13_shl}; 
  assign cfiType_23_shl={cfiType_23,11'h0}; 
  assign cfiType_23_pad={7'h0,cfiType_23_shl}; 
  assign cfiType_4_shl={cfiType_4,11'h0}; 
  assign cfiType_4_pad={7'h0,cfiType_4_shl}; 
  assign cfiType_1_shl={cfiType_1,11'h0}; 
  assign cfiType_1_pad={7'h0,cfiType_1_shl}; 
  assign tgtPages_21_shl={tgtPages_21,15'h0}; 
  assign tgtPages_21_pad={2'h0,tgtPages_21_shl}; 
  assign cfiType_8_shl={cfiType_8,11'h0}; 
  assign cfiType_8_pad={7'h0,cfiType_8_shl}; 
  assign tgtPages_23_shl={tgtPages_23,15'h0}; 
  assign tgtPages_23_pad={2'h0,tgtPages_23_shl}; 
  assign tgtPages_19_shl={tgtPages_19,15'h0}; 
  assign tgtPages_19_pad={2'h0,tgtPages_19_shl}; 
  assign cfiType_11_shl={cfiType_11,11'h0}; 
  assign cfiType_11_pad={7'h0,cfiType_11_shl}; 
  assign tgtPages_12_shl={tgtPages_12,15'h0}; 
  assign tgtPages_12_pad={2'h0,tgtPages_12_shl}; 
  assign cfiType_9_shl={cfiType_9,11'h0}; 
  assign cfiType_9_pad={7'h0,cfiType_9_shl}; 
  assign cfiType_14_shl={cfiType_14,11'h0}; 
  assign cfiType_14_pad={7'h0,cfiType_14_shl}; 
  assign cfiType_7_shl={cfiType_7,11'h0}; 
  assign cfiType_7_pad={7'h0,cfiType_7_shl}; 
  assign cfiType_26_shl={cfiType_26,11'h0}; 
  assign cfiType_26_pad={7'h0,cfiType_26_shl}; 
  assign cfiType_15_shl={cfiType_15,11'h0}; 
  assign cfiType_15_pad={7'h0,cfiType_15_shl}; 
  assign BTB_xor31=nextPageRepl_pad^r_respPipe_bits_taken_pad; 
  assign BTB_xor66=count_pad^r_respPipe_valid_pad; 
  assign BTB_xor32=r_btb_updatePipe_valid_pad^BTB_xor66; 
  assign BTB_xor15=BTB_xor31^BTB_xor32; 
  assign BTB_xor68=pageValid_pad^r_btb_updatePipe_bits_isValid_pad; 
  assign BTB_xor33=pos_pad^BTB_xor68; 
  assign BTB_xor70=mux_cond_1_pad^mux_cond_2_pad; 
  assign BTB_xor34=mux_cond_0_pad^BTB_xor70; 
  assign BTB_xor16=BTB_xor33^BTB_xor34; 
  assign BTB_xor7=BTB_xor15^BTB_xor16; 
  assign BTB_xor72=mux_cond_4_pad^mux_cond_5_pad; 
  assign BTB_xor35=mux_cond_3_pad^BTB_xor72; 
  assign BTB_xor74=mux_cond_7_pad^mux_cond_8_pad; 
  assign BTB_xor36=mux_cond_6_pad^BTB_xor74; 
  assign BTB_xor17=BTB_xor35^BTB_xor36; 
  assign BTB_xor76=mux_cond_10_pad^mux_cond_11_pad; 
  assign BTB_xor37=mux_cond_9_pad^BTB_xor76; 
  assign BTB_xor78=mux_cond_13_pad^mux_cond_14_pad; 
  assign BTB_xor38=mux_cond_12_pad^BTB_xor78; 
  assign BTB_xor18=BTB_xor37^BTB_xor38; 
  assign BTB_xor8=BTB_xor17^BTB_xor18; 
  assign BTB_xor3=BTB_xor7^BTB_xor8; 
  assign BTB_xor39=mux_cond_15_pad^mux_cond_16_pad; 
  assign BTB_xor82=mux_cond_18_pad^mux_cond_19_pad; 
  assign BTB_xor40=mux_cond_17_pad^BTB_xor82; 
  assign BTB_xor19=BTB_xor39^BTB_xor40; 
  assign BTB_xor84=mux_cond_21_pad^mux_cond_22_pad; 
  assign BTB_xor41=mux_cond_20_pad^BTB_xor84; 
  assign BTB_xor86=mux_cond_24_pad^mux_cond_25_pad; 
  assign BTB_xor42=mux_cond_23_pad^BTB_xor86; 
  assign BTB_xor20=BTB_xor41^BTB_xor42; 
  assign BTB_xor9=BTB_xor19^BTB_xor20; 
  assign BTB_xor88=mux_cond_27_pad^mux_cond_28_pad; 
  assign BTB_xor43=mux_cond_26_pad^BTB_xor88; 
  assign BTB_xor90=cfiType_22_pad^cfiType_21_pad; 
  assign BTB_xor44=cfiType_17_pad^BTB_xor90; 
  assign BTB_xor21=BTB_xor43^BTB_xor44; 
  assign BTB_xor92=tgtPages_6_pad^tgtPages_11_pad; 
  assign BTB_xor45=tgtPages_4_pad^BTB_xor92; 
  assign BTB_xor94=tgtPages_20_pad^cfiType_3_pad; 
  assign BTB_xor46=tgtPages_7_pad^BTB_xor94; 
  assign BTB_xor22=BTB_xor45^BTB_xor46; 
  assign BTB_xor10=BTB_xor21^BTB_xor22; 
  assign BTB_xor4=BTB_xor9^BTB_xor10; 
  assign BTB_xor1=BTB_xor3^BTB_xor4; 
  assign BTB_xor47=tgtPages_16_pad^cfiType_24_pad; 
  assign BTB_xor98=cfiType_6_pad^tgtPages_9_pad; 
  assign BTB_xor48=tgtPages_17_pad^BTB_xor98; 
  assign BTB_xor23=BTB_xor47^BTB_xor48; 
  assign BTB_xor100=cfiType_10_pad^tgtPages_18_pad; 
  assign BTB_xor49=tgtPages_2_pad^BTB_xor100; 
  assign BTB_xor102=tgtPages_25_pad^tgtPages_22_pad; 
  assign BTB_xor50=tgtPages_0_pad^BTB_xor102; 
  assign BTB_xor24=BTB_xor49^BTB_xor50; 
  assign BTB_xor11=BTB_xor23^BTB_xor24; 
  assign BTB_xor104=cfiType_12_pad^cfiType_18_pad; 
  assign BTB_xor51=cfiType_5_pad^BTB_xor104; 
  assign BTB_xor106=tgtPages_26_pad^tgtPages_1_pad; 
  assign BTB_xor52=tgtPages_24_pad^BTB_xor106; 
  assign BTB_xor25=BTB_xor51^BTB_xor52; 
  assign BTB_xor108=cfiType_25_pad^cfiType_16_pad; 
  assign BTB_xor53=tgtPages_10_pad^BTB_xor108; 
  assign BTB_xor110=cfiType_19_pad^cfiType_2_pad; 
  assign BTB_xor54=tgtPages_13_pad^BTB_xor110; 
  assign BTB_xor26=BTB_xor53^BTB_xor54; 
  assign BTB_xor12=BTB_xor25^BTB_xor26; 
  assign BTB_xor5=BTB_xor11^BTB_xor12; 
  assign BTB_xor112=tgtPages_15_pad^tgtPages_8_pad; 
  assign BTB_xor55=cfiType_20_pad^BTB_xor112; 
  assign BTB_xor114=cfiType_0_pad^tgtPages_3_pad; 
  assign BTB_xor56=tgtPages_5_pad^BTB_xor114; 
  assign BTB_xor27=BTB_xor55^BTB_xor56; 
  assign BTB_xor116=cfiType_27_pad^tgtPages_14_pad; 
  assign BTB_xor57=tgtPages_27_pad^BTB_xor116; 
  assign BTB_xor118=cfiType_23_pad^cfiType_4_pad; 
  assign BTB_xor58=cfiType_13_pad^BTB_xor118; 
  assign BTB_xor28=BTB_xor57^BTB_xor58; 
  assign BTB_xor13=BTB_xor27^BTB_xor28; 
  assign BTB_xor120=tgtPages_21_pad^cfiType_8_pad; 
  assign BTB_xor59=cfiType_1_pad^BTB_xor120; 
  assign BTB_xor122=tgtPages_19_pad^cfiType_11_pad; 
  assign BTB_xor60=tgtPages_23_pad^BTB_xor122; 
  assign BTB_xor29=BTB_xor59^BTB_xor60; 
  assign BTB_xor124=cfiType_9_pad^cfiType_14_pad; 
  assign BTB_xor61=tgtPages_12_pad^BTB_xor124; 
  assign BTB_xor126=cfiType_26_pad^cfiType_15_pad; 
  assign BTB_xor62=cfiType_7_pad^BTB_xor126; 
  assign BTB_xor30=BTB_xor61^BTB_xor62; 
  assign BTB_xor14=BTB_xor29^BTB_xor30; 
  assign BTB_xor6=BTB_xor13^BTB_xor14; 
  assign BTB_xor2=BTB_xor5^BTB_xor6; 
  assign BTB_xor0=BTB_xor1^BTB_xor2; 
  assign io_covSum=BTB_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (table__MPORT_en&table__MPORT_mask)
            begin 
              table_ [table__MPORT_addr]<=table__MPORT_data;
            end 
         if (metaReset)
            begin 
              idxs_0 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h0==waddr)
                    begin 
                      idxs_0 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_1 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1==waddr)
                    begin 
                      idxs_1 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_2 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h2==waddr)
                    begin 
                      idxs_2 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_3 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h3==waddr)
                    begin 
                      idxs_3 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_4 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h4==waddr)
                    begin 
                      idxs_4 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_5 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h5==waddr)
                    begin 
                      idxs_5 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_6 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h6==waddr)
                    begin 
                      idxs_6 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_7 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h7==waddr)
                    begin 
                      idxs_7 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_8 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h8==waddr)
                    begin 
                      idxs_8 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_9 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h9==waddr)
                    begin 
                      idxs_9 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_10 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'ha==waddr)
                    begin 
                      idxs_10 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_11 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hb==waddr)
                    begin 
                      idxs_11 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_12 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hc==waddr)
                    begin 
                      idxs_12 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_13 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hd==waddr)
                    begin 
                      idxs_13 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_14 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'he==waddr)
                    begin 
                      idxs_14 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_15 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hf==waddr)
                    begin 
                      idxs_15 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_16 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h10==waddr)
                    begin 
                      idxs_16 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_17 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h11==waddr)
                    begin 
                      idxs_17 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_18 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h12==waddr)
                    begin 
                      idxs_18 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_19 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h13==waddr)
                    begin 
                      idxs_19 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_20 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h14==waddr)
                    begin 
                      idxs_20 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_21 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h15==waddr)
                    begin 
                      idxs_21 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_22 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h16==waddr)
                    begin 
                      idxs_22 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_23 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h17==waddr)
                    begin 
                      idxs_23 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_24 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h18==waddr)
                    begin 
                      idxs_24 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_25 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h19==waddr)
                    begin 
                      idxs_25 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_26 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1a==waddr)
                    begin 
                      idxs_26 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxs_27 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1b==waddr)
                    begin 
                      idxs_27 <=r_btb_updatePipe_bits_pc[13:1];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_0 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h0==waddr)
                    begin 
                      idxPages_0 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_1 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1==waddr)
                    begin 
                      idxPages_1 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_2 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h2==waddr)
                    begin 
                      idxPages_2 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_3 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h3==waddr)
                    begin 
                      idxPages_3 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_4 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h4==waddr)
                    begin 
                      idxPages_4 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_5 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h5==waddr)
                    begin 
                      idxPages_5 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_6 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h6==waddr)
                    begin 
                      idxPages_6 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_7 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h7==waddr)
                    begin 
                      idxPages_7 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_8 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h8==waddr)
                    begin 
                      idxPages_8 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_9 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h9==waddr)
                    begin 
                      idxPages_9 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_10 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'ha==waddr)
                    begin 
                      idxPages_10 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_11 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hb==waddr)
                    begin 
                      idxPages_11 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_12 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hc==waddr)
                    begin 
                      idxPages_12 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_13 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hd==waddr)
                    begin 
                      idxPages_13 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_14 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'he==waddr)
                    begin 
                      idxPages_14 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_15 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hf==waddr)
                    begin 
                      idxPages_15 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_16 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h10==waddr)
                    begin 
                      idxPages_16 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_17 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h11==waddr)
                    begin 
                      idxPages_17 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_18 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h12==waddr)
                    begin 
                      idxPages_18 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_19 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h13==waddr)
                    begin 
                      idxPages_19 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_20 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h14==waddr)
                    begin 
                      idxPages_20 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_21 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h15==waddr)
                    begin 
                      idxPages_21 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_22 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h16==waddr)
                    begin 
                      idxPages_22 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_23 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h17==waddr)
                    begin 
                      idxPages_23 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_24 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h18==waddr)
                    begin 
                      idxPages_24 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_25 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h19==waddr)
                    begin 
                      idxPages_25 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_26 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1a==waddr)
                    begin 
                      idxPages_26 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              idxPages_27 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1b==waddr)
                    begin 
                      idxPages_27 <=_idxPages_T[2:0];
                    end 
               end 
         if (metaReset)
            begin 
              tgts_0 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h0==waddr)
                    begin 
                      tgts_0 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_1 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1==waddr)
                    begin 
                      tgts_1 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_2 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h2==waddr)
                    begin 
                      tgts_2 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_3 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h3==waddr)
                    begin 
                      tgts_3 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_4 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h4==waddr)
                    begin 
                      tgts_4 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_5 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h5==waddr)
                    begin 
                      tgts_5 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_6 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h6==waddr)
                    begin 
                      tgts_6 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_7 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h7==waddr)
                    begin 
                      tgts_7 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_8 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h8==waddr)
                    begin 
                      tgts_8 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_9 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h9==waddr)
                    begin 
                      tgts_9 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_10 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'ha==waddr)
                    begin 
                      tgts_10 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_11 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hb==waddr)
                    begin 
                      tgts_11 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_12 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hc==waddr)
                    begin 
                      tgts_12 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_13 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hd==waddr)
                    begin 
                      tgts_13 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_14 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'he==waddr)
                    begin 
                      tgts_14 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_15 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hf==waddr)
                    begin 
                      tgts_15 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_16 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h10==waddr)
                    begin 
                      tgts_16 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_17 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h11==waddr)
                    begin 
                      tgts_17 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_18 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h12==waddr)
                    begin 
                      tgts_18 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_19 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h13==waddr)
                    begin 
                      tgts_19 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_20 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h14==waddr)
                    begin 
                      tgts_20 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_21 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h15==waddr)
                    begin 
                      tgts_21 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_22 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h16==waddr)
                    begin 
                      tgts_22 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_23 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h17==waddr)
                    begin 
                      tgts_23 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_24 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h18==waddr)
                    begin 
                      tgts_24 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_25 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h19==waddr)
                    begin 
                      tgts_25 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_26 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1a==waddr)
                    begin 
                      tgts_26 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgts_27 <=13'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1b==waddr)
                    begin 
                      tgts_27 <=idxHit_idx;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_0 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h0==waddr)
                    begin 
                      tgtPages_0 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_1 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1==waddr)
                    begin 
                      tgtPages_1 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_2 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h2==waddr)
                    begin 
                      tgtPages_2 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_3 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h3==waddr)
                    begin 
                      tgtPages_3 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_4 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h4==waddr)
                    begin 
                      tgtPages_4 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_5 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h5==waddr)
                    begin 
                      tgtPages_5 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_6 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h6==waddr)
                    begin 
                      tgtPages_6 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_7 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h7==waddr)
                    begin 
                      tgtPages_7 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_8 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h8==waddr)
                    begin 
                      tgtPages_8 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_9 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h9==waddr)
                    begin 
                      tgtPages_9 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_10 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'ha==waddr)
                    begin 
                      tgtPages_10 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_11 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hb==waddr)
                    begin 
                      tgtPages_11 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_12 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hc==waddr)
                    begin 
                      tgtPages_12 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_13 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hd==waddr)
                    begin 
                      tgtPages_13 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_14 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'he==waddr)
                    begin 
                      tgtPages_14 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_15 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hf==waddr)
                    begin 
                      tgtPages_15 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_16 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h10==waddr)
                    begin 
                      tgtPages_16 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_17 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h11==waddr)
                    begin 
                      tgtPages_17 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_18 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h12==waddr)
                    begin 
                      tgtPages_18 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_19 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h13==waddr)
                    begin 
                      tgtPages_19 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_20 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h14==waddr)
                    begin 
                      tgtPages_20 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_21 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h15==waddr)
                    begin 
                      tgtPages_21 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_22 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h16==waddr)
                    begin 
                      tgtPages_22 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_23 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h17==waddr)
                    begin 
                      tgtPages_23 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_24 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h18==waddr)
                    begin 
                      tgtPages_24 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_25 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h19==waddr)
                    begin 
                      tgtPages_25 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_26 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1a==waddr)
                    begin 
                      tgtPages_26 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              tgtPages_27 <=3'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1b==waddr)
                    begin 
                      tgtPages_27 <=tgtPageUpdate;
                    end 
               end 
         if (metaReset)
            begin 
              pages_0 <=25'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (_T_5[0])
                    begin 
                      if (idxWritesEven)
                         begin 
                           pages_0 <=updatePageHit_p;
                         end 
                       else 
                         begin 
                           pages_0 <=pageHit_p;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              pages_1 <=25'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (_T_12[1])
                    begin 
                      if (idxWritesEven)
                         begin 
                           pages_1 <=pageHit_p;
                         end 
                       else 
                         begin 
                           pages_1 <=updatePageHit_p;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              pages_2 <=25'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (_T_5[2])
                    begin 
                      if (idxWritesEven)
                         begin 
                           pages_2 <=updatePageHit_p;
                         end 
                       else 
                         begin 
                           pages_2 <=pageHit_p;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              pages_3 <=25'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (_T_12[3])
                    begin 
                      if (idxWritesEven)
                         begin 
                           pages_3 <=pageHit_p;
                         end 
                       else 
                         begin 
                           pages_3 <=updatePageHit_p;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              pages_4 <=25'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (_T_5[4])
                    begin 
                      if (idxWritesEven)
                         begin 
                           pages_4 <=updatePageHit_p;
                         end 
                       else 
                         begin 
                           pages_4 <=pageHit_p;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              pages_5 <=25'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (_T_12[5])
                    begin 
                      if (idxWritesEven)
                         begin 
                           pages_5 <=pageHit_p;
                         end 
                       else 
                         begin 
                           pages_5 <=updatePageHit_p;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              pageValid <=6'h0;
            end 
          else 
            if (reset)
               begin 
                 pageValid <=6'h0;
               end 
             else 
               begin 
                 pageValid <=_GEN_373[5:0];
               end 
         if (metaReset)
            begin 
              isValid <=28'h0;
            end 
          else 
            if (reset)
               begin 
                 isValid <=28'h0;
               end 
             else 
               begin 
                 isValid <=_GEN_375[27:0];
               end 
         if (metaReset)
            begin 
              cfiType_0 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h0==waddr)
                    begin 
                      cfiType_0 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_1 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1==waddr)
                    begin 
                      cfiType_1 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_2 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h2==waddr)
                    begin 
                      cfiType_2 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_3 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h3==waddr)
                    begin 
                      cfiType_3 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_4 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h4==waddr)
                    begin 
                      cfiType_4 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_5 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h5==waddr)
                    begin 
                      cfiType_5 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_6 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h6==waddr)
                    begin 
                      cfiType_6 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_7 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h7==waddr)
                    begin 
                      cfiType_7 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_8 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h8==waddr)
                    begin 
                      cfiType_8 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_9 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h9==waddr)
                    begin 
                      cfiType_9 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_10 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'ha==waddr)
                    begin 
                      cfiType_10 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_11 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hb==waddr)
                    begin 
                      cfiType_11 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_12 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hc==waddr)
                    begin 
                      cfiType_12 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_13 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hd==waddr)
                    begin 
                      cfiType_13 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_14 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'he==waddr)
                    begin 
                      cfiType_14 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_15 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hf==waddr)
                    begin 
                      cfiType_15 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_16 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h10==waddr)
                    begin 
                      cfiType_16 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_17 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h11==waddr)
                    begin 
                      cfiType_17 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_18 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h12==waddr)
                    begin 
                      cfiType_18 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_19 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h13==waddr)
                    begin 
                      cfiType_19 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_20 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h14==waddr)
                    begin 
                      cfiType_20 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_21 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h15==waddr)
                    begin 
                      cfiType_21 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_22 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h16==waddr)
                    begin 
                      cfiType_22 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_23 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h17==waddr)
                    begin 
                      cfiType_23 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_24 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h18==waddr)
                    begin 
                      cfiType_24 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_25 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h19==waddr)
                    begin 
                      cfiType_25 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_26 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1a==waddr)
                    begin 
                      cfiType_26 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              cfiType_27 <=2'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1b==waddr)
                    begin 
                      cfiType_27 <=r_btb_updatePipe_bits_cfiType;
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_0 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h0==waddr)
                    begin 
                      brIdx_0 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_1 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1==waddr)
                    begin 
                      brIdx_1 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_2 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h2==waddr)
                    begin 
                      brIdx_2 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_3 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h3==waddr)
                    begin 
                      brIdx_3 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_4 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h4==waddr)
                    begin 
                      brIdx_4 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_5 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h5==waddr)
                    begin 
                      brIdx_5 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_6 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h6==waddr)
                    begin 
                      brIdx_6 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_7 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h7==waddr)
                    begin 
                      brIdx_7 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_8 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h8==waddr)
                    begin 
                      brIdx_8 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_9 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h9==waddr)
                    begin 
                      brIdx_9 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_10 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'ha==waddr)
                    begin 
                      brIdx_10 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_11 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hb==waddr)
                    begin 
                      brIdx_11 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_12 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hc==waddr)
                    begin 
                      brIdx_12 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_13 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hd==waddr)
                    begin 
                      brIdx_13 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_14 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'he==waddr)
                    begin 
                      brIdx_14 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_15 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'hf==waddr)
                    begin 
                      brIdx_15 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_16 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h10==waddr)
                    begin 
                      brIdx_16 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_17 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h11==waddr)
                    begin 
                      brIdx_17 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_18 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h12==waddr)
                    begin 
                      brIdx_18 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_19 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h13==waddr)
                    begin 
                      brIdx_19 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_20 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h14==waddr)
                    begin 
                      brIdx_20 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_21 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h15==waddr)
                    begin 
                      brIdx_21 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_22 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h16==waddr)
                    begin 
                      brIdx_22 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_23 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h17==waddr)
                    begin 
                      brIdx_23 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_24 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h18==waddr)
                    begin 
                      brIdx_24 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_25 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h19==waddr)
                    begin 
                      brIdx_25 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_26 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1a==waddr)
                    begin 
                      brIdx_26 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              brIdx_27 <=1'h0;
            end 
          else 
            if (r_btb_updatePipe_valid)
               begin 
                 if (5'h1b==waddr)
                    begin 
                      brIdx_27 <=r_btb_updatePipe_bits_br_pc[1];
                    end 
               end 
         if (metaReset)
            begin 
              r_btb_updatePipe_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 r_btb_updatePipe_valid <=1'h0;
               end 
             else 
               begin 
                 r_btb_updatePipe_valid <=io_btb_update_valid;
               end 
         if (metaReset)
            begin 
              r_btb_updatePipe_bits_prediction_entry <=5'h0;
            end 
          else 
            if (io_btb_update_valid)
               begin 
                 r_btb_updatePipe_bits_prediction_entry <=io_btb_update_bits_prediction_entry;
               end 
         if (metaReset)
            begin 
              r_btb_updatePipe_bits_pc <=39'h0;
            end 
          else 
            if (io_btb_update_valid)
               begin 
                 r_btb_updatePipe_bits_pc <=io_btb_update_bits_pc;
               end 
         if (metaReset)
            begin 
              r_btb_updatePipe_bits_isValid <=1'h0;
            end 
          else 
            if (io_btb_update_valid)
               begin 
                 r_btb_updatePipe_bits_isValid <=io_btb_update_bits_isValid;
               end 
         if (metaReset)
            begin 
              r_btb_updatePipe_bits_br_pc <=39'h0;
            end 
          else 
            if (io_btb_update_valid)
               begin 
                 r_btb_updatePipe_bits_br_pc <=io_btb_update_bits_br_pc;
               end 
         if (metaReset)
            begin 
              r_btb_updatePipe_bits_cfiType <=2'h0;
            end 
          else 
            if (io_btb_update_valid)
               begin 
                 r_btb_updatePipe_bits_cfiType <=io_btb_update_bits_cfiType;
               end 
         if (metaReset)
            begin 
              nextPageRepl <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 nextPageRepl <=3'h0;
               end 
             else 
               if (_T_1)
                  begin 
                    if (_nextPageRepl_T)
                       begin 
                         nextPageRepl <={2'b0,next[0]};
                       end 
                     else 
                       begin 
                         nextPageRepl <=next;
                       end 
                  end 
         if (metaReset)
            begin 
              state_reg <=27'h0;
            end 
          else 
            if (reset)
               begin 
                 state_reg <=27'h0;
               end 
             else 
               if (_T_3)
                  begin 
                    state_reg <=_state_reg_T_66;
                  end 
         if (metaReset)
            begin 
              r_respPipe_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 r_respPipe_valid <=1'h0;
               end 
             else 
               begin 
                 r_respPipe_valid <=io_resp_valid;
               end 
         if (metaReset)
            begin 
              r_respPipe_bits_taken <=1'h0;
            end 
          else 
            if (io_resp_valid)
               begin 
                 r_respPipe_bits_taken <=io_resp_bits_taken;
               end 
         if (metaReset)
            begin 
              r_respPipe_bits_entry <=5'h0;
            end 
          else 
            if (io_resp_valid)
               begin 
                 r_respPipe_bits_entry <=io_resp_bits_entry;
               end 
         if (metaReset)
            begin 
              history <=8'h0;
            end 
          else 
            if (reset)
               begin 
                 history <=8'h0;
               end 
             else 
               if (io_bht_update_valid)
                  begin 
                    if (io_bht_update_bits_branch)
                       begin 
                         if (io_bht_update_bits_mispredict)
                            begin 
                              history <=_history_T_1;
                            end 
                          else 
                            if (io_bht_advance_valid)
                               begin 
                                 history <=_history_T;
                               end 
                       end 
                     else 
                       if (io_bht_update_bits_mispredict)
                          begin 
                            history <=io_bht_update_bits_prediction_history;
                          end 
                        else 
                          if (io_bht_advance_valid)
                             begin 
                               history <=_history_T;
                             end 
                  end 
                else 
                  if (io_bht_advance_valid)
                     begin 
                       history <=_history_T;
                     end 
         if (metaReset)
            begin 
              reset_waddr <=10'h0;
            end 
          else 
            if (reset)
               begin 
                 reset_waddr <=10'h0;
               end 
             else 
               if (resetting)
                  begin 
                    reset_waddr <=_reset_waddr_T_1;
                  end 
         if (metaReset)
            begin 
              count <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 count <=3'h0;
               end 
             else 
               if (io_ras_update_valid)
                  begin 
                    if (_T_138)
                       begin 
                         if (_T_139)
                            begin 
                              count <=_count_T_1;
                            end 
                       end 
                     else 
                       if (_T_140)
                          begin 
                            if (~_io_ras_head_valid_T)
                               begin 
                                 count <=_count_T_3;
                               end 
                          end 
                  end 
         if (metaReset)
            begin 
              pos <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 pos <=3'h0;
               end 
             else 
               if (io_ras_update_valid)
                  begin 
                    if (_T_138)
                       begin 
                         if (_nextPos_T)
                            begin 
                              pos <=_nextPos_T_3;
                            end 
                          else 
                            begin 
                              pos <=3'h0;
                            end 
                       end 
                     else 
                       if (_T_140)
                          begin 
                            if (~_io_ras_head_valid_T)
                               begin 
                                 if (_pos_T)
                                    begin 
                                      pos <=_pos_T_3;
                                    end 
                                  else 
                                    begin 
                                      pos <=3'h5;
                                    end 
                               end 
                          end 
                  end 
         if (metaReset)
            begin 
              stack_0 <=39'h0;
            end 
          else 
            if (io_ras_update_valid)
               begin 
                 if (_T_138)
                    begin 
                      if (3'h0==nextPos)
                         begin 
                           stack_0 <=io_ras_update_bits_returnAddr;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              stack_1 <=39'h0;
            end 
          else 
            if (io_ras_update_valid)
               begin 
                 if (_T_138)
                    begin 
                      if (3'h1==nextPos)
                         begin 
                           stack_1 <=io_ras_update_bits_returnAddr;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              stack_2 <=39'h0;
            end 
          else 
            if (io_ras_update_valid)
               begin 
                 if (_T_138)
                    begin 
                      if (3'h2==nextPos)
                         begin 
                           stack_2 <=io_ras_update_bits_returnAddr;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              stack_3 <=39'h0;
            end 
          else 
            if (io_ras_update_valid)
               begin 
                 if (_T_138)
                    begin 
                      if (3'h3==nextPos)
                         begin 
                           stack_3 <=io_ras_update_bits_returnAddr;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              stack_4 <=39'h0;
            end 
          else 
            if (io_ras_update_valid)
               begin 
                 if (_T_138)
                    begin 
                      if (3'h4==nextPos)
                         begin 
                           stack_4 <=io_ras_update_bits_returnAddr;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              stack_5 <=39'h0;
            end 
          else 
            if (io_ras_update_valid)
               begin 
                 if (_T_138)
                    begin 
                      if (3'h5==nextPos)
                         begin 
                           stack_5 <=io_ras_update_bits_returnAddr;
                         end 
                    end 
               end 
         BTB_state <=BTB_xor0;
         if (!(BTB_cov_read_data))
            begin 
              BTB_covSum <=BTB_covSum+1'h1;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (BTB_cov_write_en&BTB_cov_write_mask)
            begin 
              BTB_cov [BTB_cov_write_addr]<=BTB_cov_write_data;
            end 
       end
  
endmodule
 
module FPUDecoder (
  input [31:0] io_inst,
  output io_sigs_wen,
  output io_sigs_ren1,
  output io_sigs_ren2,
  output io_sigs_ren3,
  output io_sigs_swap12,
  output io_sigs_swap23,
  output [1:0] io_sigs_typeTagIn,
  output [1:0] io_sigs_typeTagOut,
  output io_sigs_fromint,
  output io_sigs_toint,
  output io_sigs_fastpipe,
  output io_sigs_fma,
  output io_sigs_div,
  output io_sigs_sqrt,
  output io_sigs_wflags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [31:0] _decoder_T ;  
   wire decoder_0 ;  
   wire [31:0] _decoder_T_2 ;  
   wire _decoder_T_3 ;  
   wire [31:0] _decoder_T_4 ;  
   wire _decoder_T_5 ;  
   wire [31:0] _decoder_T_6 ;  
   wire _decoder_T_7 ;  
   wire _decoder_T_9 ;  
   wire [31:0] _decoder_T_10 ;  
   wire _decoder_T_11 ;  
   wire [31:0] _decoder_T_12 ;  
   wire _decoder_T_13 ;  
   wire [31:0] _decoder_T_14 ;  
   wire decoder_4 ;  
   wire _decoder_T_17 ;  
   wire [31:0] _decoder_T_18 ;  
   wire _decoder_T_19 ;  
   wire [31:0] _decoder_T_20 ;  
   wire _decoder_T_21 ;  
   wire _decoder_T_23 ;  
   wire [31:0] _decoder_T_24 ;  
   wire [31:0] _decoder_T_26 ;  
   wire _decoder_T_27 ;  
   wire [31:0] _decoder_T_28 ;  
   wire _decoder_T_29 ;  
   wire [31:0] _decoder_T_30 ;  
   wire _decoder_T_31 ;  
   wire [31:0] _decoder_T_32 ;  
   wire _decoder_T_33 ;  
   wire [31:0] _decoder_T_34 ;  
   wire _decoder_T_35 ;  
   wire [31:0] _decoder_T_36 ;  
   wire _decoder_T_37 ;  
   wire _decoder_T_39 ;  
   wire _decoder_T_40 ;  
   wire _decoder_T_41 ;  
   wire _decoder_T_42 ;  
   wire _decoder_T_43 ;  
   wire decoder_7 ;  
   wire [31:0] _decoder_T_44 ;  
   wire _decoder_T_45 ;  
   wire [31:0] _decoder_T_46 ;  
   wire _decoder_T_47 ;  
   wire _decoder_T_49 ;  
   wire _decoder_T_51 ;  
   wire decoder_8 ;  
   wire [31:0] _decoder_T_52 ;  
   wire _decoder_T_55 ;  
   wire [31:0] _decoder_T_57 ;  
   wire _decoder_T_58 ;  
   wire [31:0] _decoder_T_59 ;  
   wire _decoder_T_60 ;  
   wire [31:0] _decoder_T_62 ;  
   wire _decoder_T_63 ;  
   wire [31:0] _decoder_T_64 ;  
   wire _decoder_T_65 ;  
   wire _decoder_T_67 ;  
   wire [31:0] _decoder_T_68 ;  
   wire [31:0] _decoder_T_72 ;  
   wire _decoder_T_73 ;  
   wire [31:0] _decoder_T_74 ;  
   wire _decoder_T_75 ;  
   wire [31:0] _decoder_T_76 ;  
   wire _decoder_T_77 ;  
   wire _decoder_T_79 ;  
   wire _decoder_T_80 ;  
   wire [29:0] FPUDecoder_covSum ;  
  assign _decoder_T=io_inst&32'h40; 
  assign decoder_0=_decoder_T==32'h0; 
  assign _decoder_T_2=io_inst&32'h80000020; 
  assign _decoder_T_3=_decoder_T_2==32'h0; 
  assign _decoder_T_4=io_inst&32'h30; 
  assign _decoder_T_5=_decoder_T_4==32'h0; 
  assign _decoder_T_6=io_inst&32'h10000020; 
  assign _decoder_T_7=_decoder_T_6==32'h10000000; 
  assign _decoder_T_9=_decoder_T_3|_decoder_T_5; 
  assign _decoder_T_10=io_inst&32'h80000004; 
  assign _decoder_T_11=_decoder_T_10==32'h0; 
  assign _decoder_T_12=io_inst&32'h10000004; 
  assign _decoder_T_13=_decoder_T_12==32'h0; 
  assign _decoder_T_14=io_inst&32'h50; 
  assign decoder_4=_decoder_T_14==32'h40; 
  assign _decoder_T_17=_decoder_T_11|_decoder_T_13; 
  assign _decoder_T_18=io_inst&32'h40000004; 
  assign _decoder_T_19=_decoder_T_18==32'h0; 
  assign _decoder_T_20=io_inst&32'h20; 
  assign _decoder_T_21=_decoder_T_20==32'h20; 
  assign _decoder_T_23=_decoder_T_19|_decoder_T_21; 
  assign _decoder_T_24=io_inst&32'h30000010; 
  assign _decoder_T_26=io_inst&32'h42000000; 
  assign _decoder_T_27=_decoder_T_26==32'h2000000; 
  assign _decoder_T_28=io_inst&32'h2000010; 
  assign _decoder_T_29=_decoder_T_28==32'h2000000; 
  assign _decoder_T_30=io_inst&32'h12000000; 
  assign _decoder_T_31=_decoder_T_30==32'h12000000; 
  assign _decoder_T_32=io_inst&32'hd2000010; 
  assign _decoder_T_33=_decoder_T_32==32'h40000010; 
  assign _decoder_T_34=io_inst&32'h70001010; 
  assign _decoder_T_35=_decoder_T_34==32'h60000010; 
  assign _decoder_T_36=io_inst&32'h82000000; 
  assign _decoder_T_37=_decoder_T_36==32'h82000000; 
  assign _decoder_T_39=decoder_0|_decoder_T_27; 
  assign _decoder_T_40=_decoder_T_39|_decoder_T_29; 
  assign _decoder_T_41=_decoder_T_40|_decoder_T_31; 
  assign _decoder_T_42=_decoder_T_41|_decoder_T_33; 
  assign _decoder_T_43=_decoder_T_42|_decoder_T_35; 
  assign decoder_7=_decoder_T_43|_decoder_T_37; 
  assign _decoder_T_44=io_inst&32'h1040; 
  assign _decoder_T_45=_decoder_T_44==32'h1000; 
  assign _decoder_T_46=io_inst&32'h2000020; 
  assign _decoder_T_47=_decoder_T_46==32'h2000000; 
  assign _decoder_T_49=_decoder_T_24==32'h30000010; 
  assign _decoder_T_51=_decoder_T_45|_decoder_T_47; 
  assign decoder_8=_decoder_T_51|_decoder_T_49; 
  assign _decoder_T_52=io_inst&32'h90000010; 
  assign _decoder_T_55=_decoder_T_52==32'h80000010; 
  assign _decoder_T_57=io_inst&32'ha0000010; 
  assign _decoder_T_58=_decoder_T_57==32'h20000010; 
  assign _decoder_T_59=io_inst&32'hd0000010; 
  assign _decoder_T_60=_decoder_T_59==32'h40000010; 
  assign _decoder_T_62=io_inst&32'h70000004; 
  assign _decoder_T_63=_decoder_T_62==32'h0; 
  assign _decoder_T_64=io_inst&32'h68000004; 
  assign _decoder_T_65=_decoder_T_64==32'h0; 
  assign _decoder_T_67=_decoder_T_63|_decoder_T_65; 
  assign _decoder_T_68=io_inst&32'h58000010; 
  assign _decoder_T_72=io_inst&32'h20000004; 
  assign _decoder_T_73=_decoder_T_72==32'h0; 
  assign _decoder_T_74=io_inst&32'h8002000; 
  assign _decoder_T_75=_decoder_T_74==32'h8000000; 
  assign _decoder_T_76=io_inst&32'hc0000004; 
  assign _decoder_T_77=_decoder_T_76==32'h80000000; 
  assign _decoder_T_79=_decoder_T_73|decoder_4; 
  assign _decoder_T_80=_decoder_T_79|_decoder_T_75; 
  assign io_sigs_wen=_decoder_T_9|_decoder_T_7; 
  assign io_sigs_ren1=_decoder_T_17|decoder_4; 
  assign io_sigs_ren2=_decoder_T_23|decoder_4; 
  assign io_sigs_ren3=_decoder_T_14==32'h40; 
  assign io_sigs_swap12=_decoder_T==32'h0; 
  assign io_sigs_swap23=_decoder_T_24==32'h10; 
  assign io_sigs_typeTagIn={1'b0,decoder_7}; 
  assign io_sigs_typeTagOut={1'b0,decoder_8}; 
  assign io_sigs_fromint=_decoder_T_52==32'h90000010; 
  assign io_sigs_toint=_decoder_T_21|_decoder_T_55; 
  assign io_sigs_fastpipe=_decoder_T_58|_decoder_T_60; 
  assign io_sigs_fma=_decoder_T_67|decoder_4; 
  assign io_sigs_div=_decoder_T_68==32'h18000010; 
  assign io_sigs_sqrt=_decoder_T_59==32'h50000010; 
  assign io_sigs_wflags=_decoder_T_80|_decoder_T_77; 
  assign FPUDecoder_covSum=30'h0; 
  assign io_covSum=FPUDecoder_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module FPUFMAPipe (
  input clock,
  input reset,
  input io_in_valid,
  input io_in_bits_ren3,
  input io_in_bits_swap23,
  input [2:0] io_in_bits_rm,
  input [1:0] io_in_bits_fmaCmd,
  input [64:0] io_in_bits_in1,
  input [64:0] io_in_bits_in2,
  input [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input fma_halt) ; 
   wire fma_clock ;  
   wire fma_reset ;  
   wire fma_io_validin ;  
   wire [1:0] fma_io_op ;  
   wire [32:0] fma_io_a ;  
   wire [32:0] fma_io_b ;  
   wire [32:0] fma_io_c ;  
   wire [2:0] fma_io_roundingMode ;  
   wire [32:0] fma_io_out ;  
   wire [4:0] fma_io_exceptionFlags ;  
   wire [29:0] fma_io_covSum ;  
   wire fma_metaAssert ;  
   wire fma_metaReset ;  
   reg valid ;  
   reg [31:0] _RAND_0 ;  
   reg [2:0] in_rm ;  
   reg [31:0] _RAND_1 ;  
   reg [1:0] in_fmaCmd ;  
   reg [31:0] _RAND_2 ;  
   reg [64:0] in_in1 ;  
   reg [95:0] _RAND_3 ;  
   reg [64:0] in_in2 ;  
   reg [95:0] _RAND_4 ;  
   reg [64:0] in_in3 ;  
   reg [95:0] _RAND_5 ;  
   wire [64:0] _zero_T ;  
   wire [64:0] zero ;  
   wire _T ;  
   wire [29:0] FPUFMAPipe_covSum ;  
   wire [29:0] fma_sum ;  
   wire fma_metaAssert_wire ;  
   reg FPUFMAPipe_metaAssert ;  
   reg [31:0] _RAND_6 ;  
  MulAddRecFNPipe fma(.clock(fma_clock),.reset(fma_reset),.io_validin(fma_io_validin),.io_op(fma_io_op),.io_a(fma_io_a),.io_b(fma_io_b),.io_c(fma_io_c),.io_roundingMode(fma_io_roundingMode),.io_out(fma_io_out),.io_exceptionFlags(fma_io_exceptionFlags),.io_covSum(fma_io_covSum),.metaAssert(fma_metaAssert),.metaReset(fma_metaReset)); 
  assign _zero_T=io_in_bits_in1^io_in_bits_in2; 
  assign zero=_zero_T&65'h100000000; 
  assign _T=io_in_bits_ren3|io_in_bits_swap23; 
  assign io_out_bits_data={32'b0,fma_io_out}; 
  assign io_out_bits_exc=fma_io_exceptionFlags; 
  assign fma_clock=clock; 
  assign fma_reset=reset; 
  assign fma_io_validin=valid; 
  assign fma_io_op=in_fmaCmd; 
  assign fma_io_a=in_in1[32:0]; 
  assign fma_io_b=in_in2[32:0]; 
  assign fma_io_c=in_in3[32:0]; 
  assign fma_io_roundingMode=in_rm; 
  assign FPUFMAPipe_covSum=30'h0; 
  assign fma_sum=FPUFMAPipe_covSum+fma_io_covSum; 
  assign io_covSum=fma_sum; 
  assign fma_metaAssert_wire=fma_metaAssert; 
  assign metaAssert=FPUFMAPipe_metaAssert; 
  assign fma_metaReset=metaReset|fma_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              valid <=1'h0;
            end 
          else 
            begin 
              valid <=io_in_valid;
            end 
         if (metaReset)
            begin 
              in_rm <=3'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_rm <=io_in_bits_rm;
               end 
         if (metaReset)
            begin 
              in_fmaCmd <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_fmaCmd <=io_in_bits_fmaCmd;
               end 
         if (metaReset)
            begin 
              in_in1 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_in1 <=io_in_bits_in1;
               end 
         if (metaReset)
            begin 
              in_in2 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 if (io_in_bits_swap23)
                    begin 
                      in_in2 <=65'h80000000;
                    end 
                  else 
                    begin 
                      in_in2 <=io_in_bits_in2;
                    end 
               end 
         if (metaReset)
            begin 
              in_in3 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 if (~_T)
                    begin 
                      in_in3 <=zero;
                    end 
                  else 
                    begin 
                      in_in3 <=io_in_bits_in3;
                    end 
               end 
         if (metaReset)
            begin 
              FPUFMAPipe_metaAssert <=1'h0;
            end 
          else 
            begin 
              FPUFMAPipe_metaAssert <=FPUFMAPipe_metaAssert|fma_metaAssert_wire;
            end 
       end
  
endmodule
 
module FPToInt (
  input clock,
  input io_in_valid,
  input io_in_bits_ren2,
  input [1:0] io_in_bits_typeTagIn,
  input [1:0] io_in_bits_typeTagOut,
  input io_in_bits_wflags,
  input [2:0] io_in_bits_rm,
  input [1:0] io_in_bits_typ,
  input [1:0] io_in_bits_fmt,
  input [64:0] io_in_bits_in1,
  input [64:0] io_in_bits_in2,
  output [2:0] io_out_bits_in_rm,
  output [64:0] io_out_bits_in_in1,
  output [64:0] io_out_bits_in_in2,
  output io_out_bits_lt,
  output [63:0] io_out_bits_store,
  output [63:0] io_out_bits_toint,
  output [4:0] io_out_bits_exc,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [64:0] dcmp_io_a ;  
   wire [64:0] dcmp_io_b ;  
   wire dcmp_io_signaling ;  
   wire dcmp_io_lt ;  
   wire dcmp_io_eq ;  
   wire [4:0] dcmp_io_exceptionFlags ;  
   wire [29:0] dcmp_io_covSum ;  
   wire dcmp_metaAssert ;  
   wire [64:0] conv_io_in ;  
   wire [2:0] conv_io_roundingMode ;  
   wire conv_io_signedOut ;  
   wire [63:0] conv_io_out ;  
   wire [2:0] conv_io_intExceptionFlags ;  
   wire [29:0] conv_io_covSum ;  
   wire conv_metaAssert ;  
   wire [64:0] narrow_io_in ;  
   wire [2:0] narrow_io_roundingMode ;  
   wire narrow_io_signedOut ;  
   wire [2:0] narrow_io_intExceptionFlags ;  
   wire [29:0] narrow_io_covSum ;  
   wire narrow_metaAssert ;  
   reg in_ren2 ;  
   reg [31:0] _RAND_0 ;  
   reg [1:0] in_typeTagOut ;  
   reg [31:0] _RAND_1 ;  
   reg in_wflags ;  
   reg [31:0] _RAND_2 ;  
   reg [2:0] in_rm ;  
   reg [31:0] _RAND_3 ;  
   reg [1:0] in_typ ;  
   reg [31:0] _RAND_4 ;  
   reg [1:0] in_fmt ;  
   reg [31:0] _RAND_5 ;  
   reg [64:0] in_in1 ;  
   reg [95:0] _RAND_6 ;  
   reg [64:0] in_in2 ;  
   reg [95:0] _RAND_7 ;  
   wire [11:0] store_unrecoded_rawIn_exp ;  
   wire store_unrecoded_rawIn_isZero ;  
   wire store_unrecoded_rawIn_isSpecial ;  
   wire store_unrecoded_rawIn__isNaN ;  
   wire store_unrecoded_rawIn__isInf ;  
   wire store_unrecoded_rawIn__sign ;  
   wire [12:0] store_unrecoded_rawIn__sExp ;  
   wire store_unrecoded_rawIn_out_sig_hi_lo ;  
   wire [51:0] store_unrecoded_rawIn_out_sig_lo ;  
   wire [53:0] store_unrecoded_rawIn__sig ;  
   wire store_unrecoded_isSubnormal ;  
   wire [5:0] store_unrecoded_denormShiftDist ;  
   wire [52:0] _store_unrecoded_denormFract_T_1 ;  
   wire [51:0] store_unrecoded_denormFract ;  
   wire [10:0] _store_unrecoded_expOut_T_2 ;  
   wire [10:0] _store_unrecoded_expOut_T_3 ;  
   wire _store_unrecoded_expOut_T_4 ;  
   wire [10:0] _store_unrecoded_expOut_T_6 ;  
   wire [10:0] store_unrecoded_hi_lo ;  
   wire [51:0] _store_unrecoded_fractOut_T_1 ;  
   wire [51:0] store_unrecoded_lo ;  
   wire [63:0] store_unrecoded ;  
   wire store_prevRecoded_hi_hi ;  
   wire store_prevRecoded_hi_lo ;  
   wire [30:0] store_prevRecoded_lo ;  
   wire [32:0] store_prevRecoded ;  
   wire [8:0] store_prevUnrecoded_rawIn_exp ;  
   wire store_prevUnrecoded_rawIn_isZero ;  
   wire store_prevUnrecoded_rawIn_isSpecial ;  
   wire store_prevUnrecoded_rawIn__isNaN ;  
   wire store_prevUnrecoded_rawIn__isInf ;  
   wire store_prevUnrecoded_rawIn__sign ;  
   wire [9:0] store_prevUnrecoded_rawIn__sExp ;  
   wire store_prevUnrecoded_rawIn_out_sig_hi_lo ;  
   wire [22:0] store_prevUnrecoded_rawIn_out_sig_lo ;  
   wire [24:0] store_prevUnrecoded_rawIn__sig ;  
   wire store_prevUnrecoded_isSubnormal ;  
   wire [4:0] store_prevUnrecoded_denormShiftDist ;  
   wire [23:0] _store_prevUnrecoded_denormFract_T_1 ;  
   wire [22:0] store_prevUnrecoded_denormFract ;  
   wire [7:0] _store_prevUnrecoded_expOut_T_2 ;  
   wire [7:0] _store_prevUnrecoded_expOut_T_3 ;  
   wire _store_prevUnrecoded_expOut_T_4 ;  
   wire [7:0] _store_prevUnrecoded_expOut_T_6 ;  
   wire [7:0] store_prevUnrecoded_hi_lo ;  
   wire [22:0] _store_prevUnrecoded_fractOut_T_1 ;  
   wire [22:0] store_prevUnrecoded_lo ;  
   wire [31:0] store_prevUnrecoded ;  
   wire [31:0] store_hi ;  
   wire _store_T_1 ;  
   wire [31:0] store_lo ;  
   wire [63:0] _store_T_3 ;  
   wire [31:0] store_hi_1 ;  
   wire [63:0] _store_T_4 ;  
   wire store_truncIdx ;  
   wire [63:0] store ;  
   wire intType_x6 ;  
   wire cvtType ;  
   wire io_out_bits_exc_hi_hi_1 ;  
   wire [31:0] toint_hi ;  
   wire excSign ;  
   wire excOut_hi ;  
   wire [30:0] excOut_lo ;  
   wire [63:0] _toint_T_10 ;  
   wire [63:0] _GEN_25 ;  
   wire [63:0] _GEN_26 ;  
   wire [1:0] _toint_T_4 ;  
   wire [2:0] _GEN_34 ;  
   wire [2:0] _toint_T_5 ;  
   wire _toint_T_6 ;  
   wire [63:0] _toint_T_8 ;  
   wire [63:0] _GEN_35 ;  
   wire [63:0] _toint_T_9 ;  
   wire [63:0] _GEN_29 ;  
   wire classify_out_hi_hi_hi_hi_1 ;  
   wire classify_out_hi_hi_hi_lo_1 ;  
   wire [1:0] classify_out_codeHi_1 ;  
   wire classify_out_isSpecial_1 ;  
   wire classify_out_isInf_1 ;  
   wire classify_out_hi_hi_lo_1 ;  
   wire _classify_out_isNormal_T_4 ;  
   wire classify_out_isHighSubnormalIn_1 ;  
   wire _classify_out_isNormal_T_6 ;  
   wire _classify_out_isNormal_T_7 ;  
   wire classify_out_isNormal_1 ;  
   wire classify_out_hi_lo_hi_1 ;  
   wire _classify_out_isSubnormal_T_3 ;  
   wire _classify_out_isSubnormal_T_5 ;  
   wire classify_out_isSubnormal_1 ;  
   wire classify_out_hi_lo_lo_1 ;  
   wire classify_out_isZero_1 ;  
   wire classify_out_lo_hi_hi_hi_1 ;  
   wire classify_out_lo_hi_hi_lo_1 ;  
   wire classify_out_lo_hi_lo_1 ;  
   wire classify_out_lo_lo_hi_1 ;  
   wire classify_out_lo_lo_lo_1 ;  
   wire [9:0] _classify_out_T_10 ;  
   wire _classify_out_expOut_T_1 ;  
   wire _classify_out_expOut_T_2 ;  
   wire [11:0] _classify_out_expOut_commonCase_T_1 ;  
   wire [11:0] classify_out_expOut_commonCase ;  
   wire [5:0] classify_out_expOut_lo ;  
   wire [8:0] _classify_out_expOut_T_3 ;  
   wire [8:0] classify_out_hi_lo ;  
   wire [75:0] _classify_out_fractOut_T ;  
   wire [22:0] classify_out_lo ;  
   wire [32:0] _classify_out_T ;  
   wire [2:0] classify_out_code ;  
   wire classify_out_isNaN ;  
   wire classify_out_hi_hi_hi_hi ;  
   wire classify_out_hi_hi_hi_lo ;  
   wire [1:0] classify_out_codeHi ;  
   wire classify_out_isSpecial ;  
   wire classify_out_isInf ;  
   wire classify_out_sign ;  
   wire classify_out_hi_hi_lo ;  
   wire _classify_out_isNormal_T ;  
   wire classify_out_isHighSubnormalIn ;  
   wire _classify_out_isNormal_T_2 ;  
   wire _classify_out_isNormal_T_3 ;  
   wire classify_out_isNormal ;  
   wire classify_out_hi_lo_hi ;  
   wire _classify_out_isSubnormal_T ;  
   wire _classify_out_isSubnormal_T_2 ;  
   wire classify_out_isSubnormal ;  
   wire classify_out_hi_lo_lo ;  
   wire classify_out_isZero ;  
   wire classify_out_lo_hi_hi_hi ;  
   wire classify_out_lo_hi_hi_lo ;  
   wire classify_out_lo_hi_lo ;  
   wire classify_out_lo_lo_hi ;  
   wire classify_out_lo_lo_lo ;  
   wire [9:0] _classify_out_T_5 ;  
   wire [9:0] classify_out ;  
   wire [63:0] _GEN_36 ;  
   wire [63:0] _toint_T_2 ;  
   wire [63:0] _GEN_23 ;  
   wire [63:0] toint ;  
   wire [31:0] io_out_bits_toint_lo ;  
   wire [31:0] io_out_bits_toint_hi ;  
   wire [63:0] _io_out_bits_toint_T_2 ;  
   wire _GEN_28 ;  
   wire _GEN_24 ;  
   wire intType ;  
   wire io_out_bits_exc_hi_hi ;  
   wire io_out_bits_exc_lo ;  
   wire [4:0] _io_out_bits_exc_T_1 ;  
   wire io_out_bits_exc_lo_1 ;  
   wire [4:0] _io_out_bits_exc_T_4 ;  
   wire [4:0] _GEN_27 ;  
   wire [4:0] _GEN_30 ;  
   wire _io_out_bits_lt_T_1 ;  
   wire _io_out_bits_lt_T_3 ;  
   wire _io_out_bits_lt_T_4 ;  
   reg [3:0] FPToInt_state ;  
   reg [31:0] _RAND_8 ;  
   reg FPToInt_cov[0:15] ;  
   reg [31:0] _RAND_9 ;  
   wire FPToInt_cov_read_data ;  
   wire [3:0] FPToInt_cov_read_addr ;  
   wire FPToInt_cov_write_data ;  
   wire [3:0] FPToInt_cov_write_addr ;  
   wire FPToInt_cov_write_mask ;  
   wire FPToInt_cov_write_en ;  
   reg [29:0] FPToInt_covSum ;  
   reg [31:0] _RAND_10 ;  
   wire in_wflags_shl ;  
   wire [3:0] in_wflags_pad ;  
   wire [2:0] in_typ_shl ;  
   wire [3:0] in_typ_pad ;  
   wire [3:0] in_ren2_shl ;  
   wire [3:0] in_ren2_pad ;  
   wire [3:0] FPToInt_xor2 ;  
   wire [3:0] FPToInt_xor0 ;  
   wire [29:0] dcmp_sum ;  
   wire [29:0] conv_sum ;  
   wire [29:0] narrow_sum ;  
   wire dcmp_metaAssert_wire ;  
   wire conv_metaAssert_wire ;  
   wire narrow_metaAssert_wire ;  
   wire FPToInt_or2 ;  
   wire FPToInt_or0 ;  
  CompareRecFN dcmp(.io_a(dcmp_io_a),.io_b(dcmp_io_b),.io_signaling(dcmp_io_signaling),.io_lt(dcmp_io_lt),.io_eq(dcmp_io_eq),.io_exceptionFlags(dcmp_io_exceptionFlags),.io_covSum(dcmp_io_covSum),.metaAssert(dcmp_metaAssert)); 
  RecFNToIN conv(.io_in(conv_io_in),.io_roundingMode(conv_io_roundingMode),.io_signedOut(conv_io_signedOut),.io_out(conv_io_out),.io_intExceptionFlags(conv_io_intExceptionFlags),.io_covSum(conv_io_covSum),.metaAssert(conv_metaAssert)); 
  RecFNToIN_1 narrow(.io_in(narrow_io_in),.io_roundingMode(narrow_io_roundingMode),.io_signedOut(narrow_io_signedOut),.io_intExceptionFlags(narrow_io_intExceptionFlags),.io_covSum(narrow_io_covSum),.metaAssert(narrow_metaAssert)); 
  assign store_unrecoded_rawIn_exp=in_in1[63:52]; 
  assign store_unrecoded_rawIn_isZero=store_unrecoded_rawIn_exp[11:9]==3'h0; 
  assign store_unrecoded_rawIn_isSpecial=store_unrecoded_rawIn_exp[11:10]==2'h3; 
  assign store_unrecoded_rawIn__isNaN=store_unrecoded_rawIn_isSpecial&store_unrecoded_rawIn_exp[9]; 
  assign store_unrecoded_rawIn__isInf=store_unrecoded_rawIn_isSpecial&~store_unrecoded_rawIn_exp[9]; 
  assign store_unrecoded_rawIn__sign=in_in1[64]; 
  assign store_unrecoded_rawIn__sExp={1'b0,$signed(store_unrecoded_rawIn_exp)}; 
  assign store_unrecoded_rawIn_out_sig_hi_lo=~store_unrecoded_rawIn_isZero; 
  assign store_unrecoded_rawIn_out_sig_lo=in_in1[51:0]; 
  assign store_unrecoded_rawIn__sig={1'h0,store_unrecoded_rawIn_out_sig_hi_lo,store_unrecoded_rawIn_out_sig_lo}; 
  assign store_unrecoded_isSubnormal=$signed(store_unrecoded_rawIn__sExp)<13'sh402; 
  assign store_unrecoded_denormShiftDist=6'h1-store_unrecoded_rawIn__sExp[5:0]; 
  assign _store_unrecoded_denormFract_T_1=store_unrecoded_rawIn__sig[53:1]>>store_unrecoded_denormShiftDist; 
  assign store_unrecoded_denormFract=_store_unrecoded_denormFract_T_1[51:0]; 
  assign _store_unrecoded_expOut_T_2=store_unrecoded_rawIn__sExp[10:0]-11'h401; 
  assign _store_unrecoded_expOut_T_3=store_unrecoded_isSubnormal ? 11'h0:_store_unrecoded_expOut_T_2; 
  assign _store_unrecoded_expOut_T_4=store_unrecoded_rawIn__isNaN|store_unrecoded_rawIn__isInf; 
  assign _store_unrecoded_expOut_T_6=_store_unrecoded_expOut_T_4 ? 11'h7ff:11'h0; 
  assign store_unrecoded_hi_lo=_store_unrecoded_expOut_T_3|_store_unrecoded_expOut_T_6; 
  assign _store_unrecoded_fractOut_T_1=store_unrecoded_rawIn__isInf ? 52'h0:store_unrecoded_rawIn__sig[51:0]; 
  assign store_unrecoded_lo=store_unrecoded_isSubnormal ? store_unrecoded_denormFract:_store_unrecoded_fractOut_T_1; 
  assign store_unrecoded={store_unrecoded_rawIn__sign,store_unrecoded_hi_lo,store_unrecoded_lo}; 
  assign store_prevRecoded_hi_hi=in_in1[31]; 
  assign store_prevRecoded_hi_lo=in_in1[52]; 
  assign store_prevRecoded_lo=in_in1[30:0]; 
  assign store_prevRecoded={store_prevRecoded_hi_hi,store_prevRecoded_hi_lo,store_prevRecoded_lo}; 
  assign store_prevUnrecoded_rawIn_exp=store_prevRecoded[31:23]; 
  assign store_prevUnrecoded_rawIn_isZero=store_prevUnrecoded_rawIn_exp[8:6]==3'h0; 
  assign store_prevUnrecoded_rawIn_isSpecial=store_prevUnrecoded_rawIn_exp[8:7]==2'h3; 
  assign store_prevUnrecoded_rawIn__isNaN=store_prevUnrecoded_rawIn_isSpecial&store_prevUnrecoded_rawIn_exp[6]; 
  assign store_prevUnrecoded_rawIn__isInf=store_prevUnrecoded_rawIn_isSpecial&~store_prevUnrecoded_rawIn_exp[6]; 
  assign store_prevUnrecoded_rawIn__sign=store_prevRecoded[32]; 
  assign store_prevUnrecoded_rawIn__sExp={1'b0,$signed(store_prevUnrecoded_rawIn_exp)}; 
  assign store_prevUnrecoded_rawIn_out_sig_hi_lo=~store_prevUnrecoded_rawIn_isZero; 
  assign store_prevUnrecoded_rawIn_out_sig_lo=store_prevRecoded[22:0]; 
  assign store_prevUnrecoded_rawIn__sig={1'h0,store_prevUnrecoded_rawIn_out_sig_hi_lo,store_prevUnrecoded_rawIn_out_sig_lo}; 
  assign store_prevUnrecoded_isSubnormal=$signed(store_prevUnrecoded_rawIn__sExp)<10'sh82; 
  assign store_prevUnrecoded_denormShiftDist=5'h1-store_prevUnrecoded_rawIn__sExp[4:0]; 
  assign _store_prevUnrecoded_denormFract_T_1=store_prevUnrecoded_rawIn__sig[24:1]>>store_prevUnrecoded_denormShiftDist; 
  assign store_prevUnrecoded_denormFract=_store_prevUnrecoded_denormFract_T_1[22:0]; 
  assign _store_prevUnrecoded_expOut_T_2=store_prevUnrecoded_rawIn__sExp[7:0]-8'h81; 
  assign _store_prevUnrecoded_expOut_T_3=store_prevUnrecoded_isSubnormal ? 8'h0:_store_prevUnrecoded_expOut_T_2; 
  assign _store_prevUnrecoded_expOut_T_4=store_prevUnrecoded_rawIn__isNaN|store_prevUnrecoded_rawIn__isInf; 
  assign _store_prevUnrecoded_expOut_T_6=_store_prevUnrecoded_expOut_T_4 ? 8'hff:8'h0; 
  assign store_prevUnrecoded_hi_lo=_store_prevUnrecoded_expOut_T_3|_store_prevUnrecoded_expOut_T_6; 
  assign _store_prevUnrecoded_fractOut_T_1=store_prevUnrecoded_rawIn__isInf ? 23'h0:store_prevUnrecoded_rawIn__sig[22:0]; 
  assign store_prevUnrecoded_lo=store_prevUnrecoded_isSubnormal ? store_prevUnrecoded_denormFract:_store_prevUnrecoded_fractOut_T_1; 
  assign store_prevUnrecoded={store_prevUnrecoded_rawIn__sign,store_prevUnrecoded_hi_lo,store_prevUnrecoded_lo}; 
  assign store_hi=store_unrecoded[63:32]; 
  assign _store_T_1=&in_in1[63:61]; 
  assign store_lo=_store_T_1 ? store_prevUnrecoded:store_unrecoded[31:0]; 
  assign _store_T_3={store_hi,store_lo}; 
  assign store_hi_1=_store_T_3[31:0]; 
  assign _store_T_4={store_hi_1,store_hi_1}; 
  assign store_truncIdx=in_typeTagOut[0]; 
  assign store=store_truncIdx ? _store_T_3:_store_T_4; 
  assign intType_x6=in_fmt[0]; 
  assign cvtType=in_typ[1]; 
  assign io_out_bits_exc_hi_hi_1=conv_io_intExceptionFlags[2]|narrow_io_intExceptionFlags[1]; 
  assign toint_hi=conv_io_out[63:32]; 
  assign excSign=store_unrecoded_rawIn__sign&~_store_T_1; 
  assign excOut_hi=conv_io_signedOut==excSign; 
  assign excOut_lo=excSign ? 31'h0:31'h7fffffff; 
  assign _toint_T_10={toint_hi,excOut_hi,excOut_lo}; 
  assign _GEN_25=io_out_bits_exc_hi_hi_1 ? _toint_T_10:conv_io_out; 
  assign _GEN_26=cvtType ? conv_io_out:_GEN_25; 
  assign _toint_T_4={dcmp_io_lt,dcmp_io_eq}; 
  assign _GEN_34={1'b0,_toint_T_4}; 
  assign _toint_T_5=~in_rm&_GEN_34; 
  assign _toint_T_6=|_toint_T_5; 
  assign _toint_T_8={store[63:32],32'h0}; 
  assign _GEN_35={63'b0,_toint_T_6}; 
  assign _toint_T_9=_GEN_35|_toint_T_8; 
  assign _GEN_29=in_ren2 ? _toint_T_9:_GEN_26; 
  assign classify_out_hi_hi_hi_hi_1=_store_T_1&in_in1[51]; 
  assign classify_out_hi_hi_hi_lo_1=_store_T_1&~in_in1[51]; 
  assign classify_out_codeHi_1=in_in1[63:62]; 
  assign classify_out_isSpecial_1=classify_out_codeHi_1==2'h3; 
  assign classify_out_isInf_1=classify_out_isSpecial_1&~in_in1[61]; 
  assign classify_out_hi_hi_lo_1=classify_out_isInf_1&~store_unrecoded_rawIn__sign; 
  assign _classify_out_isNormal_T_4=classify_out_codeHi_1==2'h1; 
  assign classify_out_isHighSubnormalIn_1=in_in1[61:52]<10'h2; 
  assign _classify_out_isNormal_T_6=_classify_out_isNormal_T_4&~classify_out_isHighSubnormalIn_1; 
  assign _classify_out_isNormal_T_7=classify_out_codeHi_1==2'h2; 
  assign classify_out_isNormal_1=_classify_out_isNormal_T_6|_classify_out_isNormal_T_7; 
  assign classify_out_hi_lo_hi_1=classify_out_isNormal_1&~store_unrecoded_rawIn__sign; 
  assign _classify_out_isSubnormal_T_3=in_in1[63:61]==3'h1; 
  assign _classify_out_isSubnormal_T_5=_classify_out_isNormal_T_4&classify_out_isHighSubnormalIn_1; 
  assign classify_out_isSubnormal_1=_classify_out_isSubnormal_T_3|_classify_out_isSubnormal_T_5; 
  assign classify_out_hi_lo_lo_1=classify_out_isSubnormal_1&~store_unrecoded_rawIn__sign; 
  assign classify_out_isZero_1=in_in1[63:61]==3'h0; 
  assign classify_out_lo_hi_hi_hi_1=classify_out_isZero_1&~store_unrecoded_rawIn__sign; 
  assign classify_out_lo_hi_hi_lo_1=classify_out_isZero_1&store_unrecoded_rawIn__sign; 
  assign classify_out_lo_hi_lo_1=classify_out_isSubnormal_1&store_unrecoded_rawIn__sign; 
  assign classify_out_lo_lo_hi_1=classify_out_isNormal_1&store_unrecoded_rawIn__sign; 
  assign classify_out_lo_lo_lo_1=classify_out_isInf_1&store_unrecoded_rawIn__sign; 
  assign _classify_out_T_10={classify_out_hi_hi_hi_hi_1,classify_out_hi_hi_hi_lo_1,classify_out_hi_hi_lo_1,classify_out_hi_lo_hi_1,classify_out_hi_lo_lo_1,classify_out_lo_hi_hi_hi_1,classify_out_lo_hi_hi_lo_1,classify_out_lo_hi_lo_1,classify_out_lo_lo_hi_1,classify_out_lo_lo_lo_1}; 
  assign _classify_out_expOut_T_1=store_unrecoded_rawIn_exp[11:9]>=3'h6; 
  assign _classify_out_expOut_T_2=store_unrecoded_rawIn_isZero|_classify_out_expOut_T_1; 
  assign _classify_out_expOut_commonCase_T_1=store_unrecoded_rawIn_exp+12'h100; 
  assign classify_out_expOut_commonCase=_classify_out_expOut_commonCase_T_1-12'h800; 
  assign classify_out_expOut_lo=classify_out_expOut_commonCase[5:0]; 
  assign _classify_out_expOut_T_3={store_unrecoded_rawIn_exp[11:9],classify_out_expOut_lo}; 
  assign classify_out_hi_lo=_classify_out_expOut_T_2 ? _classify_out_expOut_T_3:classify_out_expOut_commonCase[8:0]; 
  assign _classify_out_fractOut_T={store_unrecoded_rawIn_out_sig_lo,24'h0}; 
  assign classify_out_lo=_classify_out_fractOut_T[75:53]; 
  assign _classify_out_T={store_unrecoded_rawIn__sign,classify_out_hi_lo,classify_out_lo}; 
  assign classify_out_code=_classify_out_T[31:29]; 
  assign classify_out_isNaN=&classify_out_code; 
  assign classify_out_hi_hi_hi_hi=classify_out_isNaN&_classify_out_T[22]; 
  assign classify_out_hi_hi_hi_lo=classify_out_isNaN&~_classify_out_T[22]; 
  assign classify_out_codeHi=classify_out_code[2:1]; 
  assign classify_out_isSpecial=classify_out_codeHi==2'h3; 
  assign classify_out_isInf=classify_out_isSpecial&~classify_out_code[0]; 
  assign classify_out_sign=_classify_out_T[32]; 
  assign classify_out_hi_hi_lo=classify_out_isInf&~classify_out_sign; 
  assign _classify_out_isNormal_T=classify_out_codeHi==2'h1; 
  assign classify_out_isHighSubnormalIn=_classify_out_T[29:23]<7'h2; 
  assign _classify_out_isNormal_T_2=_classify_out_isNormal_T&~classify_out_isHighSubnormalIn; 
  assign _classify_out_isNormal_T_3=classify_out_codeHi==2'h2; 
  assign classify_out_isNormal=_classify_out_isNormal_T_2|_classify_out_isNormal_T_3; 
  assign classify_out_hi_lo_hi=classify_out_isNormal&~classify_out_sign; 
  assign _classify_out_isSubnormal_T=classify_out_code==3'h1; 
  assign _classify_out_isSubnormal_T_2=_classify_out_isNormal_T&classify_out_isHighSubnormalIn; 
  assign classify_out_isSubnormal=_classify_out_isSubnormal_T|_classify_out_isSubnormal_T_2; 
  assign classify_out_hi_lo_lo=classify_out_isSubnormal&~classify_out_sign; 
  assign classify_out_isZero=classify_out_code==3'h0; 
  assign classify_out_lo_hi_hi_hi=classify_out_isZero&~classify_out_sign; 
  assign classify_out_lo_hi_hi_lo=classify_out_isZero&classify_out_sign; 
  assign classify_out_lo_hi_lo=classify_out_isSubnormal&classify_out_sign; 
  assign classify_out_lo_lo_hi=classify_out_isNormal&classify_out_sign; 
  assign classify_out_lo_lo_lo=classify_out_isInf&classify_out_sign; 
  assign _classify_out_T_5={classify_out_hi_hi_hi_hi,classify_out_hi_hi_hi_lo,classify_out_hi_hi_lo,classify_out_hi_lo_hi,classify_out_hi_lo_lo,classify_out_lo_hi_hi_hi,classify_out_lo_hi_hi_lo,classify_out_lo_hi_lo,classify_out_lo_lo_hi,classify_out_lo_lo_lo}; 
  assign classify_out=store_truncIdx ? _classify_out_T_10:_classify_out_T_5; 
  assign _GEN_36={54'b0,classify_out}; 
  assign _toint_T_2=_GEN_36|_toint_T_8; 
  assign _GEN_23=in_rm[0] ? _toint_T_2:store; 
  assign toint=in_wflags ? _GEN_29:_GEN_23; 
  assign io_out_bits_toint_lo=toint[31:0]; 
  assign io_out_bits_toint_hi=io_out_bits_toint_lo[31] ? 32'hffffffff:32'h0; 
  assign _io_out_bits_toint_T_2={io_out_bits_toint_hi,io_out_bits_toint_lo}; 
  assign _GEN_28=~in_ren2&cvtType; 
  assign _GEN_24=in_rm[0] ? 1'h0:intType_x6; 
  assign intType=in_wflags ? _GEN_28:_GEN_24; 
  assign io_out_bits_exc_hi_hi=|conv_io_intExceptionFlags[2:1]; 
  assign io_out_bits_exc_lo=conv_io_intExceptionFlags[0]; 
  assign _io_out_bits_exc_T_1={io_out_bits_exc_hi_hi,3'h0,io_out_bits_exc_lo}; 
  assign io_out_bits_exc_lo_1=~io_out_bits_exc_hi_hi_1&io_out_bits_exc_lo; 
  assign _io_out_bits_exc_T_4={io_out_bits_exc_hi_hi_1,3'h0,io_out_bits_exc_lo_1}; 
  assign _GEN_27=cvtType ? _io_out_bits_exc_T_1:_io_out_bits_exc_T_4; 
  assign _GEN_30=in_ren2 ? dcmp_io_exceptionFlags:_GEN_27; 
  assign _io_out_bits_lt_T_1=$signed(dcmp_io_a)<65'sh0; 
  assign _io_out_bits_lt_T_3=$signed(dcmp_io_b)>=65'sh0; 
  assign _io_out_bits_lt_T_4=_io_out_bits_lt_T_1&_io_out_bits_lt_T_3; 
  assign io_out_bits_in_rm=in_rm; 
  assign io_out_bits_in_in1=in_in1; 
  assign io_out_bits_in_in2=in_in2; 
  assign io_out_bits_lt=dcmp_io_lt|_io_out_bits_lt_T_4; 
  assign io_out_bits_store=store_truncIdx ? _store_T_3:_store_T_4; 
  assign io_out_bits_toint=intType ? toint:_io_out_bits_toint_T_2; 
  assign io_out_bits_exc=in_wflags ? _GEN_30:5'h0; 
  assign dcmp_io_a=in_in1; 
  assign dcmp_io_b=in_in2; 
  assign dcmp_io_signaling=~in_rm[1]; 
  assign conv_io_in=in_in1; 
  assign conv_io_roundingMode=in_rm; 
  assign conv_io_signedOut=~in_typ[0]; 
  assign narrow_io_in=in_in1; 
  assign narrow_io_roundingMode=in_rm; 
  assign narrow_io_signedOut=~in_typ[0]; 
  assign FPToInt_cov_read_addr=FPToInt_state; 
  assign FPToInt_cov_read_data=FPToInt_cov[FPToInt_cov_read_addr]; 
  assign FPToInt_cov_write_data=1'h1; 
  assign FPToInt_cov_write_addr=FPToInt_state; 
  assign FPToInt_cov_write_mask=1'h1; 
  assign FPToInt_cov_write_en=1'h1; 
  assign in_wflags_shl=in_wflags; 
  assign in_wflags_pad={3'h0,in_wflags_shl}; 
  assign in_typ_shl={in_typ,1'h0}; 
  assign in_typ_pad={1'h0,in_typ_shl}; 
  assign in_ren2_shl={in_ren2,3'h0}; 
  assign in_ren2_pad=in_ren2_shl; 
  assign FPToInt_xor2=in_typ_pad^in_ren2_pad; 
  assign FPToInt_xor0=in_wflags_pad^FPToInt_xor2; 
  assign dcmp_sum=FPToInt_covSum+dcmp_io_covSum; 
  assign conv_sum=dcmp_sum+conv_io_covSum; 
  assign narrow_sum=conv_sum+narrow_io_covSum; 
  assign io_covSum=narrow_sum; 
  assign dcmp_metaAssert_wire=dcmp_metaAssert; 
  assign conv_metaAssert_wire=conv_metaAssert; 
  assign narrow_metaAssert_wire=narrow_metaAssert; 
  assign FPToInt_or2=conv_metaAssert_wire|narrow_metaAssert_wire; 
  assign FPToInt_or0=dcmp_metaAssert_wire|FPToInt_or2; 
  assign metaAssert=FPToInt_or0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              in_ren2 <=1'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_ren2 <=io_in_bits_ren2;
               end 
         if (metaReset)
            begin 
              in_typeTagOut <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_typeTagOut <=io_in_bits_typeTagOut;
               end 
         if (metaReset)
            begin 
              in_wflags <=1'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_wflags <=io_in_bits_wflags;
               end 
         if (metaReset)
            begin 
              in_rm <=3'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_rm <=io_in_bits_rm;
               end 
         if (metaReset)
            begin 
              in_typ <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_typ <=io_in_bits_typ;
               end 
         if (metaReset)
            begin 
              in_fmt <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_fmt <=io_in_bits_fmt;
               end 
         if (metaReset)
            begin 
              in_in1 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_in1 <=io_in_bits_in1;
               end 
         if (metaReset)
            begin 
              in_in2 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_in2 <=io_in_bits_in2;
               end 
         FPToInt_state <=FPToInt_xor0;
         if (!(FPToInt_cov_read_data))
            begin 
              FPToInt_covSum <=FPToInt_covSum+1'h1;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (FPToInt_cov_write_en&FPToInt_cov_write_mask)
            begin 
              FPToInt_cov [FPToInt_cov_write_addr]<=FPToInt_cov_write_data;
            end 
       end
  
endmodule
 
module IntToFP (
  input clock,
  input reset,
  input io_in_valid,
  input [1:0] io_in_bits_typeTagIn,
  input io_in_bits_wflags,
  input [2:0] io_in_bits_rm,
  input [1:0] io_in_bits_typ,
  input [63:0] io_in_bits_in1,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire i2f_io_signedIn ;  
   wire [63:0] i2f_io_in ;  
   wire [2:0] i2f_io_roundingMode ;  
   wire [32:0] i2f_io_out ;  
   wire [4:0] i2f_io_exceptionFlags ;  
   wire [29:0] i2f_io_covSum ;  
   wire i2f_metaAssert ;  
   wire i2f_1_io_signedIn ;  
   wire [63:0] i2f_1_io_in ;  
   wire [2:0] i2f_1_io_roundingMode ;  
   wire [64:0] i2f_1_io_out ;  
   wire [4:0] i2f_1_io_exceptionFlags ;  
   wire [29:0] i2f_1_io_covSum ;  
   wire i2f_1_metaAssert ;  
   reg inPipe_valid ;  
   reg [31:0] _RAND_0 ;  
   reg [1:0] inPipe_bits_typeTagIn ;  
   reg [31:0] _RAND_1 ;  
   reg inPipe_bits_wflags ;  
   reg [31:0] _RAND_2 ;  
   reg [2:0] inPipe_bits_rm ;  
   reg [31:0] _RAND_3 ;  
   reg [1:0] inPipe_bits_typ ;  
   reg [31:0] _RAND_4 ;  
   reg [63:0] inPipe_bits_in1 ;  
   reg [63:0] _RAND_5 ;  
   wire mux_data_truncIdx ;  
   wire [63:0] _mux_data_T_1 ;  
   wire [63:0] _mux_data_T_2 ;  
   wire mux_data_rawIn_sign ;  
   wire [10:0] mux_data_rawIn_expIn ;  
   wire [51:0] mux_data_rawIn_fractIn ;  
   wire mux_data_rawIn_isZeroExpIn ;  
   wire mux_data_rawIn_isZeroFractIn ;  
   wire [5:0] _mux_data_rawIn_normDist_T_52 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_53 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_54 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_55 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_56 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_57 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_58 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_59 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_60 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_61 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_62 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_63 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_64 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_65 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_66 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_67 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_68 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_69 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_70 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_71 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_72 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_73 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_74 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_75 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_76 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_77 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_78 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_79 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_80 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_81 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_82 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_83 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_84 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_85 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_86 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_87 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_88 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_89 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_90 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_91 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_92 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_93 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_94 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_95 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_96 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_97 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_98 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_99 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_100 ;  
   wire [5:0] _mux_data_rawIn_normDist_T_101 ;  
   wire [5:0] mux_data_rawIn_normDist ;  
   wire [114:0] _GEN_24 ;  
   wire [114:0] _mux_data_rawIn_subnormFract_T ;  
   wire [51:0] mux_data_rawIn_subnormFract ;  
   wire [11:0] _GEN_25 ;  
   wire [11:0] _mux_data_rawIn_adjustedExp_T ;  
   wire [11:0] _mux_data_rawIn_adjustedExp_T_1 ;  
   wire [1:0] _mux_data_rawIn_adjustedExp_T_2 ;  
   wire [10:0] _GEN_26 ;  
   wire [10:0] _mux_data_rawIn_adjustedExp_T_3 ;  
   wire [11:0] _GEN_27 ;  
   wire [11:0] mux_data_rawIn_adjustedExp ;  
   wire mux_data_rawIn_isZero ;  
   wire mux_data_rawIn_isSpecial ;  
   wire mux_data_rawIn__isNaN ;  
   wire [12:0] mux_data_rawIn__sExp ;  
   wire mux_data_rawIn_out_sig_hi_lo ;  
   wire [51:0] mux_data_rawIn_out_sig_lo ;  
   wire [53:0] mux_data_rawIn__sig ;  
   wire [2:0] _mux_data_T_4 ;  
   wire [2:0] _GEN_28 ;  
   wire [2:0] mux_data_hi_lo ;  
   wire [8:0] mux_data_lo_hi ;  
   wire [51:0] mux_data_lo_lo ;  
   wire [64:0] _mux_data_T_6 ;  
   wire mux_data_rawIn_sign_1 ;  
   wire [7:0] mux_data_rawIn_expIn_1 ;  
   wire [22:0] mux_data_rawIn_fractIn_1 ;  
   wire mux_data_rawIn_isZeroExpIn_1 ;  
   wire mux_data_rawIn_isZeroFractIn_1 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_125 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_126 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_127 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_128 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_129 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_130 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_131 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_132 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_133 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_134 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_135 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_136 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_137 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_138 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_139 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_140 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_141 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_142 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_143 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_144 ;  
   wire [4:0] _mux_data_rawIn_normDist_T_145 ;  
   wire [4:0] mux_data_rawIn_normDist_1 ;  
   wire [53:0] _GEN_29 ;  
   wire [53:0] _mux_data_rawIn_subnormFract_T_2 ;  
   wire [22:0] mux_data_rawIn_subnormFract_1 ;  
   wire [8:0] _GEN_30 ;  
   wire [8:0] _mux_data_rawIn_adjustedExp_T_5 ;  
   wire [8:0] _mux_data_rawIn_adjustedExp_T_6 ;  
   wire [1:0] _mux_data_rawIn_adjustedExp_T_7 ;  
   wire [7:0] _GEN_31 ;  
   wire [7:0] _mux_data_rawIn_adjustedExp_T_8 ;  
   wire [8:0] _GEN_32 ;  
   wire [8:0] mux_data_rawIn_adjustedExp_1 ;  
   wire mux_data_rawIn_isZero_1 ;  
   wire mux_data_rawIn_isSpecial_1 ;  
   wire mux_data_rawIn_1_isNaN ;  
   wire [9:0] mux_data_rawIn_1_sExp ;  
   wire mux_data_rawIn_out_sig_hi_lo_1 ;  
   wire [22:0] mux_data_rawIn_out_sig_lo_1 ;  
   wire [24:0] mux_data_rawIn_1_sig ;  
   wire [2:0] _mux_data_T_8 ;  
   wire [2:0] _GEN_33 ;  
   wire [2:0] mux_data_hi_lo_1 ;  
   wire [5:0] mux_data_lo_hi_1 ;  
   wire [22:0] mux_data_lo_lo_1 ;  
   wire [32:0] _mux_data_T_10 ;  
   wire [3:0] mux_data_swizzledNaN_hi_hi_hi ;  
   wire mux_data_swizzledNaN_hi_hi_lo ;  
   wire [6:0] mux_data_swizzledNaN_hi_lo_hi ;  
   wire mux_data_swizzledNaN_hi_lo_lo ;  
   wire mux_data_swizzledNaN_lo_hi_lo ;  
   wire [30:0] mux_data_swizzledNaN_lo_lo ;  
   wire [64:0] mux_data_swizzledNaN ;  
   wire _mux_data_T_12 ;  
   wire [31:0] intValue_smallInt ;  
   wire [32:0] _intValue_res_T_1 ;  
   wire [31:0] _intValue_res_T_2 ;  
   wire [32:0] _intValue_res_T_3 ;  
   wire [64:0] maskedNaN ;  
   wire _T_1 ;  
   wire [64:0] _T_2 ;  
   wire [31:0] dataPadded_hi ;  
   wire [64:0] dataPadded_0 ;  
   reg [64:0] io_out_b_data ;  
   reg [95:0] _RAND_6 ;  
   reg [4:0] io_out_b_exc ;  
   reg [31:0] _RAND_7 ;  
   reg [3:0] IntToFP_state ;  
   reg [31:0] _RAND_8 ;  
   reg IntToFP_cov[0:15] ;  
   reg [31:0] _RAND_9 ;  
   wire IntToFP_cov_read_data ;  
   wire [3:0] IntToFP_cov_read_addr ;  
   wire IntToFP_cov_write_data ;  
   wire [3:0] IntToFP_cov_write_addr ;  
   wire IntToFP_cov_write_mask ;  
   wire IntToFP_cov_write_en ;  
   reg [29:0] IntToFP_covSum ;  
   reg [31:0] _RAND_10 ;  
   wire inPipe_valid_shl ;  
   wire [3:0] inPipe_valid_pad ;  
   wire [1:0] inPipe_bits_wflags_shl ;  
   wire [3:0] inPipe_bits_wflags_pad ;  
   wire [3:0] inPipe_bits_typ_shl ;  
   wire [3:0] inPipe_bits_typ_pad ;  
   wire [3:0] IntToFP_xor2 ;  
   wire [3:0] IntToFP_xor0 ;  
   wire [29:0] i2f_sum ;  
   wire [29:0] i2f_1_sum ;  
   wire i2f_metaAssert_wire ;  
   wire i2f_1_metaAssert_wire ;  
   wire IntToFP_or0 ;  
   reg IntToFP_metaAssert ;  
   reg [31:0] _RAND_11 ;  
  INToRecFN i2f(.io_signedIn(i2f_io_signedIn),.io_in(i2f_io_in),.io_roundingMode(i2f_io_roundingMode),.io_out(i2f_io_out),.io_exceptionFlags(i2f_io_exceptionFlags),.io_covSum(i2f_io_covSum),.metaAssert(i2f_metaAssert)); 
  INToRecFN_1 i2f_1(.io_signedIn(i2f_1_io_signedIn),.io_in(i2f_1_io_in),.io_roundingMode(i2f_1_io_roundingMode),.io_out(i2f_1_io_out),.io_exceptionFlags(i2f_1_io_exceptionFlags),.io_covSum(i2f_1_io_covSum),.metaAssert(i2f_1_metaAssert)); 
  assign mux_data_truncIdx=inPipe_bits_typeTagIn[0]; 
  assign _mux_data_T_1=mux_data_truncIdx ? 64'h0:64'hffffffff00000000; 
  assign _mux_data_T_2=_mux_data_T_1|inPipe_bits_in1; 
  assign mux_data_rawIn_sign=_mux_data_T_2[63]; 
  assign mux_data_rawIn_expIn=_mux_data_T_2[62:52]; 
  assign mux_data_rawIn_fractIn=_mux_data_T_2[51:0]; 
  assign mux_data_rawIn_isZeroExpIn=mux_data_rawIn_expIn==11'h0; 
  assign mux_data_rawIn_isZeroFractIn=mux_data_rawIn_fractIn==52'h0; 
  assign _mux_data_rawIn_normDist_T_52=mux_data_rawIn_fractIn[1] ? 6'h32:6'h33; 
  assign _mux_data_rawIn_normDist_T_53=mux_data_rawIn_fractIn[2] ? 6'h31:_mux_data_rawIn_normDist_T_52; 
  assign _mux_data_rawIn_normDist_T_54=mux_data_rawIn_fractIn[3] ? 6'h30:_mux_data_rawIn_normDist_T_53; 
  assign _mux_data_rawIn_normDist_T_55=mux_data_rawIn_fractIn[4] ? 6'h2f:_mux_data_rawIn_normDist_T_54; 
  assign _mux_data_rawIn_normDist_T_56=mux_data_rawIn_fractIn[5] ? 6'h2e:_mux_data_rawIn_normDist_T_55; 
  assign _mux_data_rawIn_normDist_T_57=mux_data_rawIn_fractIn[6] ? 6'h2d:_mux_data_rawIn_normDist_T_56; 
  assign _mux_data_rawIn_normDist_T_58=mux_data_rawIn_fractIn[7] ? 6'h2c:_mux_data_rawIn_normDist_T_57; 
  assign _mux_data_rawIn_normDist_T_59=mux_data_rawIn_fractIn[8] ? 6'h2b:_mux_data_rawIn_normDist_T_58; 
  assign _mux_data_rawIn_normDist_T_60=mux_data_rawIn_fractIn[9] ? 6'h2a:_mux_data_rawIn_normDist_T_59; 
  assign _mux_data_rawIn_normDist_T_61=mux_data_rawIn_fractIn[10] ? 6'h29:_mux_data_rawIn_normDist_T_60; 
  assign _mux_data_rawIn_normDist_T_62=mux_data_rawIn_fractIn[11] ? 6'h28:_mux_data_rawIn_normDist_T_61; 
  assign _mux_data_rawIn_normDist_T_63=mux_data_rawIn_fractIn[12] ? 6'h27:_mux_data_rawIn_normDist_T_62; 
  assign _mux_data_rawIn_normDist_T_64=mux_data_rawIn_fractIn[13] ? 6'h26:_mux_data_rawIn_normDist_T_63; 
  assign _mux_data_rawIn_normDist_T_65=mux_data_rawIn_fractIn[14] ? 6'h25:_mux_data_rawIn_normDist_T_64; 
  assign _mux_data_rawIn_normDist_T_66=mux_data_rawIn_fractIn[15] ? 6'h24:_mux_data_rawIn_normDist_T_65; 
  assign _mux_data_rawIn_normDist_T_67=mux_data_rawIn_fractIn[16] ? 6'h23:_mux_data_rawIn_normDist_T_66; 
  assign _mux_data_rawIn_normDist_T_68=mux_data_rawIn_fractIn[17] ? 6'h22:_mux_data_rawIn_normDist_T_67; 
  assign _mux_data_rawIn_normDist_T_69=mux_data_rawIn_fractIn[18] ? 6'h21:_mux_data_rawIn_normDist_T_68; 
  assign _mux_data_rawIn_normDist_T_70=mux_data_rawIn_fractIn[19] ? 6'h20:_mux_data_rawIn_normDist_T_69; 
  assign _mux_data_rawIn_normDist_T_71=mux_data_rawIn_fractIn[20] ? 6'h1f:_mux_data_rawIn_normDist_T_70; 
  assign _mux_data_rawIn_normDist_T_72=mux_data_rawIn_fractIn[21] ? 6'h1e:_mux_data_rawIn_normDist_T_71; 
  assign _mux_data_rawIn_normDist_T_73=mux_data_rawIn_fractIn[22] ? 6'h1d:_mux_data_rawIn_normDist_T_72; 
  assign _mux_data_rawIn_normDist_T_74=mux_data_rawIn_fractIn[23] ? 6'h1c:_mux_data_rawIn_normDist_T_73; 
  assign _mux_data_rawIn_normDist_T_75=mux_data_rawIn_fractIn[24] ? 6'h1b:_mux_data_rawIn_normDist_T_74; 
  assign _mux_data_rawIn_normDist_T_76=mux_data_rawIn_fractIn[25] ? 6'h1a:_mux_data_rawIn_normDist_T_75; 
  assign _mux_data_rawIn_normDist_T_77=mux_data_rawIn_fractIn[26] ? 6'h19:_mux_data_rawIn_normDist_T_76; 
  assign _mux_data_rawIn_normDist_T_78=mux_data_rawIn_fractIn[27] ? 6'h18:_mux_data_rawIn_normDist_T_77; 
  assign _mux_data_rawIn_normDist_T_79=mux_data_rawIn_fractIn[28] ? 6'h17:_mux_data_rawIn_normDist_T_78; 
  assign _mux_data_rawIn_normDist_T_80=mux_data_rawIn_fractIn[29] ? 6'h16:_mux_data_rawIn_normDist_T_79; 
  assign _mux_data_rawIn_normDist_T_81=mux_data_rawIn_fractIn[30] ? 6'h15:_mux_data_rawIn_normDist_T_80; 
  assign _mux_data_rawIn_normDist_T_82=mux_data_rawIn_fractIn[31] ? 6'h14:_mux_data_rawIn_normDist_T_81; 
  assign _mux_data_rawIn_normDist_T_83=mux_data_rawIn_fractIn[32] ? 6'h13:_mux_data_rawIn_normDist_T_82; 
  assign _mux_data_rawIn_normDist_T_84=mux_data_rawIn_fractIn[33] ? 6'h12:_mux_data_rawIn_normDist_T_83; 
  assign _mux_data_rawIn_normDist_T_85=mux_data_rawIn_fractIn[34] ? 6'h11:_mux_data_rawIn_normDist_T_84; 
  assign _mux_data_rawIn_normDist_T_86=mux_data_rawIn_fractIn[35] ? 6'h10:_mux_data_rawIn_normDist_T_85; 
  assign _mux_data_rawIn_normDist_T_87=mux_data_rawIn_fractIn[36] ? 6'hf:_mux_data_rawIn_normDist_T_86; 
  assign _mux_data_rawIn_normDist_T_88=mux_data_rawIn_fractIn[37] ? 6'he:_mux_data_rawIn_normDist_T_87; 
  assign _mux_data_rawIn_normDist_T_89=mux_data_rawIn_fractIn[38] ? 6'hd:_mux_data_rawIn_normDist_T_88; 
  assign _mux_data_rawIn_normDist_T_90=mux_data_rawIn_fractIn[39] ? 6'hc:_mux_data_rawIn_normDist_T_89; 
  assign _mux_data_rawIn_normDist_T_91=mux_data_rawIn_fractIn[40] ? 6'hb:_mux_data_rawIn_normDist_T_90; 
  assign _mux_data_rawIn_normDist_T_92=mux_data_rawIn_fractIn[41] ? 6'ha:_mux_data_rawIn_normDist_T_91; 
  assign _mux_data_rawIn_normDist_T_93=mux_data_rawIn_fractIn[42] ? 6'h9:_mux_data_rawIn_normDist_T_92; 
  assign _mux_data_rawIn_normDist_T_94=mux_data_rawIn_fractIn[43] ? 6'h8:_mux_data_rawIn_normDist_T_93; 
  assign _mux_data_rawIn_normDist_T_95=mux_data_rawIn_fractIn[44] ? 6'h7:_mux_data_rawIn_normDist_T_94; 
  assign _mux_data_rawIn_normDist_T_96=mux_data_rawIn_fractIn[45] ? 6'h6:_mux_data_rawIn_normDist_T_95; 
  assign _mux_data_rawIn_normDist_T_97=mux_data_rawIn_fractIn[46] ? 6'h5:_mux_data_rawIn_normDist_T_96; 
  assign _mux_data_rawIn_normDist_T_98=mux_data_rawIn_fractIn[47] ? 6'h4:_mux_data_rawIn_normDist_T_97; 
  assign _mux_data_rawIn_normDist_T_99=mux_data_rawIn_fractIn[48] ? 6'h3:_mux_data_rawIn_normDist_T_98; 
  assign _mux_data_rawIn_normDist_T_100=mux_data_rawIn_fractIn[49] ? 6'h2:_mux_data_rawIn_normDist_T_99; 
  assign _mux_data_rawIn_normDist_T_101=mux_data_rawIn_fractIn[50] ? 6'h1:_mux_data_rawIn_normDist_T_100; 
  assign mux_data_rawIn_normDist=mux_data_rawIn_fractIn[51] ? 6'h0:_mux_data_rawIn_normDist_T_101; 
  assign _GEN_24={63'b0,mux_data_rawIn_fractIn}; 
  assign _mux_data_rawIn_subnormFract_T=_GEN_24<<mux_data_rawIn_normDist; 
  assign mux_data_rawIn_subnormFract={_mux_data_rawIn_subnormFract_T[50:0],1'h0}; 
  assign _GEN_25={6'b0,mux_data_rawIn_normDist}; 
  assign _mux_data_rawIn_adjustedExp_T=_GEN_25^12'hfff; 
  assign _mux_data_rawIn_adjustedExp_T_1=mux_data_rawIn_isZeroExpIn ? _mux_data_rawIn_adjustedExp_T:{1'b0,mux_data_rawIn_expIn}; 
  assign _mux_data_rawIn_adjustedExp_T_2=mux_data_rawIn_isZeroExpIn ? 2'h2:2'h1; 
  assign _GEN_26={9'b0,_mux_data_rawIn_adjustedExp_T_2}; 
  assign _mux_data_rawIn_adjustedExp_T_3=11'h400|_GEN_26; 
  assign _GEN_27={1'b0,_mux_data_rawIn_adjustedExp_T_3}; 
  assign mux_data_rawIn_adjustedExp=_mux_data_rawIn_adjustedExp_T_1+_GEN_27; 
  assign mux_data_rawIn_isZero=mux_data_rawIn_isZeroExpIn&mux_data_rawIn_isZeroFractIn; 
  assign mux_data_rawIn_isSpecial=mux_data_rawIn_adjustedExp[11:10]==2'h3; 
  assign mux_data_rawIn__isNaN=mux_data_rawIn_isSpecial&~mux_data_rawIn_isZeroFractIn; 
  assign mux_data_rawIn__sExp={1'b0,$signed(mux_data_rawIn_adjustedExp)}; 
  assign mux_data_rawIn_out_sig_hi_lo=~mux_data_rawIn_isZero; 
  assign mux_data_rawIn_out_sig_lo=mux_data_rawIn_isZeroExpIn ? mux_data_rawIn_subnormFract:mux_data_rawIn_fractIn; 
  assign mux_data_rawIn__sig={1'h0,mux_data_rawIn_out_sig_hi_lo,mux_data_rawIn_out_sig_lo}; 
  assign _mux_data_T_4=mux_data_rawIn_isZero ? 3'h0:mux_data_rawIn__sExp[11:9]; 
  assign _GEN_28={2'b0,mux_data_rawIn__isNaN}; 
  assign mux_data_hi_lo=_mux_data_T_4|_GEN_28; 
  assign mux_data_lo_hi=mux_data_rawIn__sExp[8:0]; 
  assign mux_data_lo_lo=mux_data_rawIn__sig[51:0]; 
  assign _mux_data_T_6={mux_data_rawIn_sign,mux_data_hi_lo,mux_data_lo_hi,mux_data_lo_lo}; 
  assign mux_data_rawIn_sign_1=_mux_data_T_2[31]; 
  assign mux_data_rawIn_expIn_1=_mux_data_T_2[30:23]; 
  assign mux_data_rawIn_fractIn_1=_mux_data_T_2[22:0]; 
  assign mux_data_rawIn_isZeroExpIn_1=mux_data_rawIn_expIn_1==8'h0; 
  assign mux_data_rawIn_isZeroFractIn_1=mux_data_rawIn_fractIn_1==23'h0; 
  assign _mux_data_rawIn_normDist_T_125=mux_data_rawIn_fractIn_1[1] ? 5'h15:5'h16; 
  assign _mux_data_rawIn_normDist_T_126=mux_data_rawIn_fractIn_1[2] ? 5'h14:_mux_data_rawIn_normDist_T_125; 
  assign _mux_data_rawIn_normDist_T_127=mux_data_rawIn_fractIn_1[3] ? 5'h13:_mux_data_rawIn_normDist_T_126; 
  assign _mux_data_rawIn_normDist_T_128=mux_data_rawIn_fractIn_1[4] ? 5'h12:_mux_data_rawIn_normDist_T_127; 
  assign _mux_data_rawIn_normDist_T_129=mux_data_rawIn_fractIn_1[5] ? 5'h11:_mux_data_rawIn_normDist_T_128; 
  assign _mux_data_rawIn_normDist_T_130=mux_data_rawIn_fractIn_1[6] ? 5'h10:_mux_data_rawIn_normDist_T_129; 
  assign _mux_data_rawIn_normDist_T_131=mux_data_rawIn_fractIn_1[7] ? 5'hf:_mux_data_rawIn_normDist_T_130; 
  assign _mux_data_rawIn_normDist_T_132=mux_data_rawIn_fractIn_1[8] ? 5'he:_mux_data_rawIn_normDist_T_131; 
  assign _mux_data_rawIn_normDist_T_133=mux_data_rawIn_fractIn_1[9] ? 5'hd:_mux_data_rawIn_normDist_T_132; 
  assign _mux_data_rawIn_normDist_T_134=mux_data_rawIn_fractIn_1[10] ? 5'hc:_mux_data_rawIn_normDist_T_133; 
  assign _mux_data_rawIn_normDist_T_135=mux_data_rawIn_fractIn_1[11] ? 5'hb:_mux_data_rawIn_normDist_T_134; 
  assign _mux_data_rawIn_normDist_T_136=mux_data_rawIn_fractIn_1[12] ? 5'ha:_mux_data_rawIn_normDist_T_135; 
  assign _mux_data_rawIn_normDist_T_137=mux_data_rawIn_fractIn_1[13] ? 5'h9:_mux_data_rawIn_normDist_T_136; 
  assign _mux_data_rawIn_normDist_T_138=mux_data_rawIn_fractIn_1[14] ? 5'h8:_mux_data_rawIn_normDist_T_137; 
  assign _mux_data_rawIn_normDist_T_139=mux_data_rawIn_fractIn_1[15] ? 5'h7:_mux_data_rawIn_normDist_T_138; 
  assign _mux_data_rawIn_normDist_T_140=mux_data_rawIn_fractIn_1[16] ? 5'h6:_mux_data_rawIn_normDist_T_139; 
  assign _mux_data_rawIn_normDist_T_141=mux_data_rawIn_fractIn_1[17] ? 5'h5:_mux_data_rawIn_normDist_T_140; 
  assign _mux_data_rawIn_normDist_T_142=mux_data_rawIn_fractIn_1[18] ? 5'h4:_mux_data_rawIn_normDist_T_141; 
  assign _mux_data_rawIn_normDist_T_143=mux_data_rawIn_fractIn_1[19] ? 5'h3:_mux_data_rawIn_normDist_T_142; 
  assign _mux_data_rawIn_normDist_T_144=mux_data_rawIn_fractIn_1[20] ? 5'h2:_mux_data_rawIn_normDist_T_143; 
  assign _mux_data_rawIn_normDist_T_145=mux_data_rawIn_fractIn_1[21] ? 5'h1:_mux_data_rawIn_normDist_T_144; 
  assign mux_data_rawIn_normDist_1=mux_data_rawIn_fractIn_1[22] ? 5'h0:_mux_data_rawIn_normDist_T_145; 
  assign _GEN_29={31'b0,mux_data_rawIn_fractIn_1}; 
  assign _mux_data_rawIn_subnormFract_T_2=_GEN_29<<mux_data_rawIn_normDist_1; 
  assign mux_data_rawIn_subnormFract_1={_mux_data_rawIn_subnormFract_T_2[21:0],1'h0}; 
  assign _GEN_30={4'b0,mux_data_rawIn_normDist_1}; 
  assign _mux_data_rawIn_adjustedExp_T_5=_GEN_30^9'h1ff; 
  assign _mux_data_rawIn_adjustedExp_T_6=mux_data_rawIn_isZeroExpIn_1 ? _mux_data_rawIn_adjustedExp_T_5:{1'b0,mux_data_rawIn_expIn_1}; 
  assign _mux_data_rawIn_adjustedExp_T_7=mux_data_rawIn_isZeroExpIn_1 ? 2'h2:2'h1; 
  assign _GEN_31={6'b0,_mux_data_rawIn_adjustedExp_T_7}; 
  assign _mux_data_rawIn_adjustedExp_T_8=8'h80|_GEN_31; 
  assign _GEN_32={1'b0,_mux_data_rawIn_adjustedExp_T_8}; 
  assign mux_data_rawIn_adjustedExp_1=_mux_data_rawIn_adjustedExp_T_6+_GEN_32; 
  assign mux_data_rawIn_isZero_1=mux_data_rawIn_isZeroExpIn_1&mux_data_rawIn_isZeroFractIn_1; 
  assign mux_data_rawIn_isSpecial_1=mux_data_rawIn_adjustedExp_1[8:7]==2'h3; 
  assign mux_data_rawIn_1_isNaN=mux_data_rawIn_isSpecial_1&~mux_data_rawIn_isZeroFractIn_1; 
  assign mux_data_rawIn_1_sExp={1'b0,$signed(mux_data_rawIn_adjustedExp_1)}; 
  assign mux_data_rawIn_out_sig_hi_lo_1=~mux_data_rawIn_isZero_1; 
  assign mux_data_rawIn_out_sig_lo_1=mux_data_rawIn_isZeroExpIn_1 ? mux_data_rawIn_subnormFract_1:mux_data_rawIn_fractIn_1; 
  assign mux_data_rawIn_1_sig={1'h0,mux_data_rawIn_out_sig_hi_lo_1,mux_data_rawIn_out_sig_lo_1}; 
  assign _mux_data_T_8=mux_data_rawIn_isZero_1 ? 3'h0:mux_data_rawIn_1_sExp[8:6]; 
  assign _GEN_33={2'b0,mux_data_rawIn_1_isNaN}; 
  assign mux_data_hi_lo_1=_mux_data_T_8|_GEN_33; 
  assign mux_data_lo_hi_1=mux_data_rawIn_1_sExp[5:0]; 
  assign mux_data_lo_lo_1=mux_data_rawIn_1_sig[22:0]; 
  assign _mux_data_T_10={mux_data_rawIn_sign_1,mux_data_hi_lo_1,mux_data_lo_hi_1,mux_data_lo_lo_1}; 
  assign mux_data_swizzledNaN_hi_hi_hi=_mux_data_T_6[64:61]; 
  assign mux_data_swizzledNaN_hi_hi_lo=&_mux_data_T_6[51:32]; 
  assign mux_data_swizzledNaN_hi_lo_hi=_mux_data_T_6[59:53]; 
  assign mux_data_swizzledNaN_hi_lo_lo=_mux_data_T_10[31]; 
  assign mux_data_swizzledNaN_lo_hi_lo=_mux_data_T_10[32]; 
  assign mux_data_swizzledNaN_lo_lo=_mux_data_T_10[30:0]; 
  assign mux_data_swizzledNaN={mux_data_swizzledNaN_hi_hi_hi,mux_data_swizzledNaN_hi_hi_lo,mux_data_swizzledNaN_hi_lo_hi,mux_data_swizzledNaN_hi_lo_lo,_mux_data_T_6[51:32],mux_data_swizzledNaN_lo_hi_lo,mux_data_swizzledNaN_lo_lo}; 
  assign _mux_data_T_12=&_mux_data_T_6[63:61]; 
  assign intValue_smallInt=inPipe_bits_in1[31:0]; 
  assign _intValue_res_T_1={1'b0,$signed(intValue_smallInt)}; 
  assign _intValue_res_T_2=inPipe_bits_in1[31:0]; 
  assign _intValue_res_T_3=inPipe_bits_typ[0] ? $signed(_intValue_res_T_1):$signed({{1{_intValue_res_T_2[31]}},_intValue_res_T_2}); 
  assign maskedNaN=i2f_1_io_out&65'h1efefffffffffffff; 
  assign _T_1=&i2f_1_io_out[63:61]; 
  assign _T_2=_T_1 ? maskedNaN:i2f_1_io_out; 
  assign dataPadded_hi=_T_2[64:33]; 
  assign dataPadded_0={dataPadded_hi,i2f_io_out}; 
  assign io_out_bits_data=io_out_b_data; 
  assign io_out_bits_exc=io_out_b_exc; 
  assign i2f_io_signedIn=~inPipe_bits_typ[0]; 
  assign i2f_io_in=inPipe_bits_typ[1] ? $signed(inPipe_bits_in1):$signed({{31{_intValue_res_T_3[32]}},_intValue_res_T_3}); 
  assign i2f_io_roundingMode=inPipe_bits_rm; 
  assign i2f_1_io_signedIn=~inPipe_bits_typ[0]; 
  assign i2f_1_io_in=inPipe_bits_typ[1] ? $signed(inPipe_bits_in1):$signed({{31{_intValue_res_T_3[32]}},_intValue_res_T_3}); 
  assign i2f_1_io_roundingMode=inPipe_bits_rm; 
  assign IntToFP_cov_read_addr=IntToFP_state; 
  assign IntToFP_cov_read_data=IntToFP_cov[IntToFP_cov_read_addr]; 
  assign IntToFP_cov_write_data=1'h1; 
  assign IntToFP_cov_write_addr=IntToFP_state; 
  assign IntToFP_cov_write_mask=1'h1; 
  assign IntToFP_cov_write_en=1'h1; 
  assign inPipe_valid_shl=inPipe_valid; 
  assign inPipe_valid_pad={3'h0,inPipe_valid_shl}; 
  assign inPipe_bits_wflags_shl={inPipe_bits_wflags,1'h0}; 
  assign inPipe_bits_wflags_pad={2'h0,inPipe_bits_wflags_shl}; 
  assign inPipe_bits_typ_shl={inPipe_bits_typ,2'h0}; 
  assign inPipe_bits_typ_pad=inPipe_bits_typ_shl; 
  assign IntToFP_xor2=inPipe_bits_wflags_pad^inPipe_bits_typ_pad; 
  assign IntToFP_xor0=inPipe_valid_pad^IntToFP_xor2; 
  assign i2f_sum=IntToFP_covSum+i2f_io_covSum; 
  assign i2f_1_sum=i2f_sum+i2f_1_io_covSum; 
  assign io_covSum=i2f_1_sum; 
  assign i2f_metaAssert_wire=i2f_metaAssert; 
  assign i2f_1_metaAssert_wire=i2f_1_metaAssert; 
  assign IntToFP_or0=i2f_metaAssert_wire|i2f_1_metaAssert_wire; 
  assign metaAssert=IntToFP_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              inPipe_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 inPipe_valid <=1'h0;
               end 
             else 
               begin 
                 inPipe_valid <=io_in_valid;
               end 
         if (metaReset)
            begin 
              inPipe_bits_typeTagIn <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_typeTagIn <=io_in_bits_typeTagIn;
               end 
         if (metaReset)
            begin 
              inPipe_bits_wflags <=1'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_wflags <=io_in_bits_wflags;
               end 
         if (metaReset)
            begin 
              inPipe_bits_rm <=3'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_rm <=io_in_bits_rm;
               end 
         if (metaReset)
            begin 
              inPipe_bits_typ <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_typ <=io_in_bits_typ;
               end 
         if (metaReset)
            begin 
              inPipe_bits_in1 <=64'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_in1 <=io_in_bits_in1;
               end 
         if (metaReset)
            begin 
              io_out_b_data <=65'h0;
            end 
          else 
            if (inPipe_valid)
               begin 
                 if (inPipe_bits_wflags)
                    begin 
                      if (mux_data_truncIdx)
                         begin 
                           if (_T_1)
                              begin 
                                io_out_b_data <=maskedNaN;
                              end 
                            else 
                              begin 
                                io_out_b_data <=i2f_1_io_out;
                              end 
                         end 
                       else 
                         begin 
                           io_out_b_data <=dataPadded_0;
                         end 
                    end 
                  else 
                    if (_mux_data_T_12)
                       begin 
                         io_out_b_data <=mux_data_swizzledNaN;
                       end 
                     else 
                       begin 
                         io_out_b_data <=_mux_data_T_6;
                       end 
               end 
         if (metaReset)
            begin 
              io_out_b_exc <=5'h0;
            end 
          else 
            if (inPipe_valid)
               begin 
                 if (inPipe_bits_wflags)
                    begin 
                      if (mux_data_truncIdx)
                         begin 
                           io_out_b_exc <=i2f_1_io_exceptionFlags;
                         end 
                       else 
                         begin 
                           io_out_b_exc <=i2f_io_exceptionFlags;
                         end 
                    end 
                  else 
                    begin 
                      io_out_b_exc <=5'h0;
                    end 
               end 
         IntToFP_state <=IntToFP_xor0;
         if (!(IntToFP_cov_read_data))
            begin 
              IntToFP_covSum <=IntToFP_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              IntToFP_metaAssert <=1'h0;
            end 
          else 
            begin 
              IntToFP_metaAssert <=IntToFP_metaAssert|IntToFP_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (IntToFP_cov_write_en&IntToFP_cov_write_mask)
            begin 
              IntToFP_cov [IntToFP_cov_write_addr]<=IntToFP_cov_write_data;
            end 
       end
  
endmodule
 
module FPToFP (
  input clock,
  input reset,
  input io_in_valid,
  input io_in_bits_ren2,
  input [1:0] io_in_bits_typeTagOut,
  input io_in_bits_wflags,
  input [2:0] io_in_bits_rm,
  input [64:0] io_in_bits_in1,
  input [64:0] io_in_bits_in2,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc,
  input io_lt,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [64:0] narrower_io_in ;  
   wire [2:0] narrower_io_roundingMode ;  
   wire [32:0] narrower_io_out ;  
   wire [4:0] narrower_io_exceptionFlags ;  
   wire [29:0] narrower_io_covSum ;  
   wire narrower_metaAssert ;  
   reg inPipe_valid ;  
   reg [31:0] _RAND_0 ;  
   reg inPipe_bits_ren2 ;  
   reg [31:0] _RAND_1 ;  
   reg [1:0] inPipe_bits_typeTagOut ;  
   reg [31:0] _RAND_2 ;  
   reg inPipe_bits_wflags ;  
   reg [31:0] _RAND_3 ;  
   reg [2:0] inPipe_bits_rm ;  
   reg [31:0] _RAND_4 ;  
   reg [64:0] inPipe_bits_in1 ;  
   reg [95:0] _RAND_5 ;  
   reg [64:0] inPipe_bits_in2 ;  
   reg [95:0] _RAND_6 ;  
   wire [64:0] _signNum_T_1 ;  
   wire [64:0] _signNum_T_4 ;  
   wire [64:0] signNum ;  
   wire fsgnj_hi ;  
   wire [63:0] fsgnj_lo ;  
   wire [64:0] fsgnj ;  
   wire isnan1 ;  
   wire isnan2 ;  
   wire _isInvalid_T_4 ;  
   wire _isInvalid_T_9 ;  
   wire isInvalid ;  
   wire isNaNOut ;  
   wire _isLHS_T_1 ;  
   wire _isLHS_T_3 ;  
   wire isLHS ;  
   wire [4:0] _fsgnjMux_exc_T ;  
   wire [64:0] _fsgnjMux_data_T ;  
   wire [64:0] _fsgnjMux_data_T_1 ;  
   wire [64:0] _GEN_24 ;  
   wire _T ;  
   wire _T_2 ;  
   wire [64:0] widened ;  
   wire [64:0] fsgnjMux_data ;  
   wire [31:0] mux_data_hi ;  
   wire mux_data_hi_hi ;  
   wire [51:0] mux_data_fractIn ;  
   wire [11:0] mux_data_expIn ;  
   wire [75:0] _mux_data_fractOut_T ;  
   wire [22:0] mux_data_lo ;  
   wire [2:0] mux_data_expOut_hi ;  
   wire [11:0] _mux_data_expOut_commonCase_T_1 ;  
   wire [11:0] mux_data_expOut_commonCase ;  
   wire _mux_data_expOut_T ;  
   wire _mux_data_expOut_T_1 ;  
   wire _mux_data_expOut_T_2 ;  
   wire [5:0] mux_data_expOut_lo ;  
   wire [8:0] _mux_data_expOut_T_3 ;  
   wire [8:0] mux_data_hi_lo ;  
   wire [64:0] _mux_data_T ;  
   wire [4:0] _fsgnjMux_exc_T_6 ;  
   wire [64:0] _mux_data_T_1 ;  
   reg [64:0] io_out_b_data ;  
   reg [95:0] _RAND_7 ;  
   reg [4:0] io_out_b_exc ;  
   reg [31:0] _RAND_8 ;  
   reg [5:0] FPToFP_state ;  
   reg [31:0] _RAND_9 ;  
   reg FPToFP_cov[0:63] ;  
   reg [31:0] _RAND_10 ;  
   wire FPToFP_cov_read_data ;  
   wire [5:0] FPToFP_cov_read_addr ;  
   wire FPToFP_cov_write_data ;  
   wire [5:0] FPToFP_cov_write_addr ;  
   wire FPToFP_cov_write_mask ;  
   wire FPToFP_cov_write_en ;  
   reg [29:0] FPToFP_covSum ;  
   reg [31:0] _RAND_11 ;  
   wire inPipe_valid_shl ;  
   wire [5:0] inPipe_valid_pad ;  
   wire [1:0] inPipe_bits_ren2_shl ;  
   wire [5:0] inPipe_bits_ren2_pad ;  
   wire [2:0] inPipe_bits_wflags_shl ;  
   wire [5:0] inPipe_bits_wflags_pad ;  
   wire [5:0] inPipe_bits_rm_shl ;  
   wire [5:0] inPipe_bits_rm_pad ;  
   wire [5:0] FPToFP_xor1 ;  
   wire [5:0] FPToFP_xor2 ;  
   wire [5:0] FPToFP_xor0 ;  
   wire [29:0] narrower_sum ;  
   wire narrower_metaAssert_wire ;  
   reg FPToFP_metaAssert ;  
   reg [31:0] _RAND_12 ;  
  RecFNToRecFN narrower(.io_in(narrower_io_in),.io_roundingMode(narrower_io_roundingMode),.io_out(narrower_io_out),.io_exceptionFlags(narrower_io_exceptionFlags),.io_covSum(narrower_io_covSum),.metaAssert(narrower_metaAssert)); 
  assign _signNum_T_1=inPipe_bits_in1^inPipe_bits_in2; 
  assign _signNum_T_4=inPipe_bits_rm[0] ? ~inPipe_bits_in2:inPipe_bits_in2; 
  assign signNum=inPipe_bits_rm[1] ? _signNum_T_1:_signNum_T_4; 
  assign fsgnj_hi=signNum[64]; 
  assign fsgnj_lo=inPipe_bits_in1[63:0]; 
  assign fsgnj={fsgnj_hi,fsgnj_lo}; 
  assign isnan1=&inPipe_bits_in1[63:61]; 
  assign isnan2=&inPipe_bits_in2[63:61]; 
  assign _isInvalid_T_4=isnan1&~inPipe_bits_in1[51]; 
  assign _isInvalid_T_9=isnan2&~inPipe_bits_in2[51]; 
  assign isInvalid=_isInvalid_T_4|_isInvalid_T_9; 
  assign isNaNOut=isnan1&isnan2; 
  assign _isLHS_T_1=inPipe_bits_rm[0]!=io_lt; 
  assign _isLHS_T_3=_isLHS_T_1&~isnan1; 
  assign isLHS=isnan2|_isLHS_T_3; 
  assign _fsgnjMux_exc_T={isInvalid,4'h0}; 
  assign _fsgnjMux_data_T=isLHS ? inPipe_bits_in1:inPipe_bits_in2; 
  assign _fsgnjMux_data_T_1=isNaNOut ? 65'he008000000000000:_fsgnjMux_data_T; 
  assign _GEN_24=inPipe_bits_wflags ? _fsgnjMux_data_T_1:fsgnj; 
  assign _T=inPipe_bits_typeTagOut==2'h0; 
  assign _T_2=inPipe_bits_wflags&~inPipe_bits_ren2; 
  assign widened=isnan1 ? 65'he008000000000000:inPipe_bits_in1; 
  assign fsgnjMux_data=_T_2 ? widened:_GEN_24; 
  assign mux_data_hi=fsgnjMux_data[64:33]; 
  assign mux_data_hi_hi=fsgnjMux_data[64]; 
  assign mux_data_fractIn=fsgnjMux_data[51:0]; 
  assign mux_data_expIn=fsgnjMux_data[63:52]; 
  assign _mux_data_fractOut_T={mux_data_fractIn,24'h0}; 
  assign mux_data_lo=_mux_data_fractOut_T[75:53]; 
  assign mux_data_expOut_hi=mux_data_expIn[11:9]; 
  assign _mux_data_expOut_commonCase_T_1=mux_data_expIn+12'h100; 
  assign mux_data_expOut_commonCase=_mux_data_expOut_commonCase_T_1-12'h800; 
  assign _mux_data_expOut_T=mux_data_expOut_hi==3'h0; 
  assign _mux_data_expOut_T_1=mux_data_expOut_hi>=3'h6; 
  assign _mux_data_expOut_T_2=_mux_data_expOut_T|_mux_data_expOut_T_1; 
  assign mux_data_expOut_lo=mux_data_expOut_commonCase[5:0]; 
  assign _mux_data_expOut_T_3={mux_data_expOut_hi,mux_data_expOut_lo}; 
  assign mux_data_hi_lo=_mux_data_expOut_T_2 ? _mux_data_expOut_T_3:mux_data_expOut_commonCase[8:0]; 
  assign _mux_data_T={mux_data_hi,mux_data_hi_hi,mux_data_hi_lo,mux_data_lo}; 
  assign _fsgnjMux_exc_T_6={_isInvalid_T_4,4'h0}; 
  assign _mux_data_T_1={mux_data_hi,narrower_io_out}; 
  assign io_out_bits_data=io_out_b_data; 
  assign io_out_bits_exc=io_out_b_exc; 
  assign narrower_io_in=inPipe_bits_in1; 
  assign narrower_io_roundingMode=inPipe_bits_rm; 
  assign FPToFP_cov_read_addr=FPToFP_state; 
  assign FPToFP_cov_read_data=FPToFP_cov[FPToFP_cov_read_addr]; 
  assign FPToFP_cov_write_data=1'h1; 
  assign FPToFP_cov_write_addr=FPToFP_state; 
  assign FPToFP_cov_write_mask=1'h1; 
  assign FPToFP_cov_write_en=1'h1; 
  assign inPipe_valid_shl=inPipe_valid; 
  assign inPipe_valid_pad={5'h0,inPipe_valid_shl}; 
  assign inPipe_bits_ren2_shl={inPipe_bits_ren2,1'h0}; 
  assign inPipe_bits_ren2_pad={4'h0,inPipe_bits_ren2_shl}; 
  assign inPipe_bits_wflags_shl={inPipe_bits_wflags,2'h0}; 
  assign inPipe_bits_wflags_pad={3'h0,inPipe_bits_wflags_shl}; 
  assign inPipe_bits_rm_shl={inPipe_bits_rm,3'h0}; 
  assign inPipe_bits_rm_pad=inPipe_bits_rm_shl; 
  assign FPToFP_xor1=inPipe_valid_pad^inPipe_bits_ren2_pad; 
  assign FPToFP_xor2=inPipe_bits_wflags_pad^inPipe_bits_rm_pad; 
  assign FPToFP_xor0=FPToFP_xor1^FPToFP_xor2; 
  assign narrower_sum=FPToFP_covSum+narrower_io_covSum; 
  assign io_covSum=narrower_sum; 
  assign narrower_metaAssert_wire=narrower_metaAssert; 
  assign metaAssert=FPToFP_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              inPipe_valid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 inPipe_valid <=1'h0;
               end 
             else 
               begin 
                 inPipe_valid <=io_in_valid;
               end 
         if (metaReset)
            begin 
              inPipe_bits_ren2 <=1'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_ren2 <=io_in_bits_ren2;
               end 
         if (metaReset)
            begin 
              inPipe_bits_typeTagOut <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_typeTagOut <=io_in_bits_typeTagOut;
               end 
         if (metaReset)
            begin 
              inPipe_bits_wflags <=1'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_wflags <=io_in_bits_wflags;
               end 
         if (metaReset)
            begin 
              inPipe_bits_rm <=3'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_rm <=io_in_bits_rm;
               end 
         if (metaReset)
            begin 
              inPipe_bits_in1 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_in1 <=io_in_bits_in1;
               end 
         if (metaReset)
            begin 
              inPipe_bits_in2 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 inPipe_bits_in2 <=io_in_bits_in2;
               end 
         if (metaReset)
            begin 
              io_out_b_data <=65'h0;
            end 
          else 
            if (inPipe_valid)
               begin 
                 if (_T_2)
                    begin 
                      if (_T)
                         begin 
                           io_out_b_data <=_mux_data_T_1;
                         end 
                       else 
                         if (_T)
                            begin 
                              io_out_b_data <=_mux_data_T;
                            end 
                          else 
                            if (_T_2)
                               begin 
                                 if (isnan1)
                                    begin 
                                      io_out_b_data <=65'he008000000000000;
                                    end 
                                  else 
                                    begin 
                                      io_out_b_data <=inPipe_bits_in1;
                                    end 
                               end 
                             else 
                               if (inPipe_bits_wflags)
                                  begin 
                                    if (isNaNOut)
                                       begin 
                                         io_out_b_data <=65'he008000000000000;
                                       end 
                                     else 
                                       if (isLHS)
                                          begin 
                                            io_out_b_data <=inPipe_bits_in1;
                                          end 
                                        else 
                                          begin 
                                            io_out_b_data <=inPipe_bits_in2;
                                          end 
                                  end 
                                else 
                                  begin 
                                    io_out_b_data <=fsgnj;
                                  end 
                    end 
                  else 
                    if (_T)
                       begin 
                         io_out_b_data <=_mux_data_T;
                       end 
                     else 
                       if (_T_2)
                          begin 
                            if (isnan1)
                               begin 
                                 io_out_b_data <=65'he008000000000000;
                               end 
                             else 
                               begin 
                                 io_out_b_data <=inPipe_bits_in1;
                               end 
                          end 
                        else 
                          if (inPipe_bits_wflags)
                             begin 
                               if (isNaNOut)
                                  begin 
                                    io_out_b_data <=65'he008000000000000;
                                  end 
                                else 
                                  if (isLHS)
                                     begin 
                                       io_out_b_data <=inPipe_bits_in1;
                                     end 
                                   else 
                                     begin 
                                       io_out_b_data <=inPipe_bits_in2;
                                     end 
                             end 
                           else 
                             begin 
                               io_out_b_data <=fsgnj;
                             end 
               end 
         if (metaReset)
            begin 
              io_out_b_exc <=5'h0;
            end 
          else 
            if (inPipe_valid)
               begin 
                 if (_T_2)
                    begin 
                      if (_T)
                         begin 
                           io_out_b_exc <=narrower_io_exceptionFlags;
                         end 
                       else 
                         if (_T_2)
                            begin 
                              io_out_b_exc <=_fsgnjMux_exc_T_6;
                            end 
                          else 
                            if (inPipe_bits_wflags)
                               begin 
                                 io_out_b_exc <=_fsgnjMux_exc_T;
                               end 
                             else 
                               begin 
                                 io_out_b_exc <=5'h0;
                               end 
                    end 
                  else 
                    if (_T_2)
                       begin 
                         io_out_b_exc <=_fsgnjMux_exc_T_6;
                       end 
                     else 
                       if (inPipe_bits_wflags)
                          begin 
                            io_out_b_exc <=_fsgnjMux_exc_T;
                          end 
                        else 
                          begin 
                            io_out_b_exc <=5'h0;
                          end 
               end 
         FPToFP_state <=FPToFP_xor0;
         if (!(FPToFP_cov_read_data))
            begin 
              FPToFP_covSum <=FPToFP_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              FPToFP_metaAssert <=1'h0;
            end 
          else 
            begin 
              FPToFP_metaAssert <=FPToFP_metaAssert|narrower_metaAssert_wire;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (FPToFP_cov_write_en&FPToFP_cov_write_mask)
            begin 
              FPToFP_cov [FPToFP_cov_write_addr]<=FPToFP_cov_write_data;
            end 
       end
  
endmodule
 
module FPUFMAPipe_1 (
  input clock,
  input reset,
  input io_in_valid,
  input io_in_bits_ren3,
  input io_in_bits_swap23,
  input [2:0] io_in_bits_rm,
  input [1:0] io_in_bits_fmaCmd,
  input [64:0] io_in_bits_in1,
  input [64:0] io_in_bits_in2,
  input [64:0] io_in_bits_in3,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input fma_halt) ; 
   wire fma_clock ;  
   wire fma_reset ;  
   wire fma_io_validin ;  
   wire [1:0] fma_io_op ;  
   wire [64:0] fma_io_a ;  
   wire [64:0] fma_io_b ;  
   wire [64:0] fma_io_c ;  
   wire [2:0] fma_io_roundingMode ;  
   wire [64:0] fma_io_out ;  
   wire [4:0] fma_io_exceptionFlags ;  
   wire fma_io_validout ;  
   wire [29:0] fma_io_covSum ;  
   wire fma_metaAssert ;  
   wire fma_metaReset ;  
   reg valid ;  
   reg [31:0] _RAND_0 ;  
   reg [2:0] in_rm ;  
   reg [31:0] _RAND_1 ;  
   reg [1:0] in_fmaCmd ;  
   reg [31:0] _RAND_2 ;  
   reg [64:0] in_in1 ;  
   reg [95:0] _RAND_3 ;  
   reg [64:0] in_in2 ;  
   reg [95:0] _RAND_4 ;  
   reg [64:0] in_in3 ;  
   reg [95:0] _RAND_5 ;  
   wire [64:0] _zero_T ;  
   wire [64:0] zero ;  
   wire _T ;  
   wire [64:0] res_data_maskedNaN ;  
   wire _res_data_T_1 ;  
   reg [64:0] io_out_b_data ;  
   reg [95:0] _RAND_6 ;  
   reg [4:0] io_out_b_exc ;  
   reg [31:0] _RAND_7 ;  
   wire [4:0] res_exc ;  
   wire [29:0] FPUFMAPipe_1_covSum ;  
   wire [29:0] fma_sum ;  
   wire fma_metaAssert_wire ;  
   reg FPUFMAPipe_1_metaAssert ;  
   reg [31:0] _RAND_8 ;  
  MulAddRecFNPipe_1 fma(.clock(fma_clock),.reset(fma_reset),.io_validin(fma_io_validin),.io_op(fma_io_op),.io_a(fma_io_a),.io_b(fma_io_b),.io_c(fma_io_c),.io_roundingMode(fma_io_roundingMode),.io_out(fma_io_out),.io_exceptionFlags(fma_io_exceptionFlags),.io_validout(fma_io_validout),.io_covSum(fma_io_covSum),.metaAssert(fma_metaAssert),.metaReset(fma_metaReset)); 
  assign _zero_T=io_in_bits_in1^io_in_bits_in2; 
  assign zero=_zero_T&65'h10000000000000000; 
  assign _T=io_in_bits_ren3|io_in_bits_swap23; 
  assign res_data_maskedNaN=fma_io_out&65'h1efefffffffffffff; 
  assign _res_data_T_1=&fma_io_out[63:61]; 
  assign res_exc=fma_io_exceptionFlags; 
  assign io_out_bits_data=io_out_b_data; 
  assign io_out_bits_exc=io_out_b_exc; 
  assign fma_clock=clock; 
  assign fma_reset=reset; 
  assign fma_io_validin=valid; 
  assign fma_io_op=in_fmaCmd; 
  assign fma_io_a=in_in1; 
  assign fma_io_b=in_in2; 
  assign fma_io_c=in_in3; 
  assign fma_io_roundingMode=in_rm; 
  assign FPUFMAPipe_1_covSum=30'h0; 
  assign fma_sum=FPUFMAPipe_1_covSum+fma_io_covSum; 
  assign io_covSum=fma_sum; 
  assign fma_metaAssert_wire=fma_metaAssert; 
  assign metaAssert=FPUFMAPipe_1_metaAssert; 
  assign fma_metaReset=metaReset|fma_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              valid <=1'h0;
            end 
          else 
            begin 
              valid <=io_in_valid;
            end 
         if (metaReset)
            begin 
              in_rm <=3'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_rm <=io_in_bits_rm;
               end 
         if (metaReset)
            begin 
              in_fmaCmd <=2'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_fmaCmd <=io_in_bits_fmaCmd;
               end 
         if (metaReset)
            begin 
              in_in1 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 in_in1 <=io_in_bits_in1;
               end 
         if (metaReset)
            begin 
              in_in2 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 if (io_in_bits_swap23)
                    begin 
                      in_in2 <=65'h8000000000000000;
                    end 
                  else 
                    begin 
                      in_in2 <=io_in_bits_in2;
                    end 
               end 
         if (metaReset)
            begin 
              in_in3 <=65'h0;
            end 
          else 
            if (io_in_valid)
               begin 
                 if (~_T)
                    begin 
                      in_in3 <=zero;
                    end 
                  else 
                    begin 
                      in_in3 <=io_in_bits_in3;
                    end 
               end 
         if (metaReset)
            begin 
              io_out_b_data <=65'h0;
            end 
          else 
            if (fma_io_validout)
               begin 
                 if (_res_data_T_1)
                    begin 
                      io_out_b_data <=res_data_maskedNaN;
                    end 
                  else 
                    begin 
                      io_out_b_data <=fma_io_out;
                    end 
               end 
         if (metaReset)
            begin 
              io_out_b_exc <=5'h0;
            end 
          else 
            if (fma_io_validout)
               begin 
                 io_out_b_exc <=res_exc;
               end 
         if (metaReset)
            begin 
              FPUFMAPipe_1_metaAssert <=1'h0;
            end 
          else 
            begin 
              FPUFMAPipe_1_metaAssert <=FPUFMAPipe_1_metaAssert|fma_metaAssert_wire;
            end 
       end
  
endmodule
 
module DivSqrtRecFN_small (
  input clock,
  input reset,
  output io_inReady,
  input io_inValid,
  input io_sqrtOp,
  input [32:0] io_a,
  input [32:0] io_b,
  input [2:0] io_roundingMode,
  output io_outValid_div,
  output io_outValid_sqrt,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input divSqrtRecFNToRaw_halt) ; 
   wire divSqrtRecFNToRaw_clock ;  
   wire divSqrtRecFNToRaw_reset ;  
   wire divSqrtRecFNToRaw_io_inReady ;  
   wire divSqrtRecFNToRaw_io_inValid ;  
   wire divSqrtRecFNToRaw_io_sqrtOp ;  
   wire [32:0] divSqrtRecFNToRaw_io_a ;  
   wire [32:0] divSqrtRecFNToRaw_io_b ;  
   wire [2:0] divSqrtRecFNToRaw_io_roundingMode ;  
   wire divSqrtRecFNToRaw_io_rawOutValid_div ;  
   wire divSqrtRecFNToRaw_io_rawOutValid_sqrt ;  
   wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut ;  
   wire divSqrtRecFNToRaw_io_invalidExc ;  
   wire divSqrtRecFNToRaw_io_infiniteExc ;  
   wire divSqrtRecFNToRaw_io_rawOut_isNaN ;  
   wire divSqrtRecFNToRaw_io_rawOut_isInf ;  
   wire divSqrtRecFNToRaw_io_rawOut_isZero ;  
   wire divSqrtRecFNToRaw_io_rawOut_sign ;  
   wire [9:0] divSqrtRecFNToRaw_io_rawOut_sExp ;  
   wire [26:0] divSqrtRecFNToRaw_io_rawOut_sig ;  
   wire [29:0] divSqrtRecFNToRaw_io_covSum ;  
   wire divSqrtRecFNToRaw_metaAssert ;  
   wire divSqrtRecFNToRaw_metaReset ;  
   wire divSqrtRecFNToRaw_divSqrtRawFN__halt ;  
   wire roundRawFNToRecFN_io_invalidExc ;  
   wire roundRawFNToRecFN_io_infiniteExc ;  
   wire roundRawFNToRecFN_io_in_isNaN ;  
   wire roundRawFNToRecFN_io_in_isInf ;  
   wire roundRawFNToRecFN_io_in_isZero ;  
   wire roundRawFNToRecFN_io_in_sign ;  
   wire [9:0] roundRawFNToRecFN_io_in_sExp ;  
   wire [26:0] roundRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundRawFNToRecFN_io_roundingMode ;  
   wire roundRawFNToRecFN_io_detectTininess ;  
   wire [32:0] roundRawFNToRecFN_io_out ;  
   wire [4:0] roundRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundRawFNToRecFN_io_covSum ;  
   wire roundRawFNToRecFN_metaAssert ;  
   wire [29:0] DivSqrtRecFN_small_covSum ;  
   wire [29:0] divSqrtRecFNToRaw_sum ;  
   wire [29:0] roundRawFNToRecFN_sum ;  
   wire divSqrtRecFNToRaw_metaAssert_wire ;  
   wire roundRawFNToRecFN_metaAssert_wire ;  
   wire DivSqrtRecFN_small_or0 ;  
   reg DivSqrtRecFN_small_metaAssert ;  
   reg [31:0] _RAND_0 ;  
  DivSqrtRecFNToRaw_small divSqrtRecFNToRaw(.clock(divSqrtRecFNToRaw_clock),.reset(divSqrtRecFNToRaw_reset),.io_inReady(divSqrtRecFNToRaw_io_inReady),.io_inValid(divSqrtRecFNToRaw_io_inValid),.io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),.io_a(divSqrtRecFNToRaw_io_a),.io_b(divSqrtRecFNToRaw_io_b),.io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),.io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),.io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),.io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),.io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),.io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),.io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),.io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),.io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),.io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),.io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),.io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),.io_covSum(divSqrtRecFNToRaw_io_covSum),.metaAssert(divSqrtRecFNToRaw_metaAssert),.metaReset(divSqrtRecFNToRaw_metaReset),.divSqrtRawFN__halt(divSqrtRecFNToRaw_divSqrtRawFN__halt)); 
  RoundRawFNToRecFN_2 roundRawFNToRecFN(.io_invalidExc(roundRawFNToRecFN_io_invalidExc),.io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),.io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),.io_in_isInf(roundRawFNToRecFN_io_in_isInf),.io_in_isZero(roundRawFNToRecFN_io_in_isZero),.io_in_sign(roundRawFNToRecFN_io_in_sign),.io_in_sExp(roundRawFNToRecFN_io_in_sExp),.io_in_sig(roundRawFNToRecFN_io_in_sig),.io_roundingMode(roundRawFNToRecFN_io_roundingMode),.io_detectTininess(roundRawFNToRecFN_io_detectTininess),.io_out(roundRawFNToRecFN_io_out),.io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),.io_covSum(roundRawFNToRecFN_io_covSum),.metaAssert(roundRawFNToRecFN_metaAssert)); 
  assign io_inReady=divSqrtRecFNToRaw_io_inReady; 
  assign io_outValid_div=divSqrtRecFNToRaw_io_rawOutValid_div; 
  assign io_outValid_sqrt=divSqrtRecFNToRaw_io_rawOutValid_sqrt; 
  assign io_out=roundRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundRawFNToRecFN_io_exceptionFlags; 
  assign divSqrtRecFNToRaw_clock=clock; 
  assign divSqrtRecFNToRaw_reset=reset; 
  assign divSqrtRecFNToRaw_io_inValid=io_inValid; 
  assign divSqrtRecFNToRaw_io_sqrtOp=io_sqrtOp; 
  assign divSqrtRecFNToRaw_io_a=io_a; 
  assign divSqrtRecFNToRaw_io_b=io_b; 
  assign divSqrtRecFNToRaw_io_roundingMode=io_roundingMode; 
  assign roundRawFNToRecFN_io_invalidExc=divSqrtRecFNToRaw_io_invalidExc; 
  assign roundRawFNToRecFN_io_infiniteExc=divSqrtRecFNToRaw_io_infiniteExc; 
  assign roundRawFNToRecFN_io_in_isNaN=divSqrtRecFNToRaw_io_rawOut_isNaN; 
  assign roundRawFNToRecFN_io_in_isInf=divSqrtRecFNToRaw_io_rawOut_isInf; 
  assign roundRawFNToRecFN_io_in_isZero=divSqrtRecFNToRaw_io_rawOut_isZero; 
  assign roundRawFNToRecFN_io_in_sign=divSqrtRecFNToRaw_io_rawOut_sign; 
  assign roundRawFNToRecFN_io_in_sExp=divSqrtRecFNToRaw_io_rawOut_sExp; 
  assign roundRawFNToRecFN_io_in_sig=divSqrtRecFNToRaw_io_rawOut_sig; 
  assign roundRawFNToRecFN_io_roundingMode=divSqrtRecFNToRaw_io_roundingModeOut; 
  assign roundRawFNToRecFN_io_detectTininess=1'h1; 
  assign DivSqrtRecFN_small_covSum=30'h0; 
  assign divSqrtRecFNToRaw_sum=DivSqrtRecFN_small_covSum+divSqrtRecFNToRaw_io_covSum; 
  assign roundRawFNToRecFN_sum=divSqrtRecFNToRaw_sum+roundRawFNToRecFN_io_covSum; 
  assign io_covSum=roundRawFNToRecFN_sum; 
  assign divSqrtRecFNToRaw_metaAssert_wire=divSqrtRecFNToRaw_metaAssert; 
  assign roundRawFNToRecFN_metaAssert_wire=roundRawFNToRecFN_metaAssert; 
  assign DivSqrtRecFN_small_or0=divSqrtRecFNToRaw_metaAssert_wire|roundRawFNToRecFN_metaAssert_wire; 
  assign metaAssert=DivSqrtRecFN_small_metaAssert; 
  assign divSqrtRecFNToRaw_metaReset=metaReset|divSqrtRecFNToRaw_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              DivSqrtRecFN_small_metaAssert <=1'h0;
            end 
          else 
            begin 
              DivSqrtRecFN_small_metaAssert <=DivSqrtRecFN_small_metaAssert|DivSqrtRecFN_small_or0;
            end 
       end
  
endmodule
 
module DivSqrtRecFN_small_1 (
  input clock,
  input reset,
  output io_inReady,
  input io_inValid,
  input io_sqrtOp,
  input [64:0] io_a,
  input [64:0] io_b,
  input [2:0] io_roundingMode,
  output io_outValid_div,
  output io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input divSqrtRecFNToRaw_halt) ; 
   wire divSqrtRecFNToRaw_clock ;  
   wire divSqrtRecFNToRaw_reset ;  
   wire divSqrtRecFNToRaw_io_inReady ;  
   wire divSqrtRecFNToRaw_io_inValid ;  
   wire divSqrtRecFNToRaw_io_sqrtOp ;  
   wire [64:0] divSqrtRecFNToRaw_io_a ;  
   wire [64:0] divSqrtRecFNToRaw_io_b ;  
   wire [2:0] divSqrtRecFNToRaw_io_roundingMode ;  
   wire divSqrtRecFNToRaw_io_rawOutValid_div ;  
   wire divSqrtRecFNToRaw_io_rawOutValid_sqrt ;  
   wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut ;  
   wire divSqrtRecFNToRaw_io_invalidExc ;  
   wire divSqrtRecFNToRaw_io_infiniteExc ;  
   wire divSqrtRecFNToRaw_io_rawOut_isNaN ;  
   wire divSqrtRecFNToRaw_io_rawOut_isInf ;  
   wire divSqrtRecFNToRaw_io_rawOut_isZero ;  
   wire divSqrtRecFNToRaw_io_rawOut_sign ;  
   wire [12:0] divSqrtRecFNToRaw_io_rawOut_sExp ;  
   wire [55:0] divSqrtRecFNToRaw_io_rawOut_sig ;  
   wire [29:0] divSqrtRecFNToRaw_io_covSum ;  
   wire divSqrtRecFNToRaw_metaAssert ;  
   wire divSqrtRecFNToRaw_metaReset ;  
   wire divSqrtRecFNToRaw_divSqrtRawFN__halt ;  
   wire roundRawFNToRecFN_io_invalidExc ;  
   wire roundRawFNToRecFN_io_infiniteExc ;  
   wire roundRawFNToRecFN_io_in_isNaN ;  
   wire roundRawFNToRecFN_io_in_isInf ;  
   wire roundRawFNToRecFN_io_in_isZero ;  
   wire roundRawFNToRecFN_io_in_sign ;  
   wire [12:0] roundRawFNToRecFN_io_in_sExp ;  
   wire [55:0] roundRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundRawFNToRecFN_io_roundingMode ;  
   wire roundRawFNToRecFN_io_detectTininess ;  
   wire [64:0] roundRawFNToRecFN_io_out ;  
   wire [4:0] roundRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundRawFNToRecFN_io_covSum ;  
   wire roundRawFNToRecFN_metaAssert ;  
   wire [29:0] DivSqrtRecFN_small_1_covSum ;  
   wire [29:0] divSqrtRecFNToRaw_sum ;  
   wire [29:0] roundRawFNToRecFN_sum ;  
   wire divSqrtRecFNToRaw_metaAssert_wire ;  
   wire roundRawFNToRecFN_metaAssert_wire ;  
   wire DivSqrtRecFN_small_1_or0 ;  
   reg DivSqrtRecFN_small_1_metaAssert ;  
   reg [31:0] _RAND_0 ;  
  DivSqrtRecFNToRaw_small_1 divSqrtRecFNToRaw(.clock(divSqrtRecFNToRaw_clock),.reset(divSqrtRecFNToRaw_reset),.io_inReady(divSqrtRecFNToRaw_io_inReady),.io_inValid(divSqrtRecFNToRaw_io_inValid),.io_sqrtOp(divSqrtRecFNToRaw_io_sqrtOp),.io_a(divSqrtRecFNToRaw_io_a),.io_b(divSqrtRecFNToRaw_io_b),.io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),.io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),.io_rawOutValid_sqrt(divSqrtRecFNToRaw_io_rawOutValid_sqrt),.io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),.io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),.io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),.io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),.io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),.io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),.io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),.io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),.io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig),.io_covSum(divSqrtRecFNToRaw_io_covSum),.metaAssert(divSqrtRecFNToRaw_metaAssert),.metaReset(divSqrtRecFNToRaw_metaReset),.divSqrtRawFN__halt(divSqrtRecFNToRaw_divSqrtRawFN__halt)); 
  RoundRawFNToRecFN_3 roundRawFNToRecFN(.io_invalidExc(roundRawFNToRecFN_io_invalidExc),.io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),.io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),.io_in_isInf(roundRawFNToRecFN_io_in_isInf),.io_in_isZero(roundRawFNToRecFN_io_in_isZero),.io_in_sign(roundRawFNToRecFN_io_in_sign),.io_in_sExp(roundRawFNToRecFN_io_in_sExp),.io_in_sig(roundRawFNToRecFN_io_in_sig),.io_roundingMode(roundRawFNToRecFN_io_roundingMode),.io_detectTininess(roundRawFNToRecFN_io_detectTininess),.io_out(roundRawFNToRecFN_io_out),.io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),.io_covSum(roundRawFNToRecFN_io_covSum),.metaAssert(roundRawFNToRecFN_metaAssert)); 
  assign io_inReady=divSqrtRecFNToRaw_io_inReady; 
  assign io_outValid_div=divSqrtRecFNToRaw_io_rawOutValid_div; 
  assign io_outValid_sqrt=divSqrtRecFNToRaw_io_rawOutValid_sqrt; 
  assign io_out=roundRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundRawFNToRecFN_io_exceptionFlags; 
  assign divSqrtRecFNToRaw_clock=clock; 
  assign divSqrtRecFNToRaw_reset=reset; 
  assign divSqrtRecFNToRaw_io_inValid=io_inValid; 
  assign divSqrtRecFNToRaw_io_sqrtOp=io_sqrtOp; 
  assign divSqrtRecFNToRaw_io_a=io_a; 
  assign divSqrtRecFNToRaw_io_b=io_b; 
  assign divSqrtRecFNToRaw_io_roundingMode=io_roundingMode; 
  assign roundRawFNToRecFN_io_invalidExc=divSqrtRecFNToRaw_io_invalidExc; 
  assign roundRawFNToRecFN_io_infiniteExc=divSqrtRecFNToRaw_io_infiniteExc; 
  assign roundRawFNToRecFN_io_in_isNaN=divSqrtRecFNToRaw_io_rawOut_isNaN; 
  assign roundRawFNToRecFN_io_in_isInf=divSqrtRecFNToRaw_io_rawOut_isInf; 
  assign roundRawFNToRecFN_io_in_isZero=divSqrtRecFNToRaw_io_rawOut_isZero; 
  assign roundRawFNToRecFN_io_in_sign=divSqrtRecFNToRaw_io_rawOut_sign; 
  assign roundRawFNToRecFN_io_in_sExp=divSqrtRecFNToRaw_io_rawOut_sExp; 
  assign roundRawFNToRecFN_io_in_sig=divSqrtRecFNToRaw_io_rawOut_sig; 
  assign roundRawFNToRecFN_io_roundingMode=divSqrtRecFNToRaw_io_roundingModeOut; 
  assign roundRawFNToRecFN_io_detectTininess=1'h1; 
  assign DivSqrtRecFN_small_1_covSum=30'h0; 
  assign divSqrtRecFNToRaw_sum=DivSqrtRecFN_small_1_covSum+divSqrtRecFNToRaw_io_covSum; 
  assign roundRawFNToRecFN_sum=divSqrtRecFNToRaw_sum+roundRawFNToRecFN_io_covSum; 
  assign io_covSum=roundRawFNToRecFN_sum; 
  assign divSqrtRecFNToRaw_metaAssert_wire=divSqrtRecFNToRaw_metaAssert; 
  assign roundRawFNToRecFN_metaAssert_wire=roundRawFNToRecFN_metaAssert; 
  assign DivSqrtRecFN_small_1_or0=divSqrtRecFNToRaw_metaAssert_wire|roundRawFNToRecFN_metaAssert_wire; 
  assign metaAssert=DivSqrtRecFN_small_1_metaAssert; 
  assign divSqrtRecFNToRaw_metaReset=metaReset|divSqrtRecFNToRaw_halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              DivSqrtRecFN_small_1_metaAssert <=1'h0;
            end 
          else 
            begin 
              DivSqrtRecFN_small_1_metaAssert <=DivSqrtRecFN_small_1_metaAssert|DivSqrtRecFN_small_1_or0;
            end 
       end
  
endmodule
 
module Arbiter (
  output io_in_0_ready,
  input io_in_0_valid,
  input [26:0] io_in_0_bits_bits_addr,
  output io_in_1_ready,
  input io_in_1_valid,
  input io_in_1_bits_valid,
  input [26:0] io_in_1_bits_bits_addr,
  input io_out_ready,
  output io_out_valid,
  output io_out_bits_valid,
  output [26:0] io_out_bits_bits_addr,
  output io_chosen,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire grant_1 ;  
   wire [29:0] Arbiter_covSum ;  
  assign grant_1=~io_in_0_valid; 
  assign io_in_0_ready=io_out_ready; 
  assign io_in_1_ready=grant_1&io_out_ready; 
  assign io_out_valid=~grant_1|io_in_1_valid; 
  assign io_out_bits_valid=io_in_0_valid|io_in_1_bits_valid; 
  assign io_out_bits_bits_addr=io_in_0_valid ? io_in_0_bits_bits_addr:io_in_1_bits_bits_addr; 
  assign io_chosen=io_in_0_valid ? 1'h0:1'h1; 
  assign Arbiter_covSum=30'h0; 
  assign io_covSum=Arbiter_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module OptimizationBarrier_42 (
  input [2:0] io_x,
  output [2:0] io_y,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [29:0] OptimizationBarrier_42_covSum ;  
  assign io_y=io_x; 
  assign OptimizationBarrier_42_covSum=30'h0; 
  assign io_covSum=OptimizationBarrier_42_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module OptimizationBarrier_43 (
  input [53:0] io_x_ppn,
  input io_x_d,
  input io_x_a,
  input io_x_g,
  input io_x_u,
  input io_x_x,
  input io_x_w,
  input io_x_r,
  input io_x_v,
  output [53:0] io_y_ppn,
  output io_y_d,
  output io_y_a,
  output io_y_g,
  output io_y_u,
  output io_y_x,
  output io_y_w,
  output io_y_r,
  output io_y_v,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [29:0] OptimizationBarrier_43_covSum ;  
  assign io_y_ppn=io_x_ppn; 
  assign io_y_d=io_x_d; 
  assign io_y_a=io_x_a; 
  assign io_y_g=io_x_g; 
  assign io_y_u=io_x_u; 
  assign io_y_x=io_x_x; 
  assign io_y_w=io_x_w; 
  assign io_y_r=io_x_r; 
  assign io_y_v=io_x_v; 
  assign OptimizationBarrier_43_covSum=30'h0; 
  assign io_covSum=OptimizationBarrier_43_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module IBuf (
  input clock,
  input reset,
  output io_imem_ready,
  input io_imem_valid,
  input io_imem_bits_btb_taken,
  input io_imem_bits_btb_bridx,
  input [4:0] io_imem_bits_btb_entry,
  input [7:0] io_imem_bits_btb_bht_history,
  input [39:0] io_imem_bits_pc,
  input [31:0] io_imem_bits_data,
  input io_imem_bits_xcpt_pf_inst,
  input io_imem_bits_xcpt_ae_inst,
  input io_imem_bits_replay,
  input io_kill,
  output [39:0] io_pc,
  output [4:0] io_btb_resp_entry,
  output [7:0] io_btb_resp_bht_history,
  input io_inst_0_ready,
  output io_inst_0_valid,
  output io_inst_0_bits_xcpt0_pf_inst,
  output io_inst_0_bits_xcpt0_ae_inst,
  output io_inst_0_bits_xcpt1_pf_inst,
  output io_inst_0_bits_xcpt1_ae_inst,
  output io_inst_0_bits_replay,
  output io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0] io_inst_0_bits_inst_rd,
  output [4:0] io_inst_0_bits_inst_rs1,
  output [4:0] io_inst_0_bits_inst_rs2,
  output [4:0] io_inst_0_bits_inst_rs3,
  output [31:0] io_inst_0_bits_raw,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [31:0] exp_io_in ;  
   wire [31:0] exp_io_out_bits ;  
   wire [4:0] exp_io_out_rd ;  
   wire [4:0] exp_io_out_rs1 ;  
   wire [4:0] exp_io_out_rs2 ;  
   wire [4:0] exp_io_out_rs3 ;  
   wire exp_io_rvc ;  
   wire [29:0] exp_io_covSum ;  
   wire exp_metaAssert ;  
   reg nBufValid ;  
   reg [31:0] _RAND_0 ;  
   reg [39:0] buf__pc ;  
   reg [63:0] _RAND_1 ;  
   reg [31:0] buf__data ;  
   reg [31:0] _RAND_2 ;  
   reg buf__xcpt_pf_inst ;  
   reg [31:0] _RAND_3 ;  
   reg buf__xcpt_ae_inst ;  
   reg [31:0] _RAND_4 ;  
   reg buf__replay ;  
   reg [31:0] _RAND_5 ;  
   reg [4:0] ibufBTBResp_entry ;  
   reg [31:0] _RAND_6 ;  
   reg [7:0] ibufBTBResp_bht_history ;  
   reg [31:0] _RAND_7 ;  
   wire pcWordBits ;  
   wire [1:0] _nIC_T ;  
   wire [1:0] _nIC_T_1 ;  
   wire [1:0] _GEN_56 ;  
   wire [1:0] nIC ;  
   wire [1:0] _nValid_T ;  
   wire [1:0] _GEN_57 ;  
   wire [1:0] nValid ;  
   wire [3:0] _valid_T ;  
   wire [3:0] _valid_T_2 ;  
   wire [1:0] valid ;  
   wire [1:0] _full_insn_T_2 ;  
   wire _full_insn_T_4 ;  
   wire [1:0] _bufMask_T ;  
   wire [1:0] bufMask ;  
   wire [1:0] buf_replay ;  
   wire full_insn ;  
   wire [1:0] _nReady_T_4 ;  
   wire [1:0] nReady ;  
   wire [1:0] nICReady ;  
   wire _io_imem_ready_T ;  
   wire _io_imem_ready_T_1 ;  
   wire _io_imem_ready_T_2 ;  
   wire [1:0] _io_imem_ready_T_4 ;  
   wire _io_imem_ready_T_5 ;  
   wire _io_imem_ready_T_6 ;  
   wire _nBufValid_T_2 ;  
   wire [1:0] _nBufValid_T_4 ;  
   wire [1:0] _nBufValid_T_5 ;  
   wire _T_1 ;  
   wire _T_2 ;  
   wire _T_3 ;  
   wire _T_7 ;  
   wire [1:0] shamt ;  
   wire [15:0] buf_data_data_hi ;  
   wire [63:0] buf_data_data ;  
   wire [5:0] _buf_data_T ;  
   wire [63:0] _buf_data_T_1 ;  
   wire [39:0] _buf_pc_T_1 ;  
   wire [2:0] _buf_pc_T_2 ;  
   wire [39:0] _GEN_65 ;  
   wire [39:0] _buf_pc_T_4 ;  
   wire [39:0] _buf_pc_T_5 ;  
   wire [39:0] _buf_pc_T_6 ;  
   wire [1:0] _GEN_0 ;  
   wire [1:0] _GEN_23 ;  
   wire [1:0] _GEN_46 ;  
   wire [1:0] _icShiftAmt_T_1 ;  
   wire [1:0] icShiftAmt ;  
   wire [15:0] icData_hi ;  
   wire [63:0] icData_data_lo ;  
   wire [15:0] icData_data_hi ;  
   wire [127:0] icData_data ;  
   wire [5:0] _icData_T ;  
   wire [190:0] _GEN_68 ;  
   wire [190:0] _icData_T_1 ;  
   wire [31:0] icData ;  
   wire [4:0] _icMask_T_1 ;  
   wire [62:0] _icMask_T_2 ;  
   wire [31:0] icMask ;  
   wire [31:0] _inst_T ;  
   wire [31:0] _inst_T_2 ;  
   wire xcpt_1_pf_inst ;  
   wire xcpt_1_ae_inst ;  
   wire [1:0] _ic_replay_T_1 ;  
   wire [1:0] _ic_replay_T_2 ;  
   wire [1:0] ic_replay ;  
   wire _T_10 ;  
   wire _T_11 ;  
   wire _T_12 ;  
   wire _T_14 ;  
   wire _io_pc_T ;  
   wire [1:0] _replay_T_5 ;  
   wire _replay_T_7 ;  
   wire [1:0] _io_inst_0_bits_xcpt1_T_4 ;  
   wire [1:0] _io_inst_0_bits_xcpt1_T_5 ;  
   wire _T_18 ;  
   wire [1:0] _T_21 ;  
   wire _T_23 ;  
   reg [1:0] IBuf_state ;  
   reg [31:0] _RAND_8 ;  
   reg IBuf_cov[0:3] ;  
   reg [31:0] _RAND_9 ;  
   wire IBuf_cov_read_data ;  
   wire [1:0] IBuf_cov_read_addr ;  
   wire IBuf_cov_write_data ;  
   wire [1:0] IBuf_cov_write_addr ;  
   wire IBuf_cov_write_mask ;  
   wire IBuf_cov_write_en ;  
   reg [29:0] IBuf_covSum ;  
   reg [31:0] _RAND_10 ;  
   wire nBufValid_shl ;  
   wire [1:0] nBufValid_pad ;  
   wire [1:0] buf__replay_shl ;  
   wire [1:0] buf__replay_pad ;  
   wire [1:0] IBuf_xor0 ;  
   wire [29:0] exp_sum ;  
   wire stopEn0 ;  
   wire exp_metaAssert_wire ;  
   wire IBuf_or0 ;  
   reg IBuf_metaAssert ;  
   reg [31:0] _RAND_11 ;  
  RVCExpander exp(.io_in(exp_io_in),.io_out_bits(exp_io_out_bits),.io_out_rd(exp_io_out_rd),.io_out_rs1(exp_io_out_rs1),.io_out_rs2(exp_io_out_rs2),.io_out_rs3(exp_io_out_rs3),.io_rvc(exp_io_rvc),.io_covSum(exp_io_covSum),.metaAssert(exp_metaAssert)); 
  assign pcWordBits=io_imem_bits_pc[1]; 
  assign _nIC_T=io_imem_bits_btb_bridx+1'h1; 
  assign _nIC_T_1=io_imem_bits_btb_taken ? _nIC_T:2'h2; 
  assign _GEN_56={1'b0,pcWordBits}; 
  assign nIC=_nIC_T_1-_GEN_56; 
  assign _nValid_T=io_imem_valid ? nIC:2'h0; 
  assign _GEN_57={1'b0,nBufValid}; 
  assign nValid=_nValid_T+_GEN_57; 
  assign _valid_T=4'h1<<nValid; 
  assign _valid_T_2=_valid_T-4'h1; 
  assign valid=_valid_T_2[1:0]; 
  assign _full_insn_T_2={1'b0,valid[1]}; 
  assign _full_insn_T_4=exp_io_rvc|_full_insn_T_2[0]; 
  assign _bufMask_T=2'h1<<nBufValid; 
  assign bufMask=_bufMask_T-2'h1; 
  assign buf_replay=buf__replay ? bufMask:2'h0; 
  assign full_insn=_full_insn_T_4|buf_replay[0]; 
  assign _nReady_T_4=exp_io_rvc ? 2'h1:2'h2; 
  assign nReady=full_insn ? _nReady_T_4:2'h0; 
  assign nICReady=nReady-_GEN_57; 
  assign _io_imem_ready_T=nReady>=_GEN_57; 
  assign _io_imem_ready_T_1=io_inst_0_ready&_io_imem_ready_T; 
  assign _io_imem_ready_T_2=nICReady>=nIC; 
  assign _io_imem_ready_T_4=nIC-nICReady; 
  assign _io_imem_ready_T_5=2'h1>=_io_imem_ready_T_4; 
  assign _io_imem_ready_T_6=_io_imem_ready_T_2|_io_imem_ready_T_5; 
  assign _nBufValid_T_2=_io_imem_ready_T|~nBufValid; 
  assign _nBufValid_T_4=_GEN_57-nReady; 
  assign _nBufValid_T_5=_nBufValid_T_2 ? 2'h0:_nBufValid_T_4; 
  assign _T_1=io_imem_valid&_io_imem_ready_T; 
  assign _T_2=nICReady<nIC; 
  assign _T_3=_T_1&_T_2; 
  assign _T_7=_T_3&_io_imem_ready_T_5; 
  assign shamt=_GEN_56+nICReady; 
  assign buf_data_data_hi=io_imem_bits_data[31:16]; 
  assign buf_data_data={buf_data_data_hi,buf_data_data_hi,io_imem_bits_data}; 
  assign _buf_data_T={shamt,4'h0}; 
  assign _buf_data_T_1=buf_data_data>>_buf_data_T; 
  assign _buf_pc_T_1=io_imem_bits_pc&40'hfffffffffc; 
  assign _buf_pc_T_2={nICReady,1'h0}; 
  assign _GEN_65={37'b0,_buf_pc_T_2}; 
  assign _buf_pc_T_4=io_imem_bits_pc+_GEN_65; 
  assign _buf_pc_T_5=_buf_pc_T_4&40'h3; 
  assign _buf_pc_T_6=_buf_pc_T_1|_buf_pc_T_5; 
  assign _GEN_0=_T_7 ? _io_imem_ready_T_4:_nBufValid_T_5; 
  assign _GEN_23=io_inst_0_ready ? _GEN_0:{1'b0,nBufValid}; 
  assign _GEN_46=io_kill ? 2'h0:_GEN_23; 
  assign _icShiftAmt_T_1=2'h2+_GEN_57; 
  assign icShiftAmt=_icShiftAmt_T_1-_GEN_56; 
  assign icData_hi=io_imem_bits_data[15:0]; 
  assign icData_data_lo={io_imem_bits_data,icData_hi,icData_hi}; 
  assign icData_data_hi=icData_data_lo[63:48]; 
  assign icData_data={icData_data_hi,icData_data_hi,icData_data_hi,icData_data_hi,io_imem_bits_data,icData_hi,icData_hi}; 
  assign _icData_T={icShiftAmt,4'h0}; 
  assign _GEN_68={63'b0,icData_data}; 
  assign _icData_T_1=_GEN_68<<_icData_T; 
  assign icData=_icData_T_1[95:64]; 
  assign _icMask_T_1={nBufValid,4'h0}; 
  assign _icMask_T_2=63'hffffffff<<_icMask_T_1; 
  assign icMask=_icMask_T_2[31:0]; 
  assign _inst_T=icData&icMask; 
  assign _inst_T_2=buf__data&~icMask; 
  assign xcpt_1_pf_inst=bufMask[1] ? buf__xcpt_pf_inst:io_imem_bits_xcpt_pf_inst; 
  assign xcpt_1_ae_inst=bufMask[1] ? buf__xcpt_ae_inst:io_imem_bits_xcpt_ae_inst; 
  assign _ic_replay_T_1=valid&~bufMask; 
  assign _ic_replay_T_2=io_imem_bits_replay ? _ic_replay_T_1:2'h0; 
  assign ic_replay=buf_replay|_ic_replay_T_2; 
  assign _T_10=~io_imem_valid|~io_imem_bits_btb_taken; 
  assign _T_11=io_imem_bits_btb_bridx>=pcWordBits; 
  assign _T_12=_T_10|_T_11; 
  assign _T_14=_T_12|reset; 
  assign _io_pc_T=nBufValid>1'h0; 
  assign _replay_T_5={1'b0,ic_replay[1]}; 
  assign _replay_T_7=~exp_io_rvc&_replay_T_5[0]; 
  assign _io_inst_0_bits_xcpt1_T_4={xcpt_1_pf_inst,xcpt_1_ae_inst}; 
  assign _io_inst_0_bits_xcpt1_T_5=exp_io_rvc ? 2'h0:_io_inst_0_bits_xcpt1_T_4; 
  assign _T_18=bufMask[0]&exp_io_rvc; 
  assign _T_21={1'b0,bufMask[1]}; 
  assign _T_23=_T_18|_T_21[0]; 
  assign io_imem_ready=_io_imem_ready_T_1&_io_imem_ready_T_6; 
  assign io_pc=_io_pc_T ? buf__pc:io_imem_bits_pc; 
  assign io_btb_resp_entry=_T_23 ? ibufBTBResp_entry:io_imem_bits_btb_entry; 
  assign io_btb_resp_bht_history=_T_23 ? ibufBTBResp_bht_history:io_imem_bits_btb_bht_history; 
  assign io_inst_0_valid=valid[0]&full_insn; 
  assign io_inst_0_bits_xcpt0_pf_inst=bufMask[0] ? buf__xcpt_pf_inst:io_imem_bits_xcpt_pf_inst; 
  assign io_inst_0_bits_xcpt0_ae_inst=bufMask[0] ? buf__xcpt_ae_inst:io_imem_bits_xcpt_ae_inst; 
  assign io_inst_0_bits_xcpt1_pf_inst=_io_inst_0_bits_xcpt1_T_5[1]; 
  assign io_inst_0_bits_xcpt1_ae_inst=_io_inst_0_bits_xcpt1_T_5[0]; 
  assign io_inst_0_bits_replay=ic_replay[0]|_replay_T_7; 
  assign io_inst_0_bits_rvc=exp_io_rvc; 
  assign io_inst_0_bits_inst_bits=exp_io_out_bits; 
  assign io_inst_0_bits_inst_rd=exp_io_out_rd; 
  assign io_inst_0_bits_inst_rs1=exp_io_out_rs1; 
  assign io_inst_0_bits_inst_rs2=exp_io_out_rs2; 
  assign io_inst_0_bits_inst_rs3=exp_io_out_rs3; 
  assign io_inst_0_bits_raw=_inst_T|_inst_T_2; 
  assign exp_io_in=_inst_T|_inst_T_2; 
  assign IBuf_cov_read_addr=IBuf_state; 
  assign IBuf_cov_read_data=IBuf_cov[IBuf_cov_read_addr]; 
  assign IBuf_cov_write_data=1'h1; 
  assign IBuf_cov_write_addr=IBuf_state; 
  assign IBuf_cov_write_mask=1'h1; 
  assign IBuf_cov_write_en=1'h1; 
  assign nBufValid_shl=nBufValid; 
  assign nBufValid_pad={1'h0,nBufValid_shl}; 
  assign buf__replay_shl={buf__replay,1'h0}; 
  assign buf__replay_pad=buf__replay_shl; 
  assign IBuf_xor0=nBufValid_pad^buf__replay_pad; 
  assign exp_sum=IBuf_covSum+exp_io_covSum; 
  assign io_covSum=exp_sum; 
  assign stopEn0=~_T_14; 
  assign exp_metaAssert_wire=exp_metaAssert; 
  assign IBuf_or0=stopEn0|exp_metaAssert_wire; 
  assign metaAssert=IBuf_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              nBufValid <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 nBufValid <=1'h0;
               end 
             else 
               begin 
                 nBufValid <=_GEN_46[0];
               end 
         if (metaReset)
            begin 
              buf__pc <=40'h0;
            end 
          else 
            if (io_inst_0_ready)
               begin 
                 if (_T_7)
                    begin 
                      buf__pc <=_buf_pc_T_6;
                    end 
               end 
         if (metaReset)
            begin 
              buf__data <=32'h0;
            end 
          else 
            if (io_inst_0_ready)
               begin 
                 if (_T_7)
                    begin 
                      buf__data <={16'b0,_buf_data_T_1[15:0]};
                    end 
               end 
         if (metaReset)
            begin 
              buf__xcpt_pf_inst <=1'h0;
            end 
          else 
            if (io_inst_0_ready)
               begin 
                 if (_T_7)
                    begin 
                      buf__xcpt_pf_inst <=io_imem_bits_xcpt_pf_inst;
                    end 
               end 
         if (metaReset)
            begin 
              buf__xcpt_ae_inst <=1'h0;
            end 
          else 
            if (io_inst_0_ready)
               begin 
                 if (_T_7)
                    begin 
                      buf__xcpt_ae_inst <=io_imem_bits_xcpt_ae_inst;
                    end 
               end 
         if (metaReset)
            begin 
              buf__replay <=1'h0;
            end 
          else 
            if (io_inst_0_ready)
               begin 
                 if (_T_7)
                    begin 
                      buf__replay <=io_imem_bits_replay;
                    end 
               end 
         if (metaReset)
            begin 
              ibufBTBResp_entry <=5'h0;
            end 
          else 
            if (io_inst_0_ready)
               begin 
                 if (_T_7)
                    begin 
                      ibufBTBResp_entry <=io_imem_bits_btb_entry;
                    end 
               end 
         if (metaReset)
            begin 
              ibufBTBResp_bht_history <=8'h0;
            end 
          else 
            if (io_inst_0_ready)
               begin 
                 if (_T_7)
                    begin 
                      ibufBTBResp_bht_history <=io_imem_bits_btb_bht_history;
                    end 
               end 
         if (~_T_14)
            begin $display("Assertion failed\n    at IBuf.scala:79 assert(!io.imem.valid || !io.imem.bits.btb.taken || io.imem.bits.btb.bridx >= pcWordBits)\n");
            end 
         if (~_T_14)
            begin $display("fatal");
            end 
         IBuf_state <=IBuf_xor0;
         if (!(IBuf_cov_read_data))
            begin 
              IBuf_covSum <=IBuf_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              IBuf_metaAssert <=1'h0;
            end 
          else 
            begin 
              IBuf_metaAssert <=IBuf_metaAssert|IBuf_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (IBuf_cov_write_en&IBuf_cov_write_mask)
            begin 
              IBuf_cov [IBuf_cov_write_addr]<=IBuf_cov_write_data;
            end 
       end
  
endmodule
 
module CSRFile (
  input clock,
  input reset,
  input io_ungated_clock,
  input io_interrupts_debug,
  input io_interrupts_mtip,
  input io_interrupts_msip,
  input io_interrupts_meip,
  input io_interrupts_seip,
  input io_hartid,
  input [11:0] io_rw_addr,
  input [2:0] io_rw_cmd,
  output [63:0] io_rw_rdata,
  input [63:0] io_rw_wdata,
  input [11:0] io_decode_0_csr,
  output io_decode_0_fp_illegal,
  output io_decode_0_fp_csr,
  output io_decode_0_read_illegal,
  output io_decode_0_write_illegal,
  output io_decode_0_write_flush,
  output io_decode_0_system_illegal,
  output io_csr_stall,
  output io_eret,
  output io_singleStep,
  output io_status_debug,
  output io_status_cease,
  output io_status_wfi,
  output [31:0] io_status_isa,
  output [1:0] io_status_dprv,
  output [1:0] io_status_prv,
  output io_status_sd,
  output [26:0] io_status_zero2,
  output [1:0] io_status_sxl,
  output [1:0] io_status_uxl,
  output io_status_sd_rv32,
  output [7:0] io_status_zero1,
  output io_status_tsr,
  output io_status_tw,
  output io_status_tvm,
  output io_status_mxr,
  output io_status_sum,
  output io_status_mprv,
  output [1:0] io_status_xs,
  output [1:0] io_status_fs,
  output [1:0] io_status_mpp,
  output [1:0] io_status_vs,
  output io_status_spp,
  output io_status_mpie,
  output io_status_hpie,
  output io_status_spie,
  output io_status_upie,
  output io_status_mie,
  output io_status_hie,
  output io_status_sie,
  output io_status_uie,
  output [3:0] io_ptbr_mode,
  output [43:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input io_exception,
  input io_retire,
  input [63:0] io_cause,
  input [39:0] io_pc,
  input [39:0] io_tval,
  output [63:0] io_time,
  output [2:0] io_fcsr_rm,
  input io_fcsr_flags_valid,
  input [4:0] io_fcsr_flags_bits,
  output io_interrupt,
  output [63:0] io_interrupt_cause,
  output io_bp_0_control_action,
  output [1:0] io_bp_0_control_tmatch,
  output io_bp_0_control_m,
  output io_bp_0_control_s,
  output io_bp_0_control_u,
  output io_bp_0_control_x,
  output io_bp_0_control_w,
  output io_bp_0_control_r,
  output [38:0] io_bp_0_address,
  output io_pmp_0_cfg_l,
  output [1:0] io_pmp_0_cfg_a,
  output io_pmp_0_cfg_x,
  output io_pmp_0_cfg_w,
  output io_pmp_0_cfg_r,
  output [29:0] io_pmp_0_addr,
  output [31:0] io_pmp_0_mask,
  output io_pmp_1_cfg_l,
  output [1:0] io_pmp_1_cfg_a,
  output io_pmp_1_cfg_x,
  output io_pmp_1_cfg_w,
  output io_pmp_1_cfg_r,
  output [29:0] io_pmp_1_addr,
  output [31:0] io_pmp_1_mask,
  output io_pmp_2_cfg_l,
  output [1:0] io_pmp_2_cfg_a,
  output io_pmp_2_cfg_x,
  output io_pmp_2_cfg_w,
  output io_pmp_2_cfg_r,
  output [29:0] io_pmp_2_addr,
  output [31:0] io_pmp_2_mask,
  output io_pmp_3_cfg_l,
  output [1:0] io_pmp_3_cfg_a,
  output io_pmp_3_cfg_x,
  output io_pmp_3_cfg_w,
  output io_pmp_3_cfg_r,
  output [29:0] io_pmp_3_addr,
  output [31:0] io_pmp_3_mask,
  output io_pmp_4_cfg_l,
  output [1:0] io_pmp_4_cfg_a,
  output io_pmp_4_cfg_x,
  output io_pmp_4_cfg_w,
  output io_pmp_4_cfg_r,
  output [29:0] io_pmp_4_addr,
  output [31:0] io_pmp_4_mask,
  output io_pmp_5_cfg_l,
  output [1:0] io_pmp_5_cfg_a,
  output io_pmp_5_cfg_x,
  output io_pmp_5_cfg_w,
  output io_pmp_5_cfg_r,
  output [29:0] io_pmp_5_addr,
  output [31:0] io_pmp_5_mask,
  output io_pmp_6_cfg_l,
  output [1:0] io_pmp_6_cfg_a,
  output io_pmp_6_cfg_x,
  output io_pmp_6_cfg_w,
  output io_pmp_6_cfg_r,
  output [29:0] io_pmp_6_addr,
  output [31:0] io_pmp_6_mask,
  output io_pmp_7_cfg_l,
  output [1:0] io_pmp_7_cfg_a,
  output io_pmp_7_cfg_x,
  output io_pmp_7_cfg_w,
  output io_pmp_7_cfg_r,
  output [29:0] io_pmp_7_addr,
  output [31:0] io_pmp_7_mask,
  output io_inhibit_cycle,
  input [31:0] io_inst_0,
  output io_trace_0_valid,
  output [39:0] io_trace_0_iaddr,
  output [31:0] io_trace_0_insn,
  output [2:0] io_trace_0_priv,
  output io_trace_0_exception,
  output io_trace_0_interrupt,
  output [63:0] io_trace_0_cause,
  output [39:0] io_trace_0_tval,
  output [63:0] io_customCSRs_0_value,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg rv_dv ;  
   reg [1:0] reg_mstatus_prv ;  
   reg [31:0] _RAND_0 ;  
   reg reg_mstatus_tsr ;  
   reg [31:0] _RAND_1 ;  
   reg reg_mstatus_tw ;  
   reg [31:0] _RAND_2 ;  
   reg reg_mstatus_tvm ;  
   reg [31:0] _RAND_3 ;  
   reg reg_mstatus_mxr ;  
   reg [31:0] _RAND_4 ;  
   reg reg_mstatus_sum ;  
   reg [31:0] _RAND_5 ;  
   reg reg_mstatus_mprv ;  
   reg [31:0] _RAND_6 ;  
   reg [1:0] reg_mstatus_fs ;  
   reg [31:0] _RAND_7 ;  
   reg [1:0] reg_mstatus_mpp ;  
   reg [31:0] _RAND_8 ;  
   reg reg_mstatus_spp ;  
   reg [31:0] _RAND_9 ;  
   reg reg_mstatus_mpie ;  
   reg [31:0] _RAND_10 ;  
   reg reg_mstatus_spie ;  
   reg [31:0] _RAND_11 ;  
   reg reg_mstatus_mie ;  
   reg [31:0] _RAND_12 ;  
   reg reg_mstatus_sie ;  
   reg [31:0] _RAND_13 ;  
   wire system_insn ;  
   wire [31:0] _T_192 ;  
   wire [31:0] _T_199 ;  
   wire _T_200 ;  
   wire [31:0] _T_201 ;  
   wire _T_202 ;  
   wire _T_204 ;  
   wire insn_ret ;  
   wire _T_406 ;  
   reg [1:0] reg_dcsr_prv ;  
   reg [31:0] _RAND_14 ;  
   wire [1:0] _GEN_149 ;  
   wire [1:0] ret_prv ;  
   wire [31:0] _T_193 ;  
   wire _T_194 ;  
   wire insn_call ;  
   wire _T_197 ;  
   wire insn_break ;  
   wire _exception_T ;  
   wire exception ;  
   reg reg_singleStepped ;  
   reg [31:0] _RAND_15 ;  
   wire [3:0] _GEN_20 ;  
   wire [3:0] _cause_T_1 ;  
   wire [63:0] _cause_T_2 ;  
   wire [63:0] cause ;  
   wire [7:0] cause_lsbs ;  
   wire _causeIsDebugInt_T_1 ;  
   wire causeIsDebugInt ;  
   wire _trapToDebug_T ;  
   wire causeIsDebugTrigger ;  
   wire _trapToDebug_T_1 ;  
   wire _causeIsDebugBreak_T_2 ;  
   reg reg_dcsr_ebreakm ;  
   reg [31:0] _RAND_16 ;  
   reg reg_dcsr_ebreaks ;  
   reg [31:0] _RAND_17 ;  
   reg reg_dcsr_ebreaku ;  
   reg [31:0] _RAND_18 ;  
   wire [3:0] _causeIsDebugBreak_T_3 ;  
   wire [3:0] _causeIsDebugBreak_T_4 ;  
   wire causeIsDebugBreak ;  
   wire _trapToDebug_T_2 ;  
   reg reg_debug ;  
   reg [31:0] _RAND_19 ;  
   wire trapToDebug ;  
   wire [1:0] _GEN_56 ;  
   reg reg_rnmie ;  
   reg [31:0] _RAND_20 ;  
   reg reg_unmie ;  
   reg [31:0] _RAND_21 ;  
   wire _delegate_T ;  
   reg [63:0] reg_mideleg ;  
   reg [63:0] _RAND_22 ;  
   wire [63:0] read_mideleg ;  
   wire [63:0] _delegate_T_3 ;  
   reg [63:0] reg_medeleg ;  
   reg [63:0] _RAND_23 ;  
   wire [63:0] read_medeleg ;  
   wire [63:0] _delegate_T_5 ;  
   wire _delegate_T_7 ;  
   wire delegate ;  
   wire nmie ;  
   wire _T_279 ;  
   wire [1:0] _GEN_70 ;  
   wire [1:0] _GEN_100 ;  
   wire [1:0] _GEN_123 ;  
   wire [1:0] new_prv ;  
   wire _reg_mstatus_prv_T ;  
   reg [2:0] reg_dcsr_cause ;  
   reg [31:0] _RAND_24 ;  
   reg reg_dcsr_step ;  
   reg [31:0] _RAND_25 ;  
   reg [39:0] reg_dpc ;  
   reg [63:0] _RAND_26 ;  
   reg [63:0] reg_dscratch ;  
   reg [63:0] _RAND_27 ;  
   reg reg_bp_0_control_dmode ;  
   reg [31:0] _RAND_28 ;  
   reg reg_bp_0_control_action ;  
   reg [31:0] _RAND_29 ;  
   reg [1:0] reg_bp_0_control_tmatch ;  
   reg [31:0] _RAND_30 ;  
   reg reg_bp_0_control_m ;  
   reg [31:0] _RAND_31 ;  
   reg reg_bp_0_control_s ;  
   reg [31:0] _RAND_32 ;  
   reg reg_bp_0_control_u ;  
   reg [31:0] _RAND_33 ;  
   reg reg_bp_0_control_x ;  
   reg [31:0] _RAND_34 ;  
   reg reg_bp_0_control_w ;  
   reg [31:0] _RAND_35 ;  
   reg reg_bp_0_control_r ;  
   reg [31:0] _RAND_36 ;  
   reg [38:0] reg_bp_0_address ;  
   reg [63:0] _RAND_37 ;  
   reg reg_pmp_0_cfg_l ;  
   reg [31:0] _RAND_38 ;  
   reg [1:0] reg_pmp_0_cfg_a ;  
   reg [31:0] _RAND_39 ;  
   reg reg_pmp_0_cfg_x ;  
   reg [31:0] _RAND_40 ;  
   reg reg_pmp_0_cfg_w ;  
   reg [31:0] _RAND_41 ;  
   reg reg_pmp_0_cfg_r ;  
   reg [31:0] _RAND_42 ;  
   reg [29:0] reg_pmp_0_addr ;  
   reg [31:0] _RAND_43 ;  
   reg reg_pmp_1_cfg_l ;  
   reg [31:0] _RAND_44 ;  
   reg [1:0] reg_pmp_1_cfg_a ;  
   reg [31:0] _RAND_45 ;  
   reg reg_pmp_1_cfg_x ;  
   reg [31:0] _RAND_46 ;  
   reg reg_pmp_1_cfg_w ;  
   reg [31:0] _RAND_47 ;  
   reg reg_pmp_1_cfg_r ;  
   reg [31:0] _RAND_48 ;  
   reg [29:0] reg_pmp_1_addr ;  
   reg [31:0] _RAND_49 ;  
   reg reg_pmp_2_cfg_l ;  
   reg [31:0] _RAND_50 ;  
   reg [1:0] reg_pmp_2_cfg_a ;  
   reg [31:0] _RAND_51 ;  
   reg reg_pmp_2_cfg_x ;  
   reg [31:0] _RAND_52 ;  
   reg reg_pmp_2_cfg_w ;  
   reg [31:0] _RAND_53 ;  
   reg reg_pmp_2_cfg_r ;  
   reg [31:0] _RAND_54 ;  
   reg [29:0] reg_pmp_2_addr ;  
   reg [31:0] _RAND_55 ;  
   reg reg_pmp_3_cfg_l ;  
   reg [31:0] _RAND_56 ;  
   reg [1:0] reg_pmp_3_cfg_a ;  
   reg [31:0] _RAND_57 ;  
   reg reg_pmp_3_cfg_x ;  
   reg [31:0] _RAND_58 ;  
   reg reg_pmp_3_cfg_w ;  
   reg [31:0] _RAND_59 ;  
   reg reg_pmp_3_cfg_r ;  
   reg [31:0] _RAND_60 ;  
   reg [29:0] reg_pmp_3_addr ;  
   reg [31:0] _RAND_61 ;  
   reg reg_pmp_4_cfg_l ;  
   reg [31:0] _RAND_62 ;  
   reg [1:0] reg_pmp_4_cfg_a ;  
   reg [31:0] _RAND_63 ;  
   reg reg_pmp_4_cfg_x ;  
   reg [31:0] _RAND_64 ;  
   reg reg_pmp_4_cfg_w ;  
   reg [31:0] _RAND_65 ;  
   reg reg_pmp_4_cfg_r ;  
   reg [31:0] _RAND_66 ;  
   reg [29:0] reg_pmp_4_addr ;  
   reg [31:0] _RAND_67 ;  
   reg reg_pmp_5_cfg_l ;  
   reg [31:0] _RAND_68 ;  
   reg [1:0] reg_pmp_5_cfg_a ;  
   reg [31:0] _RAND_69 ;  
   reg reg_pmp_5_cfg_x ;  
   reg [31:0] _RAND_70 ;  
   reg reg_pmp_5_cfg_w ;  
   reg [31:0] _RAND_71 ;  
   reg reg_pmp_5_cfg_r ;  
   reg [31:0] _RAND_72 ;  
   reg [29:0] reg_pmp_5_addr ;  
   reg [31:0] _RAND_73 ;  
   reg reg_pmp_6_cfg_l ;  
   reg [31:0] _RAND_74 ;  
   reg [1:0] reg_pmp_6_cfg_a ;  
   reg [31:0] _RAND_75 ;  
   reg reg_pmp_6_cfg_x ;  
   reg [31:0] _RAND_76 ;  
   reg reg_pmp_6_cfg_w ;  
   reg [31:0] _RAND_77 ;  
   reg reg_pmp_6_cfg_r ;  
   reg [31:0] _RAND_78 ;  
   reg [29:0] reg_pmp_6_addr ;  
   reg [31:0] _RAND_79 ;  
   reg reg_pmp_7_cfg_l ;  
   reg [31:0] _RAND_80 ;  
   reg [1:0] reg_pmp_7_cfg_a ;  
   reg [31:0] _RAND_81 ;  
   reg reg_pmp_7_cfg_x ;  
   reg [31:0] _RAND_82 ;  
   reg reg_pmp_7_cfg_w ;  
   reg [31:0] _RAND_83 ;  
   reg reg_pmp_7_cfg_r ;  
   reg [31:0] _RAND_84 ;  
   reg [29:0] reg_pmp_7_addr ;  
   reg [31:0] _RAND_85 ;  
   reg [63:0] reg_mie ;  
   reg [63:0] _RAND_86 ;  
   reg reg_mip_seip ;  
   reg [31:0] _RAND_87 ;  
   reg reg_mip_stip ;  
   reg [31:0] _RAND_88 ;  
   reg reg_mip_ssip ;  
   reg [31:0] _RAND_89 ;  
   reg [39:0] reg_mepc ;  
   reg [63:0] _RAND_90 ;  
   reg [63:0] reg_mcause ;  
   reg [63:0] _RAND_91 ;  
   reg [39:0] reg_mtval ;  
   reg [63:0] _RAND_92 ;  
   reg [63:0] reg_mscratch ;  
   reg [63:0] _RAND_93 ;  
   reg [31:0] reg_mtvec ;  
   reg [31:0] _RAND_94 ;  
   reg [31:0] reg_mcounteren ;  
   reg [31:0] _RAND_95 ;  
   wire [31:0] read_mcounteren ;  
   reg [31:0] reg_scounteren ;  
   reg [31:0] _RAND_96 ;  
   wire [31:0] read_scounteren ;  
   reg [39:0] reg_sepc ;  
   reg [63:0] _RAND_97 ;  
   reg [63:0] reg_scause ;  
   reg [63:0] _RAND_98 ;  
   reg [39:0] reg_stval ;  
   reg [63:0] _RAND_99 ;  
   reg [63:0] reg_sscratch ;  
   reg [63:0] _RAND_100 ;  
   reg [38:0] reg_stvec ;  
   reg [63:0] _RAND_101 ;  
   reg [3:0] reg_satp_mode ;  
   reg [31:0] _RAND_102 ;  
   reg [43:0] reg_satp_ppn ;  
   reg [63:0] _RAND_103 ;  
   reg reg_wfi ;  
   reg [31:0] _RAND_104 ;  
   reg [4:0] reg_fflags ;  
   reg [31:0] _RAND_105 ;  
   reg [2:0] reg_frm ;  
   reg [31:0] _RAND_106 ;  
   reg [2:0] reg_mcountinhibit ;  
   reg [31:0] _RAND_107 ;  
   wire x67 ;  
   reg [5:0] value_lo ;  
   reg [31:0] _RAND_108 ;  
   wire [5:0] _GEN_23 ;  
   wire [6:0] nextSmall ;  
   wire [6:0] _GEN_0 ;  
   reg [57:0] value_hi ;  
   reg [63:0] _RAND_109 ;  
   wire _large_T_2 ;  
   wire [57:0] _large_r_T_1 ;  
   wire [63:0] value ;  
   reg [5:0] value_lo_1 ;  
   reg [31:0] _RAND_110 ;  
   wire [6:0] nextSmall_1 ;  
   wire [6:0] _GEN_2 ;  
   reg [57:0] value_hi_1 ;  
   reg [63:0] _RAND_111 ;  
   wire _large_T_5 ;  
   wire [57:0] _large_r_T_3 ;  
   wire [63:0] value_1 ;  
   wire mip_seip ;  
   wire [7:0] read_mip_lo ;  
   wire [15:0] _read_mip_T ;  
   wire [15:0] read_mip ;  
   wire [63:0] _GEN_45 ;  
   wire [63:0] pending_interrupts ;  
   wire [14:0] d_interrupts ;  
   wire _m_interrupts_T_1 ;  
   wire _m_interrupts_T_2 ;  
   wire [63:0] _m_interrupts_T_4 ;  
   wire [63:0] m_interrupts ;  
   wire _s_interrupts_T ;  
   wire _s_interrupts_T_1 ;  
   wire _s_interrupts_T_2 ;  
   wire _s_interrupts_T_3 ;  
   wire _s_interrupts_T_4 ;  
   wire [63:0] _s_interrupts_T_5 ;  
   wire [63:0] s_interrupts ;  
   wire _any_T_38 ;  
   wire _any_T_39 ;  
   wire _any_T_40 ;  
   wire _any_T_41 ;  
   wire _any_T_42 ;  
   wire _any_T_43 ;  
   wire _any_T_44 ;  
   wire _any_T_45 ;  
   wire _any_T_46 ;  
   wire _any_T_47 ;  
   wire _any_T_48 ;  
   wire _any_T_50 ;  
   wire _any_T_51 ;  
   wire _any_T_52 ;  
   wire _any_T_53 ;  
   wire _any_T_54 ;  
   wire _any_T_55 ;  
   wire _any_T_56 ;  
   wire _any_T_57 ;  
   wire _any_T_58 ;  
   wire _any_T_59 ;  
   wire _any_T_60 ;  
   wire _any_T_61 ;  
   wire _any_T_62 ;  
   wire _any_T_63 ;  
   wire _any_T_64 ;  
   wire _any_T_65 ;  
   wire _any_T_66 ;  
   wire _any_T_67 ;  
   wire _any_T_68 ;  
   wire _any_T_69 ;  
   wire _any_T_70 ;  
   wire _any_T_71 ;  
   wire _any_T_72 ;  
   wire _any_T_73 ;  
   wire _any_T_74 ;  
   wire anyInterrupt ;  
   wire [2:0] _which_T_38 ;  
   wire [3:0] _which_T_39 ;  
   wire [3:0] _which_T_40 ;  
   wire [3:0] _which_T_41 ;  
   wire [3:0] _which_T_42 ;  
   wire [3:0] _which_T_43 ;  
   wire [3:0] _which_T_44 ;  
   wire [3:0] _which_T_45 ;  
   wire [3:0] _which_T_46 ;  
   wire [3:0] _which_T_47 ;  
   wire [3:0] _which_T_48 ;  
   wire [3:0] _which_T_49 ;  
   wire [3:0] _which_T_50 ;  
   wire [3:0] _which_T_51 ;  
   wire [3:0] _which_T_52 ;  
   wire [3:0] _which_T_53 ;  
   wire [3:0] _which_T_54 ;  
   wire [3:0] _which_T_55 ;  
   wire [3:0] _which_T_56 ;  
   wire [3:0] _which_T_57 ;  
   wire [3:0] _which_T_58 ;  
   wire [3:0] _which_T_59 ;  
   wire [3:0] _which_T_60 ;  
   wire [3:0] _which_T_61 ;  
   wire [3:0] _which_T_62 ;  
   wire [3:0] _which_T_64 ;  
   wire [3:0] _which_T_65 ;  
   wire [3:0] _which_T_66 ;  
   wire [3:0] _which_T_67 ;  
   wire [3:0] _which_T_68 ;  
   wire [3:0] _which_T_69 ;  
   wire [3:0] _which_T_70 ;  
   wire [3:0] _which_T_71 ;  
   wire [3:0] _which_T_72 ;  
   wire [3:0] _which_T_73 ;  
   wire [3:0] _which_T_74 ;  
   wire [3:0] whichInterrupt ;  
   wire [63:0] _GEN_556 ;  
   wire _io_interrupt_T_1 ;  
   wire _io_interrupt_T_2 ;  
   wire _io_interrupt_T_3 ;  
   wire pmp_mask_base_lo ;  
   wire [30:0] pmp_mask_base ;  
   wire [30:0] _pmp_mask_T_1 ;  
   wire [30:0] pmp_mask_hi ;  
   wire [32:0] _pmp_mask_T_3 ;  
   wire pmp_mask_base_lo_1 ;  
   wire [30:0] pmp_mask_base_1 ;  
   wire [30:0] _pmp_mask_T_5 ;  
   wire [30:0] pmp_mask_hi_1 ;  
   wire [32:0] _pmp_mask_T_7 ;  
   wire pmp_mask_base_lo_2 ;  
   wire [30:0] pmp_mask_base_2 ;  
   wire [30:0] _pmp_mask_T_9 ;  
   wire [30:0] pmp_mask_hi_2 ;  
   wire [32:0] _pmp_mask_T_11 ;  
   wire pmp_mask_base_lo_3 ;  
   wire [30:0] pmp_mask_base_3 ;  
   wire [30:0] _pmp_mask_T_13 ;  
   wire [30:0] pmp_mask_hi_3 ;  
   wire [32:0] _pmp_mask_T_15 ;  
   wire pmp_mask_base_lo_4 ;  
   wire [30:0] pmp_mask_base_4 ;  
   wire [30:0] _pmp_mask_T_17 ;  
   wire [30:0] pmp_mask_hi_4 ;  
   wire [32:0] _pmp_mask_T_19 ;  
   wire pmp_mask_base_lo_5 ;  
   wire [30:0] pmp_mask_base_5 ;  
   wire [30:0] _pmp_mask_T_21 ;  
   wire [30:0] pmp_mask_hi_5 ;  
   wire [32:0] _pmp_mask_T_23 ;  
   wire pmp_mask_base_lo_6 ;  
   wire [30:0] pmp_mask_base_6 ;  
   wire [30:0] _pmp_mask_T_25 ;  
   wire [30:0] pmp_mask_hi_6 ;  
   wire [32:0] _pmp_mask_T_27 ;  
   wire pmp_mask_base_lo_7 ;  
   wire [30:0] pmp_mask_base_7 ;  
   wire [30:0] _pmp_mask_T_29 ;  
   wire [30:0] pmp_mask_hi_7 ;  
   wire [32:0] _pmp_mask_T_31 ;  
   reg [63:0] reg_misa ;  
   reg [63:0] _RAND_112 ;  
   wire [6:0] read_mstatus_lo_lo ;  
   wire [18:0] read_mstatus_lo ;  
   wire [16:0] read_mstatus_hi_lo ;  
   wire [102:0] _read_mstatus_T ;  
   wire [63:0] read_mstatus ;  
   wire [7:0] _read_mtvec_T_1 ;  
   wire [31:0] _read_mtvec_T_3 ;  
   wire [31:0] read_mtvec_lo ;  
   wire [63:0] read_mtvec ;  
   wire [7:0] _read_stvec_T_1 ;  
   wire [38:0] _read_stvec_T_3 ;  
   wire [38:0] read_stvec_lo ;  
   wire [24:0] read_stvec_hi ;  
   wire [63:0] read_stvec ;  
   wire [6:0] lo_2 ;  
   wire [63:0] _T_7 ;  
   wire [24:0] hi_3 ;  
   wire [63:0] _T_10 ;  
   wire [1:0] _T_14 ;  
   wire [39:0] _GEN_557 ;  
   wire [39:0] _T_15 ;  
   wire [39:0] lo_4 ;  
   wire [23:0] hi_5 ;  
   wire [63:0] _T_18 ;  
   wire [23:0] hi_6 ;  
   wire [63:0] _T_21 ;  
   wire [11:0] lo_5 ;  
   wire [31:0] _T_22 ;  
   wire [39:0] _T_26 ;  
   wire [39:0] lo_6 ;  
   wire [23:0] hi_8 ;  
   wire [63:0] _T_29 ;  
   wire [7:0] read_fcsr ;  
   wire [63:0] read_sie ;  
   wire [63:0] read_sip ;  
   wire [6:0] lo_lo_4 ;  
   wire [18:0] lo_7 ;  
   wire [16:0] hi_lo_4 ;  
   wire [102:0] _T_30 ;  
   wire [23:0] hi_10 ;  
   wire [63:0] _T_34 ;  
   wire [63:0] _T_35 ;  
   wire [39:0] _T_39 ;  
   wire [39:0] lo_8 ;  
   wire [23:0] hi_12 ;  
   wire [63:0] _T_42 ;  
   wire [7:0] lo_lo_lo_3 ;  
   wire [7:0] lo_hi_lo_5 ;  
   wire [7:0] hi_lo_lo_4 ;  
   wire [7:0] hi_hi_lo_5 ;  
   wire [15:0] lo_lo_5 ;  
   wire [31:0] lo_17 ;  
   wire [15:0] hi_lo_5 ;  
   wire [63:0] _T_43 ;  
   reg [63:0] reg_custom_0 ;  
   reg [63:0] _RAND_113 ;  
   wire _T_46 ;  
   wire _T_47 ;  
   wire _T_49 ;  
   wire _T_50 ;  
   wire _T_51 ;  
   wire _T_52 ;  
   wire _T_53 ;  
   wire _T_54 ;  
   wire _T_55 ;  
   wire _T_56 ;  
   wire _T_57 ;  
   wire _T_58 ;  
   wire _T_59 ;  
   wire _T_60 ;  
   wire _T_61 ;  
   wire _T_62 ;  
   wire _T_63 ;  
   wire _T_64 ;  
   wire _T_65 ;  
   wire _T_66 ;  
   wire _T_67 ;  
   wire _T_155 ;  
   wire _T_156 ;  
   wire _T_157 ;  
   wire _T_158 ;  
   wire _T_159 ;  
   wire _T_160 ;  
   wire _T_161 ;  
   wire _T_162 ;  
   wire _T_163 ;  
   wire _T_164 ;  
   wire _T_165 ;  
   wire _T_166 ;  
   wire _T_167 ;  
   wire _T_168 ;  
   wire _T_169 ;  
   wire _T_170 ;  
   wire _T_172 ;  
   wire _T_173 ;  
   wire _T_174 ;  
   wire _T_175 ;  
   wire _T_176 ;  
   wire _T_177 ;  
   wire _T_178 ;  
   wire _T_179 ;  
   wire _T_188 ;  
   wire _T_189 ;  
   wire _T_191 ;  
   wire [63:0] _wdata_T_1 ;  
   wire [63:0] _wdata_T_2 ;  
   wire _wdata_T_4 ;  
   wire [63:0] _wdata_T_5 ;  
   wire [63:0] wdata ;  
   wire [31:0] _T_205 ;  
   wire _T_206 ;  
   wire [31:0] _T_208 ;  
   wire _T_209 ;  
   wire insn_cease ;  
   wire insn_wfi ;  
   wire [31:0] _T_220 ;  
   wire [31:0] _T_227 ;  
   wire _T_228 ;  
   wire [31:0] _T_229 ;  
   wire _T_230 ;  
   wire is_ret ;  
   wire [31:0] _T_236 ;  
   wire is_wfi ;  
   wire [31:0] _T_239 ;  
   wire is_sfence ;  
   wire _allow_wfi_T ;  
   wire allow_wfi ;  
   wire allow_sfence_vma ;  
   wire allow_sret ;  
   wire [4:0] counter_addr ;  
   wire [31:0] _allow_counter_T_1 ;  
   wire _allow_counter_T_3 ;  
   wire _allow_counter_T_4 ;  
   wire [31:0] _allow_counter_T_6 ;  
   wire _allow_counter_T_8 ;  
   wire allow_counter ;  
   wire _io_decode_0_fp_illegal_T ;  
   wire [11:0] _io_decode_0_fp_csr_T ;  
   wire _io_decode_0_read_illegal_T_1 ;  
   wire _io_decode_0_read_illegal_T_2 ;  
   wire _io_decode_0_read_illegal_T_3 ;  
   wire _io_decode_0_read_illegal_T_4 ;  
   wire _io_decode_0_read_illegal_T_5 ;  
   wire _io_decode_0_read_illegal_T_6 ;  
   wire _io_decode_0_read_illegal_T_7 ;  
   wire _io_decode_0_read_illegal_T_8 ;  
   wire _io_decode_0_read_illegal_T_9 ;  
   wire _io_decode_0_read_illegal_T_10 ;  
   wire _io_decode_0_read_illegal_T_11 ;  
   wire _io_decode_0_read_illegal_T_12 ;  
   wire _io_decode_0_read_illegal_T_13 ;  
   wire _io_decode_0_read_illegal_T_14 ;  
   wire _io_decode_0_read_illegal_T_15 ;  
   wire _io_decode_0_read_illegal_T_16 ;  
   wire _io_decode_0_read_illegal_T_17 ;  
   wire _io_decode_0_read_illegal_T_18 ;  
   wire _io_decode_0_read_illegal_T_19 ;  
   wire _io_decode_0_read_illegal_T_20 ;  
   wire _io_decode_0_read_illegal_T_21 ;  
   wire _io_decode_0_read_illegal_T_22 ;  
   wire _io_decode_0_read_illegal_T_23 ;  
   wire _io_decode_0_read_illegal_T_24 ;  
   wire _io_decode_0_read_illegal_T_25 ;  
   wire _io_decode_0_read_illegal_T_26 ;  
   wire _io_decode_0_read_illegal_T_27 ;  
   wire _io_decode_0_read_illegal_T_28 ;  
   wire _io_decode_0_read_illegal_T_29 ;  
   wire _io_decode_0_read_illegal_T_30 ;  
   wire _io_decode_0_read_illegal_T_31 ;  
   wire _io_decode_0_read_illegal_T_32 ;  
   wire _io_decode_0_read_illegal_T_33 ;  
   wire _io_decode_0_read_illegal_T_34 ;  
   wire _io_decode_0_read_illegal_T_35 ;  
   wire _io_decode_0_read_illegal_T_36 ;  
   wire _io_decode_0_read_illegal_T_37 ;  
   wire _io_decode_0_read_illegal_T_38 ;  
   wire _io_decode_0_read_illegal_T_39 ;  
   wire _io_decode_0_read_illegal_T_40 ;  
   wire _io_decode_0_read_illegal_T_41 ;  
   wire _io_decode_0_read_illegal_T_42 ;  
   wire _io_decode_0_read_illegal_T_43 ;  
   wire _io_decode_0_read_illegal_T_44 ;  
   wire _io_decode_0_read_illegal_T_45 ;  
   wire _io_decode_0_read_illegal_T_46 ;  
   wire _io_decode_0_read_illegal_T_47 ;  
   wire _io_decode_0_read_illegal_T_48 ;  
   wire _io_decode_0_read_illegal_T_49 ;  
   wire _io_decode_0_read_illegal_T_50 ;  
   wire _io_decode_0_read_illegal_T_51 ;  
   wire _io_decode_0_read_illegal_T_52 ;  
   wire _io_decode_0_read_illegal_T_53 ;  
   wire _io_decode_0_read_illegal_T_54 ;  
   wire _io_decode_0_read_illegal_T_55 ;  
   wire _io_decode_0_read_illegal_T_56 ;  
   wire _io_decode_0_read_illegal_T_57 ;  
   wire _io_decode_0_read_illegal_T_58 ;  
   wire _io_decode_0_read_illegal_T_59 ;  
   wire _io_decode_0_read_illegal_T_60 ;  
   wire _io_decode_0_read_illegal_T_61 ;  
   wire _io_decode_0_read_illegal_T_62 ;  
   wire _io_decode_0_read_illegal_T_63 ;  
   wire _io_decode_0_read_illegal_T_64 ;  
   wire _io_decode_0_read_illegal_T_65 ;  
   wire _io_decode_0_read_illegal_T_66 ;  
   wire _io_decode_0_read_illegal_T_67 ;  
   wire _io_decode_0_read_illegal_T_68 ;  
   wire _io_decode_0_read_illegal_T_69 ;  
   wire _io_decode_0_read_illegal_T_70 ;  
   wire _io_decode_0_read_illegal_T_71 ;  
   wire _io_decode_0_read_illegal_T_72 ;  
   wire _io_decode_0_read_illegal_T_73 ;  
   wire _io_decode_0_read_illegal_T_74 ;  
   wire _io_decode_0_read_illegal_T_75 ;  
   wire _io_decode_0_read_illegal_T_76 ;  
   wire _io_decode_0_read_illegal_T_77 ;  
   wire _io_decode_0_read_illegal_T_78 ;  
   wire _io_decode_0_read_illegal_T_79 ;  
   wire _io_decode_0_read_illegal_T_80 ;  
   wire _io_decode_0_read_illegal_T_81 ;  
   wire _io_decode_0_read_illegal_T_82 ;  
   wire _io_decode_0_read_illegal_T_83 ;  
   wire _io_decode_0_read_illegal_T_84 ;  
   wire _io_decode_0_read_illegal_T_85 ;  
   wire _io_decode_0_read_illegal_T_86 ;  
   wire _io_decode_0_read_illegal_T_87 ;  
   wire _io_decode_0_read_illegal_T_88 ;  
   wire _io_decode_0_read_illegal_T_89 ;  
   wire _io_decode_0_read_illegal_T_90 ;  
   wire _io_decode_0_read_illegal_T_91 ;  
   wire _io_decode_0_read_illegal_T_92 ;  
   wire _io_decode_0_read_illegal_T_93 ;  
   wire _io_decode_0_read_illegal_T_94 ;  
   wire _io_decode_0_read_illegal_T_95 ;  
   wire _io_decode_0_read_illegal_T_96 ;  
   wire _io_decode_0_read_illegal_T_97 ;  
   wire _io_decode_0_read_illegal_T_98 ;  
   wire _io_decode_0_read_illegal_T_99 ;  
   wire _io_decode_0_read_illegal_T_100 ;  
   wire _io_decode_0_read_illegal_T_101 ;  
   wire _io_decode_0_read_illegal_T_102 ;  
   wire _io_decode_0_read_illegal_T_103 ;  
   wire _io_decode_0_read_illegal_T_104 ;  
   wire _io_decode_0_read_illegal_T_105 ;  
   wire _io_decode_0_read_illegal_T_106 ;  
   wire _io_decode_0_read_illegal_T_107 ;  
   wire _io_decode_0_read_illegal_T_108 ;  
   wire _io_decode_0_read_illegal_T_109 ;  
   wire _io_decode_0_read_illegal_T_110 ;  
   wire _io_decode_0_read_illegal_T_111 ;  
   wire _io_decode_0_read_illegal_T_112 ;  
   wire _io_decode_0_read_illegal_T_113 ;  
   wire _io_decode_0_read_illegal_T_114 ;  
   wire _io_decode_0_read_illegal_T_115 ;  
   wire _io_decode_0_read_illegal_T_116 ;  
   wire _io_decode_0_read_illegal_T_117 ;  
   wire _io_decode_0_read_illegal_T_118 ;  
   wire _io_decode_0_read_illegal_T_119 ;  
   wire _io_decode_0_read_illegal_T_120 ;  
   wire _io_decode_0_read_illegal_T_121 ;  
   wire _io_decode_0_read_illegal_T_122 ;  
   wire _io_decode_0_read_illegal_T_123 ;  
   wire _io_decode_0_read_illegal_T_124 ;  
   wire _io_decode_0_read_illegal_T_125 ;  
   wire _io_decode_0_read_illegal_T_126 ;  
   wire _io_decode_0_read_illegal_T_127 ;  
   wire _io_decode_0_read_illegal_T_128 ;  
   wire _io_decode_0_read_illegal_T_129 ;  
   wire _io_decode_0_read_illegal_T_130 ;  
   wire _io_decode_0_read_illegal_T_131 ;  
   wire _io_decode_0_read_illegal_T_132 ;  
   wire _io_decode_0_read_illegal_T_133 ;  
   wire _io_decode_0_read_illegal_T_134 ;  
   wire _io_decode_0_read_illegal_T_135 ;  
   wire _io_decode_0_read_illegal_T_136 ;  
   wire _io_decode_0_read_illegal_T_137 ;  
   wire _io_decode_0_read_illegal_T_138 ;  
   wire _io_decode_0_read_illegal_T_139 ;  
   wire _io_decode_0_read_illegal_T_140 ;  
   wire _io_decode_0_read_illegal_T_141 ;  
   wire _io_decode_0_read_illegal_T_142 ;  
   wire _io_decode_0_read_illegal_T_143 ;  
   wire _io_decode_0_read_illegal_T_144 ;  
   wire _io_decode_0_read_illegal_T_145 ;  
   wire _io_decode_0_read_illegal_T_146 ;  
   wire _io_decode_0_read_illegal_T_147 ;  
   wire _io_decode_0_read_illegal_T_148 ;  
   wire _io_decode_0_read_illegal_T_149 ;  
   wire _io_decode_0_read_illegal_T_150 ;  
   wire _io_decode_0_read_illegal_T_151 ;  
   wire _io_decode_0_read_illegal_T_152 ;  
   wire _io_decode_0_read_illegal_T_153 ;  
   wire _io_decode_0_read_illegal_T_154 ;  
   wire _io_decode_0_read_illegal_T_155 ;  
   wire _io_decode_0_read_illegal_T_156 ;  
   wire _io_decode_0_read_illegal_T_157 ;  
   wire _io_decode_0_read_illegal_T_158 ;  
   wire _io_decode_0_read_illegal_T_159 ;  
   wire _io_decode_0_read_illegal_T_160 ;  
   wire _io_decode_0_read_illegal_T_161 ;  
   wire _io_decode_0_read_illegal_T_162 ;  
   wire _io_decode_0_read_illegal_T_163 ;  
   wire _io_decode_0_read_illegal_T_164 ;  
   wire _io_decode_0_read_illegal_T_165 ;  
   wire _io_decode_0_read_illegal_T_166 ;  
   wire _io_decode_0_read_illegal_T_167 ;  
   wire _io_decode_0_read_illegal_T_168 ;  
   wire _io_decode_0_read_illegal_T_169 ;  
   wire _io_decode_0_read_illegal_T_170 ;  
   wire _io_decode_0_read_illegal_T_171 ;  
   wire _io_decode_0_read_illegal_T_172 ;  
   wire _io_decode_0_read_illegal_T_173 ;  
   wire _io_decode_0_read_illegal_T_174 ;  
   wire _io_decode_0_read_illegal_T_175 ;  
   wire _io_decode_0_read_illegal_T_176 ;  
   wire _io_decode_0_read_illegal_T_177 ;  
   wire _io_decode_0_read_illegal_T_178 ;  
   wire _io_decode_0_read_illegal_T_179 ;  
   wire _io_decode_0_read_illegal_T_180 ;  
   wire _io_decode_0_read_illegal_T_181 ;  
   wire _io_decode_0_read_illegal_T_182 ;  
   wire _io_decode_0_read_illegal_T_183 ;  
   wire _io_decode_0_read_illegal_T_184 ;  
   wire _io_decode_0_read_illegal_T_185 ;  
   wire _io_decode_0_read_illegal_T_186 ;  
   wire _io_decode_0_read_illegal_T_187 ;  
   wire _io_decode_0_read_illegal_T_188 ;  
   wire _io_decode_0_read_illegal_T_189 ;  
   wire _io_decode_0_read_illegal_T_190 ;  
   wire _io_decode_0_read_illegal_T_191 ;  
   wire _io_decode_0_read_illegal_T_192 ;  
   wire _io_decode_0_read_illegal_T_193 ;  
   wire _io_decode_0_read_illegal_T_194 ;  
   wire _io_decode_0_read_illegal_T_195 ;  
   wire _io_decode_0_read_illegal_T_196 ;  
   wire _io_decode_0_read_illegal_T_197 ;  
   wire _io_decode_0_read_illegal_T_198 ;  
   wire _io_decode_0_read_illegal_T_199 ;  
   wire _io_decode_0_read_illegal_T_200 ;  
   wire _io_decode_0_read_illegal_T_201 ;  
   wire _io_decode_0_read_illegal_T_202 ;  
   wire _io_decode_0_read_illegal_T_203 ;  
   wire _io_decode_0_read_illegal_T_204 ;  
   wire _io_decode_0_read_illegal_T_205 ;  
   wire _io_decode_0_read_illegal_T_206 ;  
   wire _io_decode_0_read_illegal_T_207 ;  
   wire _io_decode_0_read_illegal_T_208 ;  
   wire _io_decode_0_read_illegal_T_209 ;  
   wire _io_decode_0_read_illegal_T_210 ;  
   wire _io_decode_0_read_illegal_T_211 ;  
   wire _io_decode_0_read_illegal_T_212 ;  
   wire _io_decode_0_read_illegal_T_213 ;  
   wire _io_decode_0_read_illegal_T_214 ;  
   wire _io_decode_0_read_illegal_T_215 ;  
   wire _io_decode_0_read_illegal_T_216 ;  
   wire _io_decode_0_read_illegal_T_217 ;  
   wire _io_decode_0_read_illegal_T_218 ;  
   wire _io_decode_0_read_illegal_T_219 ;  
   wire _io_decode_0_read_illegal_T_220 ;  
   wire _io_decode_0_read_illegal_T_221 ;  
   wire _io_decode_0_read_illegal_T_222 ;  
   wire _io_decode_0_read_illegal_T_223 ;  
   wire _io_decode_0_read_illegal_T_224 ;  
   wire _io_decode_0_read_illegal_T_225 ;  
   wire _io_decode_0_read_illegal_T_226 ;  
   wire _io_decode_0_read_illegal_T_227 ;  
   wire _io_decode_0_read_illegal_T_228 ;  
   wire _io_decode_0_read_illegal_T_229 ;  
   wire _io_decode_0_read_illegal_T_230 ;  
   wire _io_decode_0_read_illegal_T_231 ;  
   wire _io_decode_0_read_illegal_T_232 ;  
   wire _io_decode_0_read_illegal_T_233 ;  
   wire _io_decode_0_read_illegal_T_234 ;  
   wire _io_decode_0_read_illegal_T_235 ;  
   wire _io_decode_0_read_illegal_T_236 ;  
   wire _io_decode_0_read_illegal_T_237 ;  
   wire _io_decode_0_read_illegal_T_238 ;  
   wire _io_decode_0_read_illegal_T_239 ;  
   wire _io_decode_0_read_illegal_T_240 ;  
   wire _io_decode_0_read_illegal_T_241 ;  
   wire _io_decode_0_read_illegal_T_242 ;  
   wire _io_decode_0_read_illegal_T_243 ;  
   wire _io_decode_0_read_illegal_T_244 ;  
   wire _io_decode_0_read_illegal_T_245 ;  
   wire _io_decode_0_read_illegal_T_246 ;  
   wire _io_decode_0_read_illegal_T_247 ;  
   wire _io_decode_0_read_illegal_T_248 ;  
   wire _io_decode_0_read_illegal_T_249 ;  
   wire _io_decode_0_read_illegal_T_250 ;  
   wire _io_decode_0_read_illegal_T_251 ;  
   wire _io_decode_0_read_illegal_T_252 ;  
   wire _io_decode_0_read_illegal_T_253 ;  
   wire _io_decode_0_read_illegal_T_254 ;  
   wire _io_decode_0_read_illegal_T_255 ;  
   wire _io_decode_0_read_illegal_T_256 ;  
   wire _io_decode_0_read_illegal_T_257 ;  
   wire _io_decode_0_read_illegal_T_258 ;  
   wire _io_decode_0_read_illegal_T_259 ;  
   wire _io_decode_0_read_illegal_T_260 ;  
   wire _io_decode_0_read_illegal_T_261 ;  
   wire _io_decode_0_read_illegal_T_262 ;  
   wire _io_decode_0_read_illegal_T_263 ;  
   wire _io_decode_0_read_illegal_T_264 ;  
   wire _io_decode_0_read_illegal_T_265 ;  
   wire _io_decode_0_read_illegal_T_266 ;  
   wire _io_decode_0_read_illegal_T_267 ;  
   wire _io_decode_0_read_illegal_T_268 ;  
   wire _io_decode_0_read_illegal_T_269 ;  
   wire _io_decode_0_read_illegal_T_270 ;  
   wire _io_decode_0_read_illegal_T_271 ;  
   wire _io_decode_0_read_illegal_T_272 ;  
   wire _io_decode_0_read_illegal_T_273 ;  
   wire _io_decode_0_read_illegal_T_274 ;  
   wire _io_decode_0_read_illegal_T_275 ;  
   wire _io_decode_0_read_illegal_T_276 ;  
   wire _io_decode_0_read_illegal_T_277 ;  
   wire _io_decode_0_read_illegal_T_278 ;  
   wire _io_decode_0_read_illegal_T_279 ;  
   wire _io_decode_0_read_illegal_T_280 ;  
   wire _io_decode_0_read_illegal_T_281 ;  
   wire _io_decode_0_read_illegal_T_282 ;  
   wire _io_decode_0_read_illegal_T_283 ;  
   wire _io_decode_0_read_illegal_T_284 ;  
   wire _io_decode_0_read_illegal_T_285 ;  
   wire _io_decode_0_read_illegal_T_286 ;  
   wire _io_decode_0_read_illegal_T_287 ;  
   wire _io_decode_0_read_illegal_T_288 ;  
   wire _io_decode_0_read_illegal_T_289 ;  
   wire _io_decode_0_read_illegal_T_290 ;  
   wire _io_decode_0_read_illegal_T_291 ;  
   wire _io_decode_0_read_illegal_T_292 ;  
   wire _io_decode_0_read_illegal_T_293 ;  
   wire _io_decode_0_read_illegal_T_294 ;  
   wire _io_decode_0_read_illegal_T_296 ;  
   wire _io_decode_0_read_illegal_T_299 ;  
   wire _io_decode_0_read_illegal_T_300 ;  
   wire _io_decode_0_read_illegal_T_301 ;  
   wire _io_decode_0_read_illegal_T_302 ;  
   wire _io_decode_0_read_illegal_T_303 ;  
   wire _io_decode_0_read_illegal_T_304 ;  
   wire _io_decode_0_read_illegal_T_305 ;  
   wire _io_decode_0_read_illegal_T_306 ;  
   wire _io_decode_0_read_illegal_T_307 ;  
   wire _io_decode_0_read_illegal_T_309 ;  
   wire _io_decode_0_read_illegal_T_310 ;  
   wire [11:0] _io_decode_0_read_illegal_T_311 ;  
   wire _io_decode_0_read_illegal_T_312 ;  
   wire _io_decode_0_read_illegal_T_316 ;  
   wire _io_decode_0_read_illegal_T_317 ;  
   wire _io_decode_0_read_illegal_T_320 ;  
   wire _io_decode_0_write_flush_T ;  
   wire _io_decode_0_write_flush_T_1 ;  
   wire _io_decode_0_write_flush_T_2 ;  
   wire _io_decode_0_write_flush_T_3 ;  
   wire _io_decode_0_write_flush_T_4 ;  
   wire _io_decode_0_write_flush_T_5 ;  
   wire _io_decode_0_write_flush_T_6 ;  
   wire _io_decode_0_system_illegal_T_3 ;  
   wire _io_decode_0_system_illegal_T_4 ;  
   wire _io_decode_0_system_illegal_T_6 ;  
   wire _io_decode_0_system_illegal_T_7 ;  
   wire _io_decode_0_system_illegal_T_9 ;  
   wire _io_decode_0_system_illegal_T_11 ;  
   wire _io_decode_0_system_illegal_T_13 ;  
   wire _io_decode_0_system_illegal_T_14 ;  
   wire _io_decode_0_system_illegal_T_16 ;  
   wire [11:0] _debugTVec_T ;  
   wire [11:0] debugTVec ;  
   wire [63:0] notDebugTVec_base ;  
   wire [7:0] notDebugTVec_interruptVec_lo ;  
   wire [55:0] notDebugTVec_interruptVec_hi ;  
   wire [63:0] notDebugTVec_interruptVec ;  
   wire _notDebugTVec_doVector_T_2 ;  
   wire _notDebugTVec_doVector_T_4 ;  
   wire notDebugTVec_doVector ;  
   wire [63:0] _notDebugTVec_T_1 ;  
   wire [63:0] notDebugTVec ;  
   wire [63:0] tvec ;  
   wire _io_status_sd_T ;  
   wire _io_status_sd_T_1 ;  
   wire _io_status_sd_T_2 ;  
   wire _io_status_sd_T_3 ;  
   wire _io_status_dprv_x87_T_1 ;  
   reg [1:0] io_status_dprv_REG ;  
   reg [31:0] _RAND_114 ;  
   wire [1:0] _T_244 ;  
   wire [1:0] _T_246 ;  
   wire [2:0] _T_248 ;  
   wire _T_250 ;  
   wire _T_252 ;  
   wire _T_255 ;  
   wire _T_257 ;  
   wire _GEN_48 ;  
   wire _T_258 ;  
   wire _T_259 ;  
   wire _T_260 ;  
   wire _T_262 ;  
   wire _GEN_50 ;  
   wire _T_272 ;  
   wire _T_274 ;  
   wire [39:0] _epc_T_1 ;  
   wire [39:0] epc ;  
   wire [1:0] _reg_dcsr_cause_T ;  
   wire [1:0] _reg_dcsr_cause_T_1 ;  
   wire _GEN_52 ;  
   wire [39:0] _GEN_53 ;  
   wire [39:0] _GEN_63 ;  
   wire _GEN_67 ;  
   wire [1:0] _GEN_68 ;  
   wire [39:0] _GEN_71 ;  
   wire _GEN_74 ;  
   wire [1:0] _GEN_75 ;  
   wire _GEN_76 ;  
   wire [39:0] _GEN_97 ;  
   wire [39:0] _GEN_106 ;  
   wire _GEN_110 ;  
   wire [1:0] _GEN_111 ;  
   wire [39:0] _GEN_113 ;  
   wire _GEN_116 ;  
   wire [1:0] _GEN_117 ;  
   wire _GEN_118 ;  
   wire [39:0] _GEN_120 ;  
   wire [39:0] _GEN_129 ;  
   wire _GEN_133 ;  
   wire [1:0] _GEN_134 ;  
   wire [39:0] _GEN_136 ;  
   wire _GEN_139 ;  
   wire [1:0] _GEN_140 ;  
   wire _GEN_141 ;  
   wire [39:0] _GEN_151 ;  
   wire _GEN_158 ;  
   wire [1:0] _GEN_159 ;  
   wire [39:0] _GEN_161 ;  
   wire _T_412 ;  
   wire [1:0] _GEN_171 ;  
   wire [63:0] _GEN_172 ;  
   reg io_status_cease_r ;  
   reg [31:0] _RAND_115 ;  
   wire _GEN_181 ;  
   wire [63:0] _io_rw_rdata_T_1 ;  
   wire [63:0] _io_rw_rdata_T_2 ;  
   wire [63:0] _io_rw_rdata_T_4 ;  
   wire [63:0] _io_rw_rdata_T_5 ;  
   wire [63:0] _io_rw_rdata_T_6 ;  
   wire [15:0] _io_rw_rdata_T_7 ;  
   wire [63:0] _io_rw_rdata_T_8 ;  
   wire [63:0] _io_rw_rdata_T_9 ;  
   wire [63:0] _io_rw_rdata_T_10 ;  
   wire [63:0] _io_rw_rdata_T_11 ;  
   wire [63:0] _io_rw_rdata_T_12 ;  
   wire _io_rw_rdata_T_13 ;  
   wire [31:0] _io_rw_rdata_T_14 ;  
   wire [63:0] _io_rw_rdata_T_15 ;  
   wire [63:0] _io_rw_rdata_T_16 ;  
   wire [4:0] _io_rw_rdata_T_17 ;  
   wire [2:0] _io_rw_rdata_T_18 ;  
   wire [7:0] _io_rw_rdata_T_19 ;  
   wire [2:0] _io_rw_rdata_T_20 ;  
   wire [63:0] _io_rw_rdata_T_21 ;  
   wire [63:0] _io_rw_rdata_T_22 ;  
   wire [31:0] _io_rw_rdata_T_110 ;  
   wire [63:0] _io_rw_rdata_T_111 ;  
   wire [63:0] _io_rw_rdata_T_112 ;  
   wire [63:0] _io_rw_rdata_T_113 ;  
   wire [63:0] _io_rw_rdata_T_114 ;  
   wire [63:0] _io_rw_rdata_T_115 ;  
   wire [63:0] _io_rw_rdata_T_116 ;  
   wire [63:0] _io_rw_rdata_T_117 ;  
   wire [63:0] _io_rw_rdata_T_118 ;  
   wire [63:0] _io_rw_rdata_T_119 ;  
   wire [63:0] _io_rw_rdata_T_120 ;  
   wire [63:0] _io_rw_rdata_T_121 ;  
   wire [31:0] _io_rw_rdata_T_122 ;  
   wire [63:0] _io_rw_rdata_T_123 ;  
   wire [63:0] _io_rw_rdata_T_124 ;  
   wire [63:0] _io_rw_rdata_T_125 ;  
   wire [29:0] _io_rw_rdata_T_127 ;  
   wire [29:0] _io_rw_rdata_T_128 ;  
   wire [29:0] _io_rw_rdata_T_129 ;  
   wire [29:0] _io_rw_rdata_T_130 ;  
   wire [29:0] _io_rw_rdata_T_131 ;  
   wire [29:0] _io_rw_rdata_T_132 ;  
   wire [29:0] _io_rw_rdata_T_133 ;  
   wire [29:0] _io_rw_rdata_T_134 ;  
   wire [63:0] _io_rw_rdata_T_143 ;  
   wire [63:0] _io_rw_rdata_T_144 ;  
   wire [63:0] _io_rw_rdata_T_146 ;  
   wire [63:0] _io_rw_rdata_T_148 ;  
   wire [63:0] _io_rw_rdata_T_150 ;  
   wire [63:0] _io_rw_rdata_T_151 ;  
   wire [63:0] _io_rw_rdata_T_152 ;  
   wire [63:0] _GEN_565 ;  
   wire [63:0] _io_rw_rdata_T_153 ;  
   wire [63:0] _io_rw_rdata_T_154 ;  
   wire [63:0] _io_rw_rdata_T_155 ;  
   wire [63:0] _io_rw_rdata_T_156 ;  
   wire [63:0] _io_rw_rdata_T_157 ;  
   wire [63:0] _io_rw_rdata_T_158 ;  
   wire [63:0] _GEN_566 ;  
   wire [63:0] _io_rw_rdata_T_159 ;  
   wire [63:0] _GEN_567 ;  
   wire [63:0] _io_rw_rdata_T_160 ;  
   wire [63:0] _io_rw_rdata_T_161 ;  
   wire [63:0] _io_rw_rdata_T_162 ;  
   wire [63:0] _GEN_568 ;  
   wire [63:0] _io_rw_rdata_T_163 ;  
   wire [63:0] _GEN_569 ;  
   wire [63:0] _io_rw_rdata_T_164 ;  
   wire [63:0] _GEN_570 ;  
   wire [63:0] _io_rw_rdata_T_165 ;  
   wire [63:0] _GEN_571 ;  
   wire [63:0] _io_rw_rdata_T_166 ;  
   wire [63:0] _io_rw_rdata_T_167 ;  
   wire [63:0] _io_rw_rdata_T_168 ;  
   wire [63:0] _GEN_572 ;  
   wire [63:0] _io_rw_rdata_T_256 ;  
   wire [63:0] _io_rw_rdata_T_257 ;  
   wire [63:0] _io_rw_rdata_T_258 ;  
   wire [63:0] _io_rw_rdata_T_259 ;  
   wire [63:0] _io_rw_rdata_T_260 ;  
   wire [63:0] _io_rw_rdata_T_261 ;  
   wire [63:0] _io_rw_rdata_T_262 ;  
   wire [63:0] _io_rw_rdata_T_263 ;  
   wire [63:0] _io_rw_rdata_T_264 ;  
   wire [63:0] _io_rw_rdata_T_265 ;  
   wire [63:0] _io_rw_rdata_T_266 ;  
   wire [63:0] _io_rw_rdata_T_267 ;  
   wire [63:0] _GEN_573 ;  
   wire [63:0] _io_rw_rdata_T_268 ;  
   wire [63:0] _io_rw_rdata_T_269 ;  
   wire [63:0] _io_rw_rdata_T_270 ;  
   wire [63:0] _io_rw_rdata_T_271 ;  
   wire [63:0] _GEN_574 ;  
   wire [63:0] _io_rw_rdata_T_273 ;  
   wire [63:0] _GEN_575 ;  
   wire [63:0] _io_rw_rdata_T_274 ;  
   wire [63:0] _GEN_576 ;  
   wire [63:0] _io_rw_rdata_T_275 ;  
   wire [63:0] _GEN_577 ;  
   wire [63:0] _io_rw_rdata_T_276 ;  
   wire [63:0] _GEN_578 ;  
   wire [63:0] _io_rw_rdata_T_277 ;  
   wire [63:0] _GEN_579 ;  
   wire [63:0] _io_rw_rdata_T_278 ;  
   wire [63:0] _GEN_580 ;  
   wire [63:0] _io_rw_rdata_T_279 ;  
   wire [63:0] _GEN_581 ;  
   wire [63:0] _io_rw_rdata_T_280 ;  
   wire [63:0] _io_rw_rdata_T_289 ;  
   wire [63:0] _io_rw_rdata_T_290 ;  
   wire _T_416 ;  
   wire _T_417 ;  
   wire _T_418 ;  
   wire [4:0] _lo_T ;  
   wire [4:0] _GEN_182 ;  
   wire _csr_wen_T_3 ;  
   wire csr_wen ;  
   wire [102:0] _new_mstatus_WIRE ;  
   wire new_mstatus_sie ;  
   wire new_mstatus_mie ;  
   wire new_mstatus_spie ;  
   wire new_mstatus_mpie ;  
   wire new_mstatus_spp ;  
   wire [1:0] new_mstatus_mpp ;  
   wire [1:0] new_mstatus_fs ;  
   wire new_mstatus_mprv ;  
   wire new_mstatus_sum ;  
   wire new_mstatus_mxr ;  
   wire new_mstatus_tvm ;  
   wire new_mstatus_tw ;  
   wire new_mstatus_tsr ;  
   wire _reg_mstatus_mpp_T_2 ;  
   wire _reg_mstatus_fs_T ;  
   wire [1:0] _GEN_188 ;  
   wire f ;  
   wire _T_1834 ;  
   wire [3:0] _reg_misa_T_2 ;  
   wire [63:0] _GEN_582 ;  
   wire [63:0] _reg_misa_T_3 ;  
   wire [63:0] _reg_misa_T_5 ;  
   wire [63:0] _reg_misa_T_7 ;  
   wire [63:0] _reg_misa_T_8 ;  
   wire [15:0] _new_mip_T ;  
   wire [15:0] _new_mip_T_2 ;  
   wire [63:0] _GEN_583 ;  
   wire [63:0] _new_mip_T_3 ;  
   wire [63:0] _new_mip_T_8 ;  
   wire new_mip_ssip ;  
   wire new_mip_stip ;  
   wire new_mip_seip ;  
   wire [63:0] _reg_mie_T ;  
   wire [63:0] _reg_mepc_T_1 ;  
   wire [63:0] _GEN_204 ;  
   wire [63:0] _GEN_206 ;  
   wire [63:0] _reg_mcause_T ;  
   wire [63:0] _reg_mcountinhibit_T_1 ;  
   wire [63:0] _GEN_209 ;  
   wire [63:0] _GEN_210 ;  
   wire [63:0] _GEN_212 ;  
   wire [63:0] _GEN_215 ;  
   wire [63:0] _GEN_217 ;  
   wire [63:0] _GEN_219 ;  
   wire [63:0] _GEN_220 ;  
   wire [1:0] new_dcsr_prv ;  
   wire new_dcsr_step ;  
   wire new_dcsr_ebreaku ;  
   wire new_dcsr_ebreaks ;  
   wire new_dcsr_ebreakm ;  
   wire _reg_dcsr_prv_T ;  
   wire [63:0] _GEN_226 ;  
   wire [1:0] _GEN_230 ;  
   wire [63:0] _new_sip_T_1 ;  
   wire [63:0] _new_sip_T_2 ;  
   wire [63:0] _new_sip_T_3 ;  
   wire new_sip_ssip ;  
   wire [43:0] new_satp_ppn ;  
   wire [3:0] new_satp_mode ;  
   wire _T_1837 ;  
   wire _T_1838 ;  
   wire _T_1839 ;  
   wire [3:0] _reg_satp_mode_T ;  
   wire [63:0] _reg_mie_T_2 ;  
   wire [63:0] _reg_mie_T_4 ;  
   wire [63:0] _GEN_242 ;  
   wire [63:0] _GEN_243 ;  
   wire [63:0] _reg_scause_T ;  
   wire [63:0] _GEN_248 ;  
   wire [63:0] _GEN_249 ;  
   wire _T_1842 ;  
   wire [63:0] _GEN_251 ;  
   wire [63:0] _newBPC_T_2 ;  
   wire [63:0] _newBPC_T_3 ;  
   wire [63:0] _newBPC_T_8 ;  
   wire newBPC_action ;  
   wire newBPC_dmode ;  
   wire dMode ;  
   wire _GEN_252 ;  
   wire [63:0] _GEN_268 ;  
   wire _T_1853 ;  
   wire newCfg_r ;  
   wire newCfg_w ;  
   wire newCfg_x ;  
   wire [1:0] newCfg_a ;  
   wire newCfg_l ;  
   wire _reg_pmp_0_cfg_w_T ;  
   wire _T_1857 ;  
   wire _T_1858 ;  
   wire _T_1859 ;  
   wire _T_1861 ;  
   wire [63:0] _GEN_323 ;  
   wire _T_1863 ;  
   wire newCfg_1_r ;  
   wire newCfg_1_w ;  
   wire newCfg_1_x ;  
   wire [1:0] newCfg_1_a ;  
   wire newCfg_1_l ;  
   wire _reg_pmp_1_cfg_w_T ;  
   wire _T_1867 ;  
   wire _T_1868 ;  
   wire _T_1869 ;  
   wire _T_1871 ;  
   wire [63:0] _GEN_330 ;  
   wire _T_1873 ;  
   wire newCfg_2_r ;  
   wire newCfg_2_w ;  
   wire newCfg_2_x ;  
   wire [1:0] newCfg_2_a ;  
   wire newCfg_2_l ;  
   wire _reg_pmp_2_cfg_w_T ;  
   wire _T_1877 ;  
   wire _T_1878 ;  
   wire _T_1879 ;  
   wire _T_1881 ;  
   wire [63:0] _GEN_337 ;  
   wire _T_1883 ;  
   wire newCfg_3_r ;  
   wire newCfg_3_w ;  
   wire newCfg_3_x ;  
   wire [1:0] newCfg_3_a ;  
   wire newCfg_3_l ;  
   wire _reg_pmp_3_cfg_w_T ;  
   wire _T_1887 ;  
   wire _T_1888 ;  
   wire _T_1889 ;  
   wire _T_1891 ;  
   wire [63:0] _GEN_344 ;  
   wire _T_1893 ;  
   wire newCfg_4_r ;  
   wire newCfg_4_w ;  
   wire newCfg_4_x ;  
   wire [1:0] newCfg_4_a ;  
   wire newCfg_4_l ;  
   wire _reg_pmp_4_cfg_w_T ;  
   wire _T_1897 ;  
   wire _T_1898 ;  
   wire _T_1899 ;  
   wire _T_1901 ;  
   wire [63:0] _GEN_351 ;  
   wire _T_1903 ;  
   wire newCfg_5_r ;  
   wire newCfg_5_w ;  
   wire newCfg_5_x ;  
   wire [1:0] newCfg_5_a ;  
   wire newCfg_5_l ;  
   wire _reg_pmp_5_cfg_w_T ;  
   wire _T_1907 ;  
   wire _T_1908 ;  
   wire _T_1909 ;  
   wire _T_1911 ;  
   wire [63:0] _GEN_358 ;  
   wire _T_1913 ;  
   wire newCfg_6_r ;  
   wire newCfg_6_w ;  
   wire newCfg_6_x ;  
   wire [1:0] newCfg_6_a ;  
   wire newCfg_6_l ;  
   wire _reg_pmp_6_cfg_w_T ;  
   wire _T_1917 ;  
   wire _T_1918 ;  
   wire _T_1919 ;  
   wire _T_1921 ;  
   wire [63:0] _GEN_365 ;  
   wire _T_1923 ;  
   wire newCfg_7_r ;  
   wire newCfg_7_w ;  
   wire newCfg_7_x ;  
   wire [1:0] newCfg_7_a ;  
   wire newCfg_7_l ;  
   wire _reg_pmp_7_cfg_w_T ;  
   wire _T_1929 ;  
   wire _T_1931 ;  
   wire [63:0] _GEN_372 ;  
   wire [63:0] _reg_custom_0_T ;  
   wire [63:0] _reg_custom_0_T_2 ;  
   wire [63:0] _reg_custom_0_T_3 ;  
   wire [1:0] _GEN_385 ;  
   wire [63:0] _GEN_400 ;  
   wire [63:0] _GEN_402 ;  
   wire [63:0] _GEN_405 ;  
   wire [63:0] _GEN_406 ;  
   wire [63:0] _GEN_408 ;  
   wire [63:0] _GEN_411 ;  
   wire [63:0] _GEN_412 ;  
   wire [63:0] _GEN_418 ;  
   wire [63:0] _GEN_423 ;  
   wire [63:0] _GEN_424 ;  
   wire [63:0] _GEN_429 ;  
   wire [63:0] _GEN_430 ;  
   wire [63:0] _GEN_432 ;  
   wire [63:0] _GEN_470 ;  
   wire [63:0] _GEN_477 ;  
   wire [63:0] _GEN_484 ;  
   wire [63:0] _GEN_491 ;  
   wire [63:0] _GEN_498 ;  
   wire [63:0] _GEN_505 ;  
   wire [63:0] _GEN_512 ;  
   wire [63:0] _GEN_519 ;  
   wire _io_trace_0_valid_T ;  
   reg [19:0] CSRFile_state ;  
   reg [31:0] _RAND_116 ;  
   reg CSRFile_cov[0:1048575] ;  
   reg [31:0] _RAND_117 ;  
   wire CSRFile_cov_read_data ;  
   wire [19:0] CSRFile_cov_read_addr ;  
   wire CSRFile_cov_write_data ;  
   wire [19:0] CSRFile_cov_write_addr ;  
   wire CSRFile_cov_write_mask ;  
   wire CSRFile_cov_write_en ;  
   reg [29:0] CSRFile_covSum ;  
   reg [31:0] _RAND_118 ;  
   wire [19:0] reg_pmp_5_cfg_l_shl ;  
   wire [19:0] reg_pmp_5_cfg_l_pad ;  
   wire [1:0] reg_debug_shl ;  
   wire [19:0] reg_debug_pad ;  
   wire [16:0] reg_mstatus_sie_shl ;  
   wire [19:0] reg_mstatus_sie_pad ;  
   wire [14:0] reg_dcsr_prv_shl ;  
   wire [19:0] reg_dcsr_prv_pad ;  
   wire [17:0] reg_mcountinhibit_shl ;  
   wire [19:0] reg_mcountinhibit_pad ;  
   wire [2:0] reg_unmie_shl ;  
   wire [19:0] reg_unmie_pad ;  
   wire [14:0] reg_pmp_7_cfg_a_shl ;  
   wire [19:0] reg_pmp_7_cfg_a_pad ;  
   wire [1:0] reg_mstatus_mpp_shl ;  
   wire [19:0] reg_mstatus_mpp_pad ;  
   wire [6:0] reg_pmp_2_cfg_l_shl ;  
   wire [19:0] reg_pmp_2_cfg_l_pad ;  
   wire [18:0] reg_pmp_1_cfg_l_shl ;  
   wire [19:0] reg_pmp_1_cfg_l_pad ;  
   wire [9:0] reg_mip_seip_shl ;  
   wire [19:0] reg_mip_seip_pad ;  
   wire [1:0] reg_rnmie_shl ;  
   wire [19:0] reg_rnmie_pad ;  
   wire [10:0] reg_mip_ssip_shl ;  
   wire [19:0] reg_mip_ssip_pad ;  
   wire [2:0] reg_bp_0_control_dmode_shl ;  
   wire [19:0] reg_bp_0_control_dmode_pad ;  
   wire [11:0] reg_pmp_4_cfg_l_shl ;  
   wire [19:0] reg_pmp_4_cfg_l_pad ;  
   wire [1:0] reg_dcsr_ebreaks_shl ;  
   wire [19:0] reg_dcsr_ebreaks_pad ;  
   wire [13:0] reg_pmp_6_cfg_l_shl ;  
   wire [19:0] reg_pmp_6_cfg_l_pad ;  
   wire [3:0] reg_mstatus_prv_shl ;  
   wire [19:0] reg_mstatus_prv_pad ;  
   wire [8:0] reg_dcsr_ebreakm_shl ;  
   wire [19:0] reg_dcsr_ebreakm_pad ;  
   wire reg_pmp_7_cfg_l_shl ;  
   wire [19:0] reg_pmp_7_cfg_l_pad ;  
   wire [18:0] reg_pmp_0_cfg_l_shl ;  
   wire [19:0] reg_pmp_0_cfg_l_pad ;  
   wire [1:0] reg_pmp_3_cfg_l_shl ;  
   wire [19:0] reg_pmp_3_cfg_l_pad ;  
   wire [13:0] reg_mstatus_spp_shl ;  
   wire [19:0] reg_mstatus_spp_pad ;  
   wire [12:0] reg_mip_stip_shl ;  
   wire [19:0] reg_mip_stip_pad ;  
   wire [13:0] reg_dcsr_ebreaku_shl ;  
   wire [19:0] reg_dcsr_ebreaku_pad ;  
   wire reg_mstatus_mprv_shl ;  
   wire [19:0] reg_mstatus_mprv_pad ;  
   wire [13:0] reg_singleStepped_shl ;  
   wire [19:0] reg_singleStepped_pad ;  
   wire [11:0] reg_mstatus_mie_shl ;  
   wire [19:0] reg_mstatus_mie_pad ;  
   wire [19:0] CSRFile_xor16 ;  
   wire [19:0] CSRFile_xor7 ;  
   wire [19:0] CSRFile_xor17 ;  
   wire [19:0] CSRFile_xor18 ;  
   wire [19:0] CSRFile_xor8 ;  
   wire [19:0] CSRFile_xor3 ;  
   wire [19:0] CSRFile_xor20 ;  
   wire [19:0] CSRFile_xor9 ;  
   wire [19:0] CSRFile_xor21 ;  
   wire [19:0] CSRFile_xor22 ;  
   wire [19:0] CSRFile_xor10 ;  
   wire [19:0] CSRFile_xor4 ;  
   wire [19:0] CSRFile_xor1 ;  
   wire [19:0] CSRFile_xor24 ;  
   wire [19:0] CSRFile_xor11 ;  
   wire [19:0] CSRFile_xor25 ;  
   wire [19:0] CSRFile_xor26 ;  
   wire [19:0] CSRFile_xor12 ;  
   wire [19:0] CSRFile_xor5 ;  
   wire [19:0] CSRFile_xor28 ;  
   wire [19:0] CSRFile_xor13 ;  
   wire [19:0] CSRFile_xor29 ;  
   wire [19:0] CSRFile_xor30 ;  
   wire [19:0] CSRFile_xor14 ;  
   wire [19:0] CSRFile_xor6 ;  
   wire [19:0] CSRFile_xor2 ;  
   wire [19:0] CSRFile_xor0 ;  
   wire stopEn0 ;  
   wire stopEn1 ;  
   wire CSRFile_or0 ;  
   reg CSRFile_metaAssert ;  
   reg [31:0] _RAND_119 ;  
  assign system_insn=io_rw_cmd==3'h4; 
  assign _T_192={io_rw_addr,20'h0}; 
  assign _T_199=_T_192&32'h12400000; 
  assign _T_200=_T_199==32'h10000000; 
  assign _T_201=_T_192&32'h40000000; 
  assign _T_202=_T_201==32'h40000000; 
  assign _T_204=_T_200|_T_202; 
  assign insn_ret=system_insn&_T_204; 
  assign _T_406=io_rw_addr[10]&io_rw_addr[7]; 
  assign _GEN_149=_T_406 ? reg_dcsr_prv:reg_mstatus_mpp; 
  assign ret_prv=io_rw_addr[9] ? _GEN_149:{1'b0,reg_mstatus_spp}; 
  assign _T_193=_T_192&32'h10100000; 
  assign _T_194=_T_193==32'h0; 
  assign insn_call=system_insn&_T_194; 
  assign _T_197=_T_193==32'h100000; 
  assign insn_break=system_insn&_T_197; 
  assign _exception_T=insn_call|insn_break; 
  assign exception=_exception_T|io_exception; 
  assign _GEN_20={2'b0,reg_mstatus_prv}; 
  assign _cause_T_1=_GEN_20+4'h8; 
  assign _cause_T_2=insn_break ? 64'h3:io_cause; 
  assign cause=insn_call ? {60'b0,_cause_T_1}:_cause_T_2; 
  assign cause_lsbs=cause[7:0]; 
  assign _causeIsDebugInt_T_1=cause_lsbs==8'he; 
  assign causeIsDebugInt=cause[63]&_causeIsDebugInt_T_1; 
  assign _trapToDebug_T=reg_singleStepped|causeIsDebugInt; 
  assign causeIsDebugTrigger=~cause[63]&_causeIsDebugInt_T_1; 
  assign _trapToDebug_T_1=_trapToDebug_T|causeIsDebugTrigger; 
  assign _causeIsDebugBreak_T_2=~cause[63]&insn_break; 
  assign _causeIsDebugBreak_T_3={reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku}; 
  assign _causeIsDebugBreak_T_4=_causeIsDebugBreak_T_3>>reg_mstatus_prv; 
  assign causeIsDebugBreak=_causeIsDebugBreak_T_2&_causeIsDebugBreak_T_4[0]; 
  assign _trapToDebug_T_2=_trapToDebug_T_1|causeIsDebugBreak; 
  assign trapToDebug=_trapToDebug_T_2|reg_debug; 
  assign _GEN_56=reg_debug ? reg_mstatus_prv:2'h3; 
  assign _delegate_T=reg_mstatus_prv<=2'h1; 
  assign read_mideleg=reg_mideleg&64'h222; 
  assign _delegate_T_3=read_mideleg>>cause_lsbs; 
  assign read_medeleg=reg_medeleg&64'hb15d; 
  assign _delegate_T_5=read_medeleg>>cause_lsbs; 
  assign _delegate_T_7=cause[63] ? _delegate_T_3[0]:_delegate_T_5[0]; 
  assign delegate=_delegate_T&_delegate_T_7; 
  assign nmie=reg_rnmie&reg_unmie; 
  assign _T_279=delegate&nmie; 
  assign _GEN_70=_T_279 ? 2'h1:2'h3; 
  assign _GEN_100=trapToDebug ? _GEN_56:_GEN_70; 
  assign _GEN_123=exception ? _GEN_100:reg_mstatus_prv; 
  assign new_prv=insn_ret ? ret_prv:_GEN_123; 
  assign _reg_mstatus_prv_T=new_prv==2'h2; 
  assign read_mcounteren=reg_mcounteren&32'h7; 
  assign read_scounteren=reg_scounteren&32'h7; 
  assign x67=reg_mcountinhibit[2]; 
  assign _GEN_23={5'b0,io_retire}; 
  assign nextSmall=value_lo+_GEN_23; 
  assign _GEN_0=x67 ? {1'b0,value_lo}:nextSmall; 
  assign _large_T_2=nextSmall[6]&~x67; 
  assign _large_r_T_1=value_hi+58'h1; 
  assign value={value_hi,value_lo}; 
  assign nextSmall_1=value_lo_1+_GEN_23; 
  assign _GEN_2=reg_mcountinhibit[0] ? {1'b0,value_lo_1}:nextSmall_1; 
  assign _large_T_5=nextSmall_1[6]&~reg_mcountinhibit[0]; 
  assign _large_r_T_3=value_hi_1+58'h1; 
  assign value_1={value_hi_1,value_lo_1}; 
  assign mip_seip=reg_mip_seip|io_interrupts_seip; 
  assign read_mip_lo={io_interrupts_mtip,1'h0,reg_mip_stip,1'h0,io_interrupts_msip,1'h0,reg_mip_ssip,1'h0}; 
  assign _read_mip_T={4'h0,io_interrupts_meip,1'h0,mip_seip,1'h0,read_mip_lo}; 
  assign read_mip=_read_mip_T&16'haaa; 
   reg [15:0] reg_mip ;  
  assign reg_mip=read_mip; 
  assign _GEN_45={48'b0,read_mip}; 
  assign pending_interrupts=_GEN_45&reg_mie; 
  assign d_interrupts={io_interrupts_debug,14'h0}; 
  assign _m_interrupts_T_1=_delegate_T|reg_mstatus_mie; 
  assign _m_interrupts_T_2=nmie&_m_interrupts_T_1; 
  assign _m_interrupts_T_4=~pending_interrupts|read_mideleg; 
  assign m_interrupts=_m_interrupts_T_2 ? ~_m_interrupts_T_4:64'h0; 
  assign _s_interrupts_T=reg_mstatus_prv<2'h1; 
  assign _s_interrupts_T_1=reg_mstatus_prv==2'h1; 
  assign _s_interrupts_T_2=_s_interrupts_T_1&reg_mstatus_sie; 
  assign _s_interrupts_T_3=_s_interrupts_T|_s_interrupts_T_2; 
  assign _s_interrupts_T_4=nmie&_s_interrupts_T_3; 
  assign _s_interrupts_T_5=pending_interrupts&read_mideleg; 
  assign s_interrupts=_s_interrupts_T_4 ? _s_interrupts_T_5:64'h0; 
  assign _any_T_38=d_interrupts[14]|d_interrupts[13]; 
  assign _any_T_39=_any_T_38|d_interrupts[12]; 
  assign _any_T_40=_any_T_39|d_interrupts[11]; 
  assign _any_T_41=_any_T_40|d_interrupts[3]; 
  assign _any_T_42=_any_T_41|d_interrupts[7]; 
  assign _any_T_43=_any_T_42|d_interrupts[9]; 
  assign _any_T_44=_any_T_43|d_interrupts[1]; 
  assign _any_T_45=_any_T_44|d_interrupts[5]; 
  assign _any_T_46=_any_T_45|d_interrupts[8]; 
  assign _any_T_47=_any_T_46|d_interrupts[0]; 
  assign _any_T_48=_any_T_47|d_interrupts[4]; 
  assign _any_T_50=_any_T_48|m_interrupts[15]; 
  assign _any_T_51=_any_T_50|m_interrupts[14]; 
  assign _any_T_52=_any_T_51|m_interrupts[13]; 
  assign _any_T_53=_any_T_52|m_interrupts[12]; 
  assign _any_T_54=_any_T_53|m_interrupts[11]; 
  assign _any_T_55=_any_T_54|m_interrupts[3]; 
  assign _any_T_56=_any_T_55|m_interrupts[7]; 
  assign _any_T_57=_any_T_56|m_interrupts[9]; 
  assign _any_T_58=_any_T_57|m_interrupts[1]; 
  assign _any_T_59=_any_T_58|m_interrupts[5]; 
  assign _any_T_60=_any_T_59|m_interrupts[8]; 
  assign _any_T_61=_any_T_60|m_interrupts[0]; 
  assign _any_T_62=_any_T_61|m_interrupts[4]; 
  assign _any_T_63=_any_T_62|s_interrupts[15]; 
  assign _any_T_64=_any_T_63|s_interrupts[14]; 
  assign _any_T_65=_any_T_64|s_interrupts[13]; 
  assign _any_T_66=_any_T_65|s_interrupts[12]; 
  assign _any_T_67=_any_T_66|s_interrupts[11]; 
  assign _any_T_68=_any_T_67|s_interrupts[3]; 
  assign _any_T_69=_any_T_68|s_interrupts[7]; 
  assign _any_T_70=_any_T_69|s_interrupts[9]; 
  assign _any_T_71=_any_T_70|s_interrupts[1]; 
  assign _any_T_72=_any_T_71|s_interrupts[5]; 
  assign _any_T_73=_any_T_72|s_interrupts[8]; 
  assign _any_T_74=_any_T_73|s_interrupts[0]; 
  assign anyInterrupt=_any_T_74|s_interrupts[4]; 
  assign _which_T_38=s_interrupts[0] ? 3'h0:3'h4; 
  assign _which_T_39=s_interrupts[8] ? 4'h8:{1'b0,_which_T_38}; 
  assign _which_T_40=s_interrupts[5] ? 4'h5:_which_T_39; 
  assign _which_T_41=s_interrupts[1] ? 4'h1:_which_T_40; 
  assign _which_T_42=s_interrupts[9] ? 4'h9:_which_T_41; 
  assign _which_T_43=s_interrupts[7] ? 4'h7:_which_T_42; 
  assign _which_T_44=s_interrupts[3] ? 4'h3:_which_T_43; 
  assign _which_T_45=s_interrupts[11] ? 4'hb:_which_T_44; 
  assign _which_T_46=s_interrupts[12] ? 4'hc:_which_T_45; 
  assign _which_T_47=s_interrupts[13] ? 4'hd:_which_T_46; 
  assign _which_T_48=s_interrupts[14] ? 4'he:_which_T_47; 
  assign _which_T_49=s_interrupts[15] ? 4'hf:_which_T_48; 
  assign _which_T_50=m_interrupts[4] ? 4'h4:_which_T_49; 
  assign _which_T_51=m_interrupts[0] ? 4'h0:_which_T_50; 
  assign _which_T_52=m_interrupts[8] ? 4'h8:_which_T_51; 
  assign _which_T_53=m_interrupts[5] ? 4'h5:_which_T_52; 
  assign _which_T_54=m_interrupts[1] ? 4'h1:_which_T_53; 
  assign _which_T_55=m_interrupts[9] ? 4'h9:_which_T_54; 
  assign _which_T_56=m_interrupts[7] ? 4'h7:_which_T_55; 
  assign _which_T_57=m_interrupts[3] ? 4'h3:_which_T_56; 
  assign _which_T_58=m_interrupts[11] ? 4'hb:_which_T_57; 
  assign _which_T_59=m_interrupts[12] ? 4'hc:_which_T_58; 
  assign _which_T_60=m_interrupts[13] ? 4'hd:_which_T_59; 
  assign _which_T_61=m_interrupts[14] ? 4'he:_which_T_60; 
  assign _which_T_62=m_interrupts[15] ? 4'hf:_which_T_61; 
  assign _which_T_64=d_interrupts[4] ? 4'h4:_which_T_62; 
  assign _which_T_65=d_interrupts[0] ? 4'h0:_which_T_64; 
  assign _which_T_66=d_interrupts[8] ? 4'h8:_which_T_65; 
  assign _which_T_67=d_interrupts[5] ? 4'h5:_which_T_66; 
  assign _which_T_68=d_interrupts[1] ? 4'h1:_which_T_67; 
  assign _which_T_69=d_interrupts[9] ? 4'h9:_which_T_68; 
  assign _which_T_70=d_interrupts[7] ? 4'h7:_which_T_69; 
  assign _which_T_71=d_interrupts[3] ? 4'h3:_which_T_70; 
  assign _which_T_72=d_interrupts[11] ? 4'hb:_which_T_71; 
  assign _which_T_73=d_interrupts[12] ? 4'hc:_which_T_72; 
  assign _which_T_74=d_interrupts[13] ? 4'hd:_which_T_73; 
  assign whichInterrupt=d_interrupts[14] ? 4'he:_which_T_74; 
  assign _GEN_556={60'b0,whichInterrupt}; 
  assign _io_interrupt_T_1=anyInterrupt&~io_singleStep; 
  assign _io_interrupt_T_2=_io_interrupt_T_1|reg_singleStepped; 
  assign _io_interrupt_T_3=reg_debug|io_status_cease; 
  assign pmp_mask_base_lo=reg_pmp_0_cfg_a[0]; 
  assign pmp_mask_base={reg_pmp_0_addr,pmp_mask_base_lo}; 
  assign _pmp_mask_T_1=pmp_mask_base+31'h1; 
  assign pmp_mask_hi=pmp_mask_base&~_pmp_mask_T_1; 
  assign _pmp_mask_T_3={pmp_mask_hi,2'h3}; 
  assign pmp_mask_base_lo_1=reg_pmp_1_cfg_a[0]; 
  assign pmp_mask_base_1={reg_pmp_1_addr,pmp_mask_base_lo_1}; 
  assign _pmp_mask_T_5=pmp_mask_base_1+31'h1; 
  assign pmp_mask_hi_1=pmp_mask_base_1&~_pmp_mask_T_5; 
  assign _pmp_mask_T_7={pmp_mask_hi_1,2'h3}; 
  assign pmp_mask_base_lo_2=reg_pmp_2_cfg_a[0]; 
  assign pmp_mask_base_2={reg_pmp_2_addr,pmp_mask_base_lo_2}; 
  assign _pmp_mask_T_9=pmp_mask_base_2+31'h1; 
  assign pmp_mask_hi_2=pmp_mask_base_2&~_pmp_mask_T_9; 
  assign _pmp_mask_T_11={pmp_mask_hi_2,2'h3}; 
  assign pmp_mask_base_lo_3=reg_pmp_3_cfg_a[0]; 
  assign pmp_mask_base_3={reg_pmp_3_addr,pmp_mask_base_lo_3}; 
  assign _pmp_mask_T_13=pmp_mask_base_3+31'h1; 
  assign pmp_mask_hi_3=pmp_mask_base_3&~_pmp_mask_T_13; 
  assign _pmp_mask_T_15={pmp_mask_hi_3,2'h3}; 
  assign pmp_mask_base_lo_4=reg_pmp_4_cfg_a[0]; 
  assign pmp_mask_base_4={reg_pmp_4_addr,pmp_mask_base_lo_4}; 
  assign _pmp_mask_T_17=pmp_mask_base_4+31'h1; 
  assign pmp_mask_hi_4=pmp_mask_base_4&~_pmp_mask_T_17; 
  assign _pmp_mask_T_19={pmp_mask_hi_4,2'h3}; 
  assign pmp_mask_base_lo_5=reg_pmp_5_cfg_a[0]; 
  assign pmp_mask_base_5={reg_pmp_5_addr,pmp_mask_base_lo_5}; 
  assign _pmp_mask_T_21=pmp_mask_base_5+31'h1; 
  assign pmp_mask_hi_5=pmp_mask_base_5&~_pmp_mask_T_21; 
  assign _pmp_mask_T_23={pmp_mask_hi_5,2'h3}; 
  assign pmp_mask_base_lo_6=reg_pmp_6_cfg_a[0]; 
  assign pmp_mask_base_6={reg_pmp_6_addr,pmp_mask_base_lo_6}; 
  assign _pmp_mask_T_25=pmp_mask_base_6+31'h1; 
  assign pmp_mask_hi_6=pmp_mask_base_6&~_pmp_mask_T_25; 
  assign _pmp_mask_T_27={pmp_mask_hi_6,2'h3}; 
  assign pmp_mask_base_lo_7=reg_pmp_7_cfg_a[0]; 
  assign pmp_mask_base_7={reg_pmp_7_addr,pmp_mask_base_lo_7}; 
  assign _pmp_mask_T_29=pmp_mask_base_7+31'h1; 
  assign pmp_mask_hi_7=pmp_mask_base_7&~_pmp_mask_T_29; 
  assign _pmp_mask_T_31={pmp_mask_hi_7,2'h3}; 
  assign read_mstatus_lo_lo={io_status_hpie,io_status_spie,io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie}; 
  assign read_mstatus_lo={io_status_sum,io_status_mprv,io_status_xs,io_status_fs,io_status_mpp,io_status_vs,io_status_spp,io_status_mpie,read_mstatus_lo_lo}; 
  assign read_mstatus_hi_lo={io_status_sxl,io_status_uxl,io_status_sd_rv32,io_status_zero1,io_status_tsr,io_status_tw,io_status_tvm,io_status_mxr}; 
  assign _read_mstatus_T={io_status_debug,io_status_cease,io_status_wfi,io_status_isa,io_status_dprv,io_status_prv,io_status_sd,io_status_zero2,read_mstatus_hi_lo,read_mstatus_lo}; 
   reg [63:0] reg_mstatus ;  
  assign reg_mstatus=read_mstatus; 
  assign read_mstatus=_read_mstatus_T[63:0]; 
  assign _read_mtvec_T_1=reg_mtvec[0] ? 8'hfe:8'h2; 
  assign _read_mtvec_T_3={24'b0,_read_mtvec_T_1}; 
  assign read_mtvec_lo=reg_mtvec&~_read_mtvec_T_3; 
  assign read_mtvec={32'h0,read_mtvec_lo}; 
  assign _read_stvec_T_1=reg_stvec[0] ? 8'hfe:8'h2; 
  assign _read_stvec_T_3={31'b0,_read_stvec_T_1}; 
  assign read_stvec_lo=reg_stvec&~_read_stvec_T_3; 
  assign read_stvec_hi=read_stvec_lo[38] ? 25'h1ffffff:25'h0; 
  assign read_stvec={read_stvec_hi,read_stvec_lo}; 
  assign lo_2={reg_bp_0_control_m,1'h0,reg_bp_0_control_s,reg_bp_0_control_u,reg_bp_0_control_x,reg_bp_0_control_w,reg_bp_0_control_r}; 
  assign _T_7={4'h2,reg_bp_0_control_dmode,46'h40000000000,reg_bp_0_control_action,1'h0,2'h0,reg_bp_0_control_tmatch,lo_2}; 
  assign hi_3=reg_bp_0_address[38] ? 25'h1ffffff:25'h0; 
  assign _T_10={hi_3,reg_bp_0_address}; 
  assign _T_14=reg_misa[2] ? 2'h1:2'h3; 
  assign _GEN_557={38'b0,_T_14}; 
  assign _T_15=~reg_mepc|_GEN_557; 
  assign lo_4=~_T_15; 
  assign hi_5=lo_4[39] ? 24'hffffff:24'h0; 
  assign _T_18={hi_5,lo_4}; 
  assign hi_6=reg_mtval[39] ? 24'hffffff:24'h0; 
  assign _T_21={hi_6,reg_mtval}; 
  assign lo_5={2'h0,1'h0,reg_dcsr_cause,3'h0,reg_dcsr_step,reg_dcsr_prv}; 
  assign _T_22={4'h4,12'h0,reg_dcsr_ebreakm,1'h0,reg_dcsr_ebreaks,reg_dcsr_ebreaku,lo_5}; 
   reg [31:0] reg_dcsr ;  
  assign reg_dcsr=_T_22; 
  assign _T_26=~reg_dpc|_GEN_557; 
  assign lo_6=~_T_26; 
  assign hi_8=lo_6[39] ? 24'hffffff:24'h0; 
  assign _T_29={hi_8,lo_6}; 
   reg [7:0] reg_fcsr ;  
  assign reg_fcsr=read_fcsr; 
  assign read_fcsr={reg_frm,reg_fflags}; 
  assign read_sie=reg_mie&read_mideleg; 
  assign read_sip=_GEN_45&read_mideleg; 
  assign lo_lo_4={1'h0,io_status_spie,2'h0,1'h0,io_status_sie,1'h0}; 
  assign lo_7={io_status_sum,1'h0,io_status_xs,io_status_fs,2'h0,io_status_vs,io_status_spp,1'h0,lo_lo_4}; 
  assign hi_lo_4={2'h0,io_status_uxl,io_status_sd_rv32,8'h0,2'h0,1'h0,io_status_mxr}; 
  assign _T_30={35'h0,4'h0,io_status_sd,27'h0,hi_lo_4,lo_7}; 
  assign hi_10=reg_stval[39] ? 24'hffffff:24'h0; 
  assign _T_34={hi_10,reg_stval}; 
   reg [63:0] reg_satp ;  
  assign reg_satp=_T_35; 
  assign _T_35={reg_satp_mode,16'h0,reg_satp_ppn}; 
  assign _T_39=~reg_sepc|_GEN_557; 
  assign lo_8=~_T_39; 
  assign hi_12=lo_8[39] ? 24'hffffff:24'h0; 
  assign _T_42={hi_12,lo_8}; 
  assign lo_lo_lo_3={reg_pmp_0_cfg_l,2'h0,reg_pmp_0_cfg_a,reg_pmp_0_cfg_x,reg_pmp_0_cfg_w,reg_pmp_0_cfg_r}; 
  assign lo_hi_lo_5={reg_pmp_2_cfg_l,2'h0,reg_pmp_2_cfg_a,reg_pmp_2_cfg_x,reg_pmp_2_cfg_w,reg_pmp_2_cfg_r}; 
  assign hi_lo_lo_4={reg_pmp_4_cfg_l,2'h0,reg_pmp_4_cfg_a,reg_pmp_4_cfg_x,reg_pmp_4_cfg_w,reg_pmp_4_cfg_r}; 
  assign hi_hi_lo_5={reg_pmp_6_cfg_l,2'h0,reg_pmp_6_cfg_a,reg_pmp_6_cfg_x,reg_pmp_6_cfg_w,reg_pmp_6_cfg_r}; 
  assign lo_lo_5={reg_pmp_1_cfg_l,2'h0,reg_pmp_1_cfg_a,reg_pmp_1_cfg_x,reg_pmp_1_cfg_w,reg_pmp_1_cfg_r,lo_lo_lo_3}; 
  assign lo_17={reg_pmp_3_cfg_l,2'h0,reg_pmp_3_cfg_a,reg_pmp_3_cfg_x,reg_pmp_3_cfg_w,reg_pmp_3_cfg_r,lo_hi_lo_5,lo_lo_5}; 
  assign hi_lo_5={reg_pmp_5_cfg_l,2'h0,reg_pmp_5_cfg_a,reg_pmp_5_cfg_x,reg_pmp_5_cfg_w,reg_pmp_5_cfg_r,hi_lo_lo_4}; 
  assign _T_43={reg_pmp_7_cfg_l,2'h0,reg_pmp_7_cfg_a,reg_pmp_7_cfg_x,reg_pmp_7_cfg_w,reg_pmp_7_cfg_r,hi_hi_lo_5,hi_lo_5,lo_17}; 
   reg [63:0] pmpcfg0 ;  
  assign pmpcfg0=_T_43; 
  assign _T_46=io_rw_addr==12'h7a1; 
  assign _T_47=io_rw_addr==12'h7a2; 
  assign _T_49=io_rw_addr==12'h301; 
  assign _T_50=io_rw_addr==12'h300; 
  assign _T_51=io_rw_addr==12'h305; 
  assign _T_52=io_rw_addr==12'h344; 
  assign _T_53=io_rw_addr==12'h304; 
  assign _T_54=io_rw_addr==12'h340; 
  assign _T_55=io_rw_addr==12'h341; 
  assign _T_56=io_rw_addr==12'h343; 
  assign _T_57=io_rw_addr==12'h342; 
  assign _T_58=io_rw_addr==12'hf14; 
  assign _T_59=io_rw_addr==12'h7b0; 
  assign _T_60=io_rw_addr==12'h7b1; 
  assign _T_61=io_rw_addr==12'h7b2; 
  assign _T_62=io_rw_addr==12'h1; 
  assign _T_63=io_rw_addr==12'h2; 
  assign _T_64=io_rw_addr==12'h3; 
  assign _T_65=io_rw_addr==12'h320; 
  assign _T_66=io_rw_addr==12'hb00; 
  assign _T_67=io_rw_addr==12'hb02; 
  assign _T_155=io_rw_addr==12'h306; 
  assign _T_156=io_rw_addr==12'hc00; 
  assign _T_157=io_rw_addr==12'hc02; 
  assign _T_158=io_rw_addr==12'h100; 
  assign _T_159=io_rw_addr==12'h144; 
  assign _T_160=io_rw_addr==12'h104; 
  assign _T_161=io_rw_addr==12'h140; 
  assign _T_162=io_rw_addr==12'h142; 
  assign _T_163=io_rw_addr==12'h143; 
  assign _T_164=io_rw_addr==12'h180; 
  assign _T_165=io_rw_addr==12'h141; 
  assign _T_166=io_rw_addr==12'h105; 
  assign _T_167=io_rw_addr==12'h106; 
  assign _T_168=io_rw_addr==12'h303; 
  assign _T_169=io_rw_addr==12'h302; 
  assign _T_170=io_rw_addr==12'h3a0; 
  assign _T_172=io_rw_addr==12'h3b0; 
  assign _T_173=io_rw_addr==12'h3b1; 
  assign _T_174=io_rw_addr==12'h3b2; 
  assign _T_175=io_rw_addr==12'h3b3; 
  assign _T_176=io_rw_addr==12'h3b4; 
  assign _T_177=io_rw_addr==12'h3b5; 
  assign _T_178=io_rw_addr==12'h3b6; 
  assign _T_179=io_rw_addr==12'h3b7; 
  assign _T_188=io_rw_addr==12'h7c1; 
  assign _T_189=io_rw_addr==12'hf12; 
  assign _T_191=io_rw_addr==12'hf13; 
  assign _wdata_T_1=io_rw_cmd[1] ? io_rw_rdata:64'h0; 
  assign _wdata_T_2=_wdata_T_1|io_rw_wdata; 
  assign _wdata_T_4=&io_rw_cmd[1:0]; 
  assign _wdata_T_5=_wdata_T_4 ? io_rw_wdata:64'h0; 
  assign wdata=_wdata_T_2&~_wdata_T_5; 
  assign _T_205=_T_192&32'h20200000; 
  assign _T_206=_T_205==32'h20000000; 
  assign _T_208=_T_192&32'h32200000; 
  assign _T_209=_T_208==32'h10000000; 
  assign insn_cease=system_insn&_T_206; 
  assign insn_wfi=system_insn&_T_209; 
  assign _T_220={io_decode_0_csr,20'h0}; 
  assign _T_227=_T_220&32'h12400000; 
  assign _T_228=_T_227==32'h10000000; 
  assign _T_229=_T_220&32'h40000000; 
  assign _T_230=_T_229==32'h40000000; 
  assign is_ret=_T_228|_T_230; 
  assign _T_236=_T_220&32'h32200000; 
  assign is_wfi=_T_236==32'h10000000; 
  assign _T_239=_T_220&32'h42000000; 
  assign is_sfence=_T_239==32'h2000000; 
  assign _allow_wfi_T=reg_mstatus_prv>2'h1; 
  assign allow_wfi=_allow_wfi_T|~reg_mstatus_tw; 
  assign allow_sfence_vma=_allow_wfi_T|~reg_mstatus_tvm; 
  assign allow_sret=_allow_wfi_T|~reg_mstatus_tsr; 
  assign counter_addr=io_decode_0_csr[4:0]; 
  assign _allow_counter_T_1=read_mcounteren>>counter_addr; 
  assign _allow_counter_T_3=_allow_wfi_T|_allow_counter_T_1[0]; 
  assign _allow_counter_T_4=reg_mstatus_prv>=2'h1; 
  assign _allow_counter_T_6=read_scounteren>>counter_addr; 
  assign _allow_counter_T_8=_allow_counter_T_4|_allow_counter_T_6[0]; 
  assign allow_counter=_allow_counter_T_3&_allow_counter_T_8; 
  assign _io_decode_0_fp_illegal_T=io_status_fs==2'h0; 
  assign _io_decode_0_fp_csr_T=io_decode_0_csr&12'h900; 
  assign _io_decode_0_read_illegal_T_1=reg_mstatus_prv<io_decode_0_csr[9:8]; 
  assign _io_decode_0_read_illegal_T_2=io_decode_0_csr==12'h7a0; 
  assign _io_decode_0_read_illegal_T_3=io_decode_0_csr==12'h7a1; 
  assign _io_decode_0_read_illegal_T_4=io_decode_0_csr==12'h7a2; 
  assign _io_decode_0_read_illegal_T_5=io_decode_0_csr==12'h7a3; 
  assign _io_decode_0_read_illegal_T_6=io_decode_0_csr==12'h301; 
  assign _io_decode_0_read_illegal_T_7=io_decode_0_csr==12'h300; 
  assign _io_decode_0_read_illegal_T_8=io_decode_0_csr==12'h305; 
  assign _io_decode_0_read_illegal_T_9=io_decode_0_csr==12'h344; 
  assign _io_decode_0_read_illegal_T_10=io_decode_0_csr==12'h304; 
  assign _io_decode_0_read_illegal_T_11=io_decode_0_csr==12'h340; 
  assign _io_decode_0_read_illegal_T_12=io_decode_0_csr==12'h341; 
  assign _io_decode_0_read_illegal_T_13=io_decode_0_csr==12'h343; 
  assign _io_decode_0_read_illegal_T_14=io_decode_0_csr==12'h342; 
  assign _io_decode_0_read_illegal_T_15=io_decode_0_csr==12'hf14; 
  assign _io_decode_0_read_illegal_T_16=io_decode_0_csr==12'h7b0; 
  assign _io_decode_0_read_illegal_T_17=io_decode_0_csr==12'h7b1; 
  assign _io_decode_0_read_illegal_T_18=io_decode_0_csr==12'h7b2; 
  assign _io_decode_0_read_illegal_T_19=io_decode_0_csr==12'h1; 
  assign _io_decode_0_read_illegal_T_20=io_decode_0_csr==12'h2; 
  assign _io_decode_0_read_illegal_T_21=io_decode_0_csr==12'h3; 
  assign _io_decode_0_read_illegal_T_22=io_decode_0_csr==12'h320; 
  assign _io_decode_0_read_illegal_T_23=io_decode_0_csr==12'hb00; 
  assign _io_decode_0_read_illegal_T_24=io_decode_0_csr==12'hb02; 
  assign _io_decode_0_read_illegal_T_25=io_decode_0_csr==12'h323; 
  assign _io_decode_0_read_illegal_T_26=io_decode_0_csr==12'hb03; 
  assign _io_decode_0_read_illegal_T_27=io_decode_0_csr==12'hc03; 
  assign _io_decode_0_read_illegal_T_28=io_decode_0_csr==12'h324; 
  assign _io_decode_0_read_illegal_T_29=io_decode_0_csr==12'hb04; 
  assign _io_decode_0_read_illegal_T_30=io_decode_0_csr==12'hc04; 
  assign _io_decode_0_read_illegal_T_31=io_decode_0_csr==12'h325; 
  assign _io_decode_0_read_illegal_T_32=io_decode_0_csr==12'hb05; 
  assign _io_decode_0_read_illegal_T_33=io_decode_0_csr==12'hc05; 
  assign _io_decode_0_read_illegal_T_34=io_decode_0_csr==12'h326; 
  assign _io_decode_0_read_illegal_T_35=io_decode_0_csr==12'hb06; 
  assign _io_decode_0_read_illegal_T_36=io_decode_0_csr==12'hc06; 
  assign _io_decode_0_read_illegal_T_37=io_decode_0_csr==12'h327; 
  assign _io_decode_0_read_illegal_T_38=io_decode_0_csr==12'hb07; 
  assign _io_decode_0_read_illegal_T_39=io_decode_0_csr==12'hc07; 
  assign _io_decode_0_read_illegal_T_40=io_decode_0_csr==12'h328; 
  assign _io_decode_0_read_illegal_T_41=io_decode_0_csr==12'hb08; 
  assign _io_decode_0_read_illegal_T_42=io_decode_0_csr==12'hc08; 
  assign _io_decode_0_read_illegal_T_43=io_decode_0_csr==12'h329; 
  assign _io_decode_0_read_illegal_T_44=io_decode_0_csr==12'hb09; 
  assign _io_decode_0_read_illegal_T_45=io_decode_0_csr==12'hc09; 
  assign _io_decode_0_read_illegal_T_46=io_decode_0_csr==12'h32a; 
  assign _io_decode_0_read_illegal_T_47=io_decode_0_csr==12'hb0a; 
  assign _io_decode_0_read_illegal_T_48=io_decode_0_csr==12'hc0a; 
  assign _io_decode_0_read_illegal_T_49=io_decode_0_csr==12'h32b; 
  assign _io_decode_0_read_illegal_T_50=io_decode_0_csr==12'hb0b; 
  assign _io_decode_0_read_illegal_T_51=io_decode_0_csr==12'hc0b; 
  assign _io_decode_0_read_illegal_T_52=io_decode_0_csr==12'h32c; 
  assign _io_decode_0_read_illegal_T_53=io_decode_0_csr==12'hb0c; 
  assign _io_decode_0_read_illegal_T_54=io_decode_0_csr==12'hc0c; 
  assign _io_decode_0_read_illegal_T_55=io_decode_0_csr==12'h32d; 
  assign _io_decode_0_read_illegal_T_56=io_decode_0_csr==12'hb0d; 
  assign _io_decode_0_read_illegal_T_57=io_decode_0_csr==12'hc0d; 
  assign _io_decode_0_read_illegal_T_58=io_decode_0_csr==12'h32e; 
  assign _io_decode_0_read_illegal_T_59=io_decode_0_csr==12'hb0e; 
  assign _io_decode_0_read_illegal_T_60=io_decode_0_csr==12'hc0e; 
  assign _io_decode_0_read_illegal_T_61=io_decode_0_csr==12'h32f; 
  assign _io_decode_0_read_illegal_T_62=io_decode_0_csr==12'hb0f; 
  assign _io_decode_0_read_illegal_T_63=io_decode_0_csr==12'hc0f; 
  assign _io_decode_0_read_illegal_T_64=io_decode_0_csr==12'h330; 
  assign _io_decode_0_read_illegal_T_65=io_decode_0_csr==12'hb10; 
  assign _io_decode_0_read_illegal_T_66=io_decode_0_csr==12'hc10; 
  assign _io_decode_0_read_illegal_T_67=io_decode_0_csr==12'h331; 
  assign _io_decode_0_read_illegal_T_68=io_decode_0_csr==12'hb11; 
  assign _io_decode_0_read_illegal_T_69=io_decode_0_csr==12'hc11; 
  assign _io_decode_0_read_illegal_T_70=io_decode_0_csr==12'h332; 
  assign _io_decode_0_read_illegal_T_71=io_decode_0_csr==12'hb12; 
  assign _io_decode_0_read_illegal_T_72=io_decode_0_csr==12'hc12; 
  assign _io_decode_0_read_illegal_T_73=io_decode_0_csr==12'h333; 
  assign _io_decode_0_read_illegal_T_74=io_decode_0_csr==12'hb13; 
  assign _io_decode_0_read_illegal_T_75=io_decode_0_csr==12'hc13; 
  assign _io_decode_0_read_illegal_T_76=io_decode_0_csr==12'h334; 
  assign _io_decode_0_read_illegal_T_77=io_decode_0_csr==12'hb14; 
  assign _io_decode_0_read_illegal_T_78=io_decode_0_csr==12'hc14; 
  assign _io_decode_0_read_illegal_T_79=io_decode_0_csr==12'h335; 
  assign _io_decode_0_read_illegal_T_80=io_decode_0_csr==12'hb15; 
  assign _io_decode_0_read_illegal_T_81=io_decode_0_csr==12'hc15; 
  assign _io_decode_0_read_illegal_T_82=io_decode_0_csr==12'h336; 
  assign _io_decode_0_read_illegal_T_83=io_decode_0_csr==12'hb16; 
  assign _io_decode_0_read_illegal_T_84=io_decode_0_csr==12'hc16; 
  assign _io_decode_0_read_illegal_T_85=io_decode_0_csr==12'h337; 
  assign _io_decode_0_read_illegal_T_86=io_decode_0_csr==12'hb17; 
  assign _io_decode_0_read_illegal_T_87=io_decode_0_csr==12'hc17; 
  assign _io_decode_0_read_illegal_T_88=io_decode_0_csr==12'h338; 
  assign _io_decode_0_read_illegal_T_89=io_decode_0_csr==12'hb18; 
  assign _io_decode_0_read_illegal_T_90=io_decode_0_csr==12'hc18; 
  assign _io_decode_0_read_illegal_T_91=io_decode_0_csr==12'h339; 
  assign _io_decode_0_read_illegal_T_92=io_decode_0_csr==12'hb19; 
  assign _io_decode_0_read_illegal_T_93=io_decode_0_csr==12'hc19; 
  assign _io_decode_0_read_illegal_T_94=io_decode_0_csr==12'h33a; 
  assign _io_decode_0_read_illegal_T_95=io_decode_0_csr==12'hb1a; 
  assign _io_decode_0_read_illegal_T_96=io_decode_0_csr==12'hc1a; 
  assign _io_decode_0_read_illegal_T_97=io_decode_0_csr==12'h33b; 
  assign _io_decode_0_read_illegal_T_98=io_decode_0_csr==12'hb1b; 
  assign _io_decode_0_read_illegal_T_99=io_decode_0_csr==12'hc1b; 
  assign _io_decode_0_read_illegal_T_100=io_decode_0_csr==12'h33c; 
  assign _io_decode_0_read_illegal_T_101=io_decode_0_csr==12'hb1c; 
  assign _io_decode_0_read_illegal_T_102=io_decode_0_csr==12'hc1c; 
  assign _io_decode_0_read_illegal_T_103=io_decode_0_csr==12'h33d; 
  assign _io_decode_0_read_illegal_T_104=io_decode_0_csr==12'hb1d; 
  assign _io_decode_0_read_illegal_T_105=io_decode_0_csr==12'hc1d; 
  assign _io_decode_0_read_illegal_T_106=io_decode_0_csr==12'h33e; 
  assign _io_decode_0_read_illegal_T_107=io_decode_0_csr==12'hb1e; 
  assign _io_decode_0_read_illegal_T_108=io_decode_0_csr==12'hc1e; 
  assign _io_decode_0_read_illegal_T_109=io_decode_0_csr==12'h33f; 
  assign _io_decode_0_read_illegal_T_110=io_decode_0_csr==12'hb1f; 
  assign _io_decode_0_read_illegal_T_111=io_decode_0_csr==12'hc1f; 
  assign _io_decode_0_read_illegal_T_112=io_decode_0_csr==12'h306; 
  assign _io_decode_0_read_illegal_T_113=io_decode_0_csr==12'hc00; 
  assign _io_decode_0_read_illegal_T_114=io_decode_0_csr==12'hc02; 
  assign _io_decode_0_read_illegal_T_115=io_decode_0_csr==12'h100; 
  assign _io_decode_0_read_illegal_T_116=io_decode_0_csr==12'h144; 
  assign _io_decode_0_read_illegal_T_117=io_decode_0_csr==12'h104; 
  assign _io_decode_0_read_illegal_T_118=io_decode_0_csr==12'h140; 
  assign _io_decode_0_read_illegal_T_119=io_decode_0_csr==12'h142; 
  assign _io_decode_0_read_illegal_T_120=io_decode_0_csr==12'h143; 
  assign _io_decode_0_read_illegal_T_121=io_decode_0_csr==12'h180; 
  assign _io_decode_0_read_illegal_T_122=io_decode_0_csr==12'h141; 
  assign _io_decode_0_read_illegal_T_123=io_decode_0_csr==12'h105; 
  assign _io_decode_0_read_illegal_T_124=io_decode_0_csr==12'h106; 
  assign _io_decode_0_read_illegal_T_125=io_decode_0_csr==12'h303; 
  assign _io_decode_0_read_illegal_T_126=io_decode_0_csr==12'h302; 
  assign _io_decode_0_read_illegal_T_127=io_decode_0_csr==12'h3a0; 
  assign _io_decode_0_read_illegal_T_128=io_decode_0_csr==12'h3a2; 
  assign _io_decode_0_read_illegal_T_129=io_decode_0_csr==12'h3b0; 
  assign _io_decode_0_read_illegal_T_130=io_decode_0_csr==12'h3b1; 
  assign _io_decode_0_read_illegal_T_131=io_decode_0_csr==12'h3b2; 
  assign _io_decode_0_read_illegal_T_132=io_decode_0_csr==12'h3b3; 
  assign _io_decode_0_read_illegal_T_133=io_decode_0_csr==12'h3b4; 
  assign _io_decode_0_read_illegal_T_134=io_decode_0_csr==12'h3b5; 
  assign _io_decode_0_read_illegal_T_135=io_decode_0_csr==12'h3b6; 
  assign _io_decode_0_read_illegal_T_136=io_decode_0_csr==12'h3b7; 
  assign _io_decode_0_read_illegal_T_137=io_decode_0_csr==12'h3b8; 
  assign _io_decode_0_read_illegal_T_138=io_decode_0_csr==12'h3b9; 
  assign _io_decode_0_read_illegal_T_139=io_decode_0_csr==12'h3ba; 
  assign _io_decode_0_read_illegal_T_140=io_decode_0_csr==12'h3bb; 
  assign _io_decode_0_read_illegal_T_141=io_decode_0_csr==12'h3bc; 
  assign _io_decode_0_read_illegal_T_142=io_decode_0_csr==12'h3bd; 
  assign _io_decode_0_read_illegal_T_143=io_decode_0_csr==12'h3be; 
  assign _io_decode_0_read_illegal_T_144=io_decode_0_csr==12'h3bf; 
  assign _io_decode_0_read_illegal_T_145=io_decode_0_csr==12'h7c1; 
  assign _io_decode_0_read_illegal_T_146=io_decode_0_csr==12'hf12; 
  assign _io_decode_0_read_illegal_T_147=io_decode_0_csr==12'hf11; 
  assign _io_decode_0_read_illegal_T_148=io_decode_0_csr==12'hf13; 
  assign _io_decode_0_read_illegal_T_149=_io_decode_0_read_illegal_T_2|_io_decode_0_read_illegal_T_3; 
  assign _io_decode_0_read_illegal_T_150=_io_decode_0_read_illegal_T_149|_io_decode_0_read_illegal_T_4; 
  assign _io_decode_0_read_illegal_T_151=_io_decode_0_read_illegal_T_150|_io_decode_0_read_illegal_T_5; 
  assign _io_decode_0_read_illegal_T_152=_io_decode_0_read_illegal_T_151|_io_decode_0_read_illegal_T_6; 
  assign _io_decode_0_read_illegal_T_153=_io_decode_0_read_illegal_T_152|_io_decode_0_read_illegal_T_7; 
  assign _io_decode_0_read_illegal_T_154=_io_decode_0_read_illegal_T_153|_io_decode_0_read_illegal_T_8; 
  assign _io_decode_0_read_illegal_T_155=_io_decode_0_read_illegal_T_154|_io_decode_0_read_illegal_T_9; 
  assign _io_decode_0_read_illegal_T_156=_io_decode_0_read_illegal_T_155|_io_decode_0_read_illegal_T_10; 
  assign _io_decode_0_read_illegal_T_157=_io_decode_0_read_illegal_T_156|_io_decode_0_read_illegal_T_11; 
  assign _io_decode_0_read_illegal_T_158=_io_decode_0_read_illegal_T_157|_io_decode_0_read_illegal_T_12; 
  assign _io_decode_0_read_illegal_T_159=_io_decode_0_read_illegal_T_158|_io_decode_0_read_illegal_T_13; 
  assign _io_decode_0_read_illegal_T_160=_io_decode_0_read_illegal_T_159|_io_decode_0_read_illegal_T_14; 
  assign _io_decode_0_read_illegal_T_161=_io_decode_0_read_illegal_T_160|_io_decode_0_read_illegal_T_15; 
  assign _io_decode_0_read_illegal_T_162=_io_decode_0_read_illegal_T_161|_io_decode_0_read_illegal_T_16; 
  assign _io_decode_0_read_illegal_T_163=_io_decode_0_read_illegal_T_162|_io_decode_0_read_illegal_T_17; 
  assign _io_decode_0_read_illegal_T_164=_io_decode_0_read_illegal_T_163|_io_decode_0_read_illegal_T_18; 
  assign _io_decode_0_read_illegal_T_165=_io_decode_0_read_illegal_T_164|_io_decode_0_read_illegal_T_19; 
  assign _io_decode_0_read_illegal_T_166=_io_decode_0_read_illegal_T_165|_io_decode_0_read_illegal_T_20; 
  assign _io_decode_0_read_illegal_T_167=_io_decode_0_read_illegal_T_166|_io_decode_0_read_illegal_T_21; 
  assign _io_decode_0_read_illegal_T_168=_io_decode_0_read_illegal_T_167|_io_decode_0_read_illegal_T_22; 
  assign _io_decode_0_read_illegal_T_169=_io_decode_0_read_illegal_T_168|_io_decode_0_read_illegal_T_23; 
  assign _io_decode_0_read_illegal_T_170=_io_decode_0_read_illegal_T_169|_io_decode_0_read_illegal_T_24; 
  assign _io_decode_0_read_illegal_T_171=_io_decode_0_read_illegal_T_170|_io_decode_0_read_illegal_T_25; 
  assign _io_decode_0_read_illegal_T_172=_io_decode_0_read_illegal_T_171|_io_decode_0_read_illegal_T_26; 
  assign _io_decode_0_read_illegal_T_173=_io_decode_0_read_illegal_T_172|_io_decode_0_read_illegal_T_27; 
  assign _io_decode_0_read_illegal_T_174=_io_decode_0_read_illegal_T_173|_io_decode_0_read_illegal_T_28; 
  assign _io_decode_0_read_illegal_T_175=_io_decode_0_read_illegal_T_174|_io_decode_0_read_illegal_T_29; 
  assign _io_decode_0_read_illegal_T_176=_io_decode_0_read_illegal_T_175|_io_decode_0_read_illegal_T_30; 
  assign _io_decode_0_read_illegal_T_177=_io_decode_0_read_illegal_T_176|_io_decode_0_read_illegal_T_31; 
  assign _io_decode_0_read_illegal_T_178=_io_decode_0_read_illegal_T_177|_io_decode_0_read_illegal_T_32; 
  assign _io_decode_0_read_illegal_T_179=_io_decode_0_read_illegal_T_178|_io_decode_0_read_illegal_T_33; 
  assign _io_decode_0_read_illegal_T_180=_io_decode_0_read_illegal_T_179|_io_decode_0_read_illegal_T_34; 
  assign _io_decode_0_read_illegal_T_181=_io_decode_0_read_illegal_T_180|_io_decode_0_read_illegal_T_35; 
  assign _io_decode_0_read_illegal_T_182=_io_decode_0_read_illegal_T_181|_io_decode_0_read_illegal_T_36; 
  assign _io_decode_0_read_illegal_T_183=_io_decode_0_read_illegal_T_182|_io_decode_0_read_illegal_T_37; 
  assign _io_decode_0_read_illegal_T_184=_io_decode_0_read_illegal_T_183|_io_decode_0_read_illegal_T_38; 
  assign _io_decode_0_read_illegal_T_185=_io_decode_0_read_illegal_T_184|_io_decode_0_read_illegal_T_39; 
  assign _io_decode_0_read_illegal_T_186=_io_decode_0_read_illegal_T_185|_io_decode_0_read_illegal_T_40; 
  assign _io_decode_0_read_illegal_T_187=_io_decode_0_read_illegal_T_186|_io_decode_0_read_illegal_T_41; 
  assign _io_decode_0_read_illegal_T_188=_io_decode_0_read_illegal_T_187|_io_decode_0_read_illegal_T_42; 
  assign _io_decode_0_read_illegal_T_189=_io_decode_0_read_illegal_T_188|_io_decode_0_read_illegal_T_43; 
  assign _io_decode_0_read_illegal_T_190=_io_decode_0_read_illegal_T_189|_io_decode_0_read_illegal_T_44; 
  assign _io_decode_0_read_illegal_T_191=_io_decode_0_read_illegal_T_190|_io_decode_0_read_illegal_T_45; 
  assign _io_decode_0_read_illegal_T_192=_io_decode_0_read_illegal_T_191|_io_decode_0_read_illegal_T_46; 
  assign _io_decode_0_read_illegal_T_193=_io_decode_0_read_illegal_T_192|_io_decode_0_read_illegal_T_47; 
  assign _io_decode_0_read_illegal_T_194=_io_decode_0_read_illegal_T_193|_io_decode_0_read_illegal_T_48; 
  assign _io_decode_0_read_illegal_T_195=_io_decode_0_read_illegal_T_194|_io_decode_0_read_illegal_T_49; 
  assign _io_decode_0_read_illegal_T_196=_io_decode_0_read_illegal_T_195|_io_decode_0_read_illegal_T_50; 
  assign _io_decode_0_read_illegal_T_197=_io_decode_0_read_illegal_T_196|_io_decode_0_read_illegal_T_51; 
  assign _io_decode_0_read_illegal_T_198=_io_decode_0_read_illegal_T_197|_io_decode_0_read_illegal_T_52; 
  assign _io_decode_0_read_illegal_T_199=_io_decode_0_read_illegal_T_198|_io_decode_0_read_illegal_T_53; 
  assign _io_decode_0_read_illegal_T_200=_io_decode_0_read_illegal_T_199|_io_decode_0_read_illegal_T_54; 
  assign _io_decode_0_read_illegal_T_201=_io_decode_0_read_illegal_T_200|_io_decode_0_read_illegal_T_55; 
  assign _io_decode_0_read_illegal_T_202=_io_decode_0_read_illegal_T_201|_io_decode_0_read_illegal_T_56; 
  assign _io_decode_0_read_illegal_T_203=_io_decode_0_read_illegal_T_202|_io_decode_0_read_illegal_T_57; 
  assign _io_decode_0_read_illegal_T_204=_io_decode_0_read_illegal_T_203|_io_decode_0_read_illegal_T_58; 
  assign _io_decode_0_read_illegal_T_205=_io_decode_0_read_illegal_T_204|_io_decode_0_read_illegal_T_59; 
  assign _io_decode_0_read_illegal_T_206=_io_decode_0_read_illegal_T_205|_io_decode_0_read_illegal_T_60; 
  assign _io_decode_0_read_illegal_T_207=_io_decode_0_read_illegal_T_206|_io_decode_0_read_illegal_T_61; 
  assign _io_decode_0_read_illegal_T_208=_io_decode_0_read_illegal_T_207|_io_decode_0_read_illegal_T_62; 
  assign _io_decode_0_read_illegal_T_209=_io_decode_0_read_illegal_T_208|_io_decode_0_read_illegal_T_63; 
  assign _io_decode_0_read_illegal_T_210=_io_decode_0_read_illegal_T_209|_io_decode_0_read_illegal_T_64; 
  assign _io_decode_0_read_illegal_T_211=_io_decode_0_read_illegal_T_210|_io_decode_0_read_illegal_T_65; 
  assign _io_decode_0_read_illegal_T_212=_io_decode_0_read_illegal_T_211|_io_decode_0_read_illegal_T_66; 
  assign _io_decode_0_read_illegal_T_213=_io_decode_0_read_illegal_T_212|_io_decode_0_read_illegal_T_67; 
  assign _io_decode_0_read_illegal_T_214=_io_decode_0_read_illegal_T_213|_io_decode_0_read_illegal_T_68; 
  assign _io_decode_0_read_illegal_T_215=_io_decode_0_read_illegal_T_214|_io_decode_0_read_illegal_T_69; 
  assign _io_decode_0_read_illegal_T_216=_io_decode_0_read_illegal_T_215|_io_decode_0_read_illegal_T_70; 
  assign _io_decode_0_read_illegal_T_217=_io_decode_0_read_illegal_T_216|_io_decode_0_read_illegal_T_71; 
  assign _io_decode_0_read_illegal_T_218=_io_decode_0_read_illegal_T_217|_io_decode_0_read_illegal_T_72; 
  assign _io_decode_0_read_illegal_T_219=_io_decode_0_read_illegal_T_218|_io_decode_0_read_illegal_T_73; 
  assign _io_decode_0_read_illegal_T_220=_io_decode_0_read_illegal_T_219|_io_decode_0_read_illegal_T_74; 
  assign _io_decode_0_read_illegal_T_221=_io_decode_0_read_illegal_T_220|_io_decode_0_read_illegal_T_75; 
  assign _io_decode_0_read_illegal_T_222=_io_decode_0_read_illegal_T_221|_io_decode_0_read_illegal_T_76; 
  assign _io_decode_0_read_illegal_T_223=_io_decode_0_read_illegal_T_222|_io_decode_0_read_illegal_T_77; 
  assign _io_decode_0_read_illegal_T_224=_io_decode_0_read_illegal_T_223|_io_decode_0_read_illegal_T_78; 
  assign _io_decode_0_read_illegal_T_225=_io_decode_0_read_illegal_T_224|_io_decode_0_read_illegal_T_79; 
  assign _io_decode_0_read_illegal_T_226=_io_decode_0_read_illegal_T_225|_io_decode_0_read_illegal_T_80; 
  assign _io_decode_0_read_illegal_T_227=_io_decode_0_read_illegal_T_226|_io_decode_0_read_illegal_T_81; 
  assign _io_decode_0_read_illegal_T_228=_io_decode_0_read_illegal_T_227|_io_decode_0_read_illegal_T_82; 
  assign _io_decode_0_read_illegal_T_229=_io_decode_0_read_illegal_T_228|_io_decode_0_read_illegal_T_83; 
  assign _io_decode_0_read_illegal_T_230=_io_decode_0_read_illegal_T_229|_io_decode_0_read_illegal_T_84; 
  assign _io_decode_0_read_illegal_T_231=_io_decode_0_read_illegal_T_230|_io_decode_0_read_illegal_T_85; 
  assign _io_decode_0_read_illegal_T_232=_io_decode_0_read_illegal_T_231|_io_decode_0_read_illegal_T_86; 
  assign _io_decode_0_read_illegal_T_233=_io_decode_0_read_illegal_T_232|_io_decode_0_read_illegal_T_87; 
  assign _io_decode_0_read_illegal_T_234=_io_decode_0_read_illegal_T_233|_io_decode_0_read_illegal_T_88; 
  assign _io_decode_0_read_illegal_T_235=_io_decode_0_read_illegal_T_234|_io_decode_0_read_illegal_T_89; 
  assign _io_decode_0_read_illegal_T_236=_io_decode_0_read_illegal_T_235|_io_decode_0_read_illegal_T_90; 
  assign _io_decode_0_read_illegal_T_237=_io_decode_0_read_illegal_T_236|_io_decode_0_read_illegal_T_91; 
  assign _io_decode_0_read_illegal_T_238=_io_decode_0_read_illegal_T_237|_io_decode_0_read_illegal_T_92; 
  assign _io_decode_0_read_illegal_T_239=_io_decode_0_read_illegal_T_238|_io_decode_0_read_illegal_T_93; 
  assign _io_decode_0_read_illegal_T_240=_io_decode_0_read_illegal_T_239|_io_decode_0_read_illegal_T_94; 
  assign _io_decode_0_read_illegal_T_241=_io_decode_0_read_illegal_T_240|_io_decode_0_read_illegal_T_95; 
  assign _io_decode_0_read_illegal_T_242=_io_decode_0_read_illegal_T_241|_io_decode_0_read_illegal_T_96; 
  assign _io_decode_0_read_illegal_T_243=_io_decode_0_read_illegal_T_242|_io_decode_0_read_illegal_T_97; 
  assign _io_decode_0_read_illegal_T_244=_io_decode_0_read_illegal_T_243|_io_decode_0_read_illegal_T_98; 
  assign _io_decode_0_read_illegal_T_245=_io_decode_0_read_illegal_T_244|_io_decode_0_read_illegal_T_99; 
  assign _io_decode_0_read_illegal_T_246=_io_decode_0_read_illegal_T_245|_io_decode_0_read_illegal_T_100; 
  assign _io_decode_0_read_illegal_T_247=_io_decode_0_read_illegal_T_246|_io_decode_0_read_illegal_T_101; 
  assign _io_decode_0_read_illegal_T_248=_io_decode_0_read_illegal_T_247|_io_decode_0_read_illegal_T_102; 
  assign _io_decode_0_read_illegal_T_249=_io_decode_0_read_illegal_T_248|_io_decode_0_read_illegal_T_103; 
  assign _io_decode_0_read_illegal_T_250=_io_decode_0_read_illegal_T_249|_io_decode_0_read_illegal_T_104; 
  assign _io_decode_0_read_illegal_T_251=_io_decode_0_read_illegal_T_250|_io_decode_0_read_illegal_T_105; 
  assign _io_decode_0_read_illegal_T_252=_io_decode_0_read_illegal_T_251|_io_decode_0_read_illegal_T_106; 
  assign _io_decode_0_read_illegal_T_253=_io_decode_0_read_illegal_T_252|_io_decode_0_read_illegal_T_107; 
  assign _io_decode_0_read_illegal_T_254=_io_decode_0_read_illegal_T_253|_io_decode_0_read_illegal_T_108; 
  assign _io_decode_0_read_illegal_T_255=_io_decode_0_read_illegal_T_254|_io_decode_0_read_illegal_T_109; 
  assign _io_decode_0_read_illegal_T_256=_io_decode_0_read_illegal_T_255|_io_decode_0_read_illegal_T_110; 
  assign _io_decode_0_read_illegal_T_257=_io_decode_0_read_illegal_T_256|_io_decode_0_read_illegal_T_111; 
  assign _io_decode_0_read_illegal_T_258=_io_decode_0_read_illegal_T_257|_io_decode_0_read_illegal_T_112; 
  assign _io_decode_0_read_illegal_T_259=_io_decode_0_read_illegal_T_258|_io_decode_0_read_illegal_T_113; 
  assign _io_decode_0_read_illegal_T_260=_io_decode_0_read_illegal_T_259|_io_decode_0_read_illegal_T_114; 
  assign _io_decode_0_read_illegal_T_261=_io_decode_0_read_illegal_T_260|_io_decode_0_read_illegal_T_115; 
  assign _io_decode_0_read_illegal_T_262=_io_decode_0_read_illegal_T_261|_io_decode_0_read_illegal_T_116; 
  assign _io_decode_0_read_illegal_T_263=_io_decode_0_read_illegal_T_262|_io_decode_0_read_illegal_T_117; 
  assign _io_decode_0_read_illegal_T_264=_io_decode_0_read_illegal_T_263|_io_decode_0_read_illegal_T_118; 
  assign _io_decode_0_read_illegal_T_265=_io_decode_0_read_illegal_T_264|_io_decode_0_read_illegal_T_119; 
  assign _io_decode_0_read_illegal_T_266=_io_decode_0_read_illegal_T_265|_io_decode_0_read_illegal_T_120; 
  assign _io_decode_0_read_illegal_T_267=_io_decode_0_read_illegal_T_266|_io_decode_0_read_illegal_T_121; 
  assign _io_decode_0_read_illegal_T_268=_io_decode_0_read_illegal_T_267|_io_decode_0_read_illegal_T_122; 
  assign _io_decode_0_read_illegal_T_269=_io_decode_0_read_illegal_T_268|_io_decode_0_read_illegal_T_123; 
  assign _io_decode_0_read_illegal_T_270=_io_decode_0_read_illegal_T_269|_io_decode_0_read_illegal_T_124; 
  assign _io_decode_0_read_illegal_T_271=_io_decode_0_read_illegal_T_270|_io_decode_0_read_illegal_T_125; 
  assign _io_decode_0_read_illegal_T_272=_io_decode_0_read_illegal_T_271|_io_decode_0_read_illegal_T_126; 
  assign _io_decode_0_read_illegal_T_273=_io_decode_0_read_illegal_T_272|_io_decode_0_read_illegal_T_127; 
  assign _io_decode_0_read_illegal_T_274=_io_decode_0_read_illegal_T_273|_io_decode_0_read_illegal_T_128; 
  assign _io_decode_0_read_illegal_T_275=_io_decode_0_read_illegal_T_274|_io_decode_0_read_illegal_T_129; 
  assign _io_decode_0_read_illegal_T_276=_io_decode_0_read_illegal_T_275|_io_decode_0_read_illegal_T_130; 
  assign _io_decode_0_read_illegal_T_277=_io_decode_0_read_illegal_T_276|_io_decode_0_read_illegal_T_131; 
  assign _io_decode_0_read_illegal_T_278=_io_decode_0_read_illegal_T_277|_io_decode_0_read_illegal_T_132; 
  assign _io_decode_0_read_illegal_T_279=_io_decode_0_read_illegal_T_278|_io_decode_0_read_illegal_T_133; 
  assign _io_decode_0_read_illegal_T_280=_io_decode_0_read_illegal_T_279|_io_decode_0_read_illegal_T_134; 
  assign _io_decode_0_read_illegal_T_281=_io_decode_0_read_illegal_T_280|_io_decode_0_read_illegal_T_135; 
  assign _io_decode_0_read_illegal_T_282=_io_decode_0_read_illegal_T_281|_io_decode_0_read_illegal_T_136; 
  assign _io_decode_0_read_illegal_T_283=_io_decode_0_read_illegal_T_282|_io_decode_0_read_illegal_T_137; 
  assign _io_decode_0_read_illegal_T_284=_io_decode_0_read_illegal_T_283|_io_decode_0_read_illegal_T_138; 
  assign _io_decode_0_read_illegal_T_285=_io_decode_0_read_illegal_T_284|_io_decode_0_read_illegal_T_139; 
  assign _io_decode_0_read_illegal_T_286=_io_decode_0_read_illegal_T_285|_io_decode_0_read_illegal_T_140; 
  assign _io_decode_0_read_illegal_T_287=_io_decode_0_read_illegal_T_286|_io_decode_0_read_illegal_T_141; 
  assign _io_decode_0_read_illegal_T_288=_io_decode_0_read_illegal_T_287|_io_decode_0_read_illegal_T_142; 
  assign _io_decode_0_read_illegal_T_289=_io_decode_0_read_illegal_T_288|_io_decode_0_read_illegal_T_143; 
  assign _io_decode_0_read_illegal_T_290=_io_decode_0_read_illegal_T_289|_io_decode_0_read_illegal_T_144; 
  assign _io_decode_0_read_illegal_T_291=_io_decode_0_read_illegal_T_290|_io_decode_0_read_illegal_T_145; 
  assign _io_decode_0_read_illegal_T_292=_io_decode_0_read_illegal_T_291|_io_decode_0_read_illegal_T_146; 
  assign _io_decode_0_read_illegal_T_293=_io_decode_0_read_illegal_T_292|_io_decode_0_read_illegal_T_147; 
  assign _io_decode_0_read_illegal_T_294=_io_decode_0_read_illegal_T_293|_io_decode_0_read_illegal_T_148; 
  assign _io_decode_0_read_illegal_T_296=_io_decode_0_read_illegal_T_1|~_io_decode_0_read_illegal_T_294; 
  assign _io_decode_0_read_illegal_T_299=_io_decode_0_read_illegal_T_121&~allow_sfence_vma; 
  assign _io_decode_0_read_illegal_T_300=_io_decode_0_read_illegal_T_296|_io_decode_0_read_illegal_T_299; 
  assign _io_decode_0_read_illegal_T_301=io_decode_0_csr>=12'hc00; 
  assign _io_decode_0_read_illegal_T_302=io_decode_0_csr<12'hc20; 
  assign _io_decode_0_read_illegal_T_303=_io_decode_0_read_illegal_T_301&_io_decode_0_read_illegal_T_302; 
  assign _io_decode_0_read_illegal_T_304=io_decode_0_csr>=12'hc80; 
  assign _io_decode_0_read_illegal_T_305=io_decode_0_csr<12'hca0; 
  assign _io_decode_0_read_illegal_T_306=_io_decode_0_read_illegal_T_304&_io_decode_0_read_illegal_T_305; 
  assign _io_decode_0_read_illegal_T_307=_io_decode_0_read_illegal_T_303|_io_decode_0_read_illegal_T_306; 
  assign _io_decode_0_read_illegal_T_309=_io_decode_0_read_illegal_T_307&~allow_counter; 
  assign _io_decode_0_read_illegal_T_310=_io_decode_0_read_illegal_T_300|_io_decode_0_read_illegal_T_309; 
  assign _io_decode_0_read_illegal_T_311=io_decode_0_csr&12'hc10; 
  assign _io_decode_0_read_illegal_T_312=_io_decode_0_read_illegal_T_311==12'h410; 
  assign _io_decode_0_read_illegal_T_316=_io_decode_0_read_illegal_T_312&~reg_debug; 
  assign _io_decode_0_read_illegal_T_317=_io_decode_0_read_illegal_T_310|_io_decode_0_read_illegal_T_316; 
  assign _io_decode_0_read_illegal_T_320=io_decode_0_fp_csr&io_decode_0_fp_illegal; 
  assign _io_decode_0_write_flush_T=io_decode_0_csr>=12'h340; 
  assign _io_decode_0_write_flush_T_1=io_decode_0_csr<=12'h343; 
  assign _io_decode_0_write_flush_T_2=_io_decode_0_write_flush_T&_io_decode_0_write_flush_T_1; 
  assign _io_decode_0_write_flush_T_3=io_decode_0_csr>=12'h140; 
  assign _io_decode_0_write_flush_T_4=io_decode_0_csr<=12'h143; 
  assign _io_decode_0_write_flush_T_5=_io_decode_0_write_flush_T_3&_io_decode_0_write_flush_T_4; 
  assign _io_decode_0_write_flush_T_6=_io_decode_0_write_flush_T_2|_io_decode_0_write_flush_T_5; 
  assign _io_decode_0_system_illegal_T_3=is_wfi&~allow_wfi; 
  assign _io_decode_0_system_illegal_T_4=_io_decode_0_read_illegal_T_1|_io_decode_0_system_illegal_T_3; 
  assign _io_decode_0_system_illegal_T_6=is_ret&~allow_sret; 
  assign _io_decode_0_system_illegal_T_7=_io_decode_0_system_illegal_T_4|_io_decode_0_system_illegal_T_6; 
  assign _io_decode_0_system_illegal_T_9=is_ret&io_decode_0_csr[10]; 
  assign _io_decode_0_system_illegal_T_11=_io_decode_0_system_illegal_T_9&io_decode_0_csr[7]; 
  assign _io_decode_0_system_illegal_T_13=_io_decode_0_system_illegal_T_11&~reg_debug; 
  assign _io_decode_0_system_illegal_T_14=_io_decode_0_system_illegal_T_7|_io_decode_0_system_illegal_T_13; 
  assign _io_decode_0_system_illegal_T_16=is_sfence&~allow_sfence_vma; 
  assign _debugTVec_T=insn_break ? 12'h800:12'h808; 
  assign debugTVec=reg_debug ? _debugTVec_T:12'h800; 
  assign notDebugTVec_base=delegate ? read_stvec:read_mtvec; 
  assign notDebugTVec_interruptVec_lo={cause[5:0],2'h0}; 
  assign notDebugTVec_interruptVec_hi=notDebugTVec_base[63:8]; 
  assign notDebugTVec_interruptVec={notDebugTVec_interruptVec_hi,notDebugTVec_interruptVec_lo}; 
  assign _notDebugTVec_doVector_T_2=notDebugTVec_base[0]&cause[63]; 
  assign _notDebugTVec_doVector_T_4=cause_lsbs[7:6]==2'h0; 
  assign notDebugTVec_doVector=_notDebugTVec_doVector_T_2&_notDebugTVec_doVector_T_4; 
  assign _notDebugTVec_T_1={notDebugTVec_base[63:2],2'h0}; 
  assign notDebugTVec=notDebugTVec_doVector ? notDebugTVec_interruptVec:_notDebugTVec_T_1; 
  assign tvec=trapToDebug ? {52'b0,debugTVec}:notDebugTVec; 
  assign _io_status_sd_T=&io_status_fs; 
  assign _io_status_sd_T_1=&io_status_xs; 
  assign _io_status_sd_T_2=_io_status_sd_T|_io_status_sd_T_1; 
  assign _io_status_sd_T_3=&io_status_vs; 
  assign _io_status_dprv_x87_T_1=reg_mstatus_mprv&~reg_debug; 
  assign _T_244=insn_ret+insn_call; 
  assign _T_246=insn_break+io_exception; 
  assign _T_248=_T_244+_T_246; 
  assign _T_250=_T_248<=3'h1; 
  assign _T_252=_T_250|reset; 
  assign _T_255=insn_wfi&~io_singleStep; 
  assign _T_257=_T_255&~reg_debug; 
  assign _GEN_48=_T_257|reg_wfi; 
  assign _T_258=|pending_interrupts; 
  assign _T_259=_T_258|io_interrupts_debug; 
  assign _T_260=_T_259|exception; 
  assign _T_262=io_retire|exception; 
  assign _GEN_50=_T_262|reg_singleStepped; 
  assign _T_272=~reg_singleStepped|~io_retire; 
  assign _T_274=_T_272|reset; 
  assign _epc_T_1=~io_pc|40'h1; 
  assign epc=~_epc_T_1; 
  assign _reg_dcsr_cause_T=causeIsDebugTrigger ? 2'h2:2'h1; 
  assign _reg_dcsr_cause_T_1=causeIsDebugInt ? 2'h3:_reg_dcsr_cause_T; 
  assign _GEN_52=~reg_debug|reg_debug; 
  assign _GEN_53=reg_debug ? reg_dpc:epc; 
  assign _GEN_63=_T_279 ? epc:reg_sepc; 
  assign _GEN_67=_T_279 ? reg_mstatus_sie:reg_mstatus_spie; 
  assign _GEN_68=_T_279 ? reg_mstatus_prv:{1'b0,reg_mstatus_spp}; 
  assign _GEN_71=_T_279 ? reg_mepc:epc; 
  assign _GEN_74=_T_279 ? reg_mstatus_mpie:reg_mstatus_mie; 
  assign _GEN_75=_T_279 ? reg_mstatus_mpp:reg_mstatus_prv; 
  assign _GEN_76=_T_279&reg_mstatus_mie; 
  assign _GEN_97=trapToDebug ? _GEN_53:reg_dpc; 
  assign _GEN_106=trapToDebug ? reg_sepc:_GEN_63; 
  assign _GEN_110=trapToDebug ? reg_mstatus_spie:_GEN_67; 
  assign _GEN_111=trapToDebug ? {1'b0,reg_mstatus_spp}:_GEN_68; 
  assign _GEN_113=trapToDebug ? reg_mepc:_GEN_71; 
  assign _GEN_116=trapToDebug ? reg_mstatus_mpie:_GEN_74; 
  assign _GEN_117=trapToDebug ? reg_mstatus_mpp:_GEN_75; 
  assign _GEN_118=trapToDebug ? reg_mstatus_mie:_GEN_76; 
  assign _GEN_120=exception ? _GEN_97:reg_dpc; 
  assign _GEN_129=exception ? _GEN_106:reg_sepc; 
  assign _GEN_133=exception ? _GEN_110:reg_mstatus_spie; 
  assign _GEN_134=exception ? _GEN_111:{1'b0,reg_mstatus_spp}; 
  assign _GEN_136=exception ? _GEN_113:reg_mepc; 
  assign _GEN_139=exception ? _GEN_116:reg_mstatus_mpie; 
  assign _GEN_140=exception ? _GEN_117:reg_mstatus_mpp; 
  assign _GEN_141=exception ? _GEN_118:reg_mstatus_mie; 
  assign _GEN_151=_T_406 ? lo_6:lo_4; 
  assign _GEN_158=~io_rw_addr[9]|_GEN_133; 
  assign _GEN_159=io_rw_addr[9] ? _GEN_134:2'h0; 
  assign _GEN_161=io_rw_addr[9] ? _GEN_151:lo_8; 
  assign _T_412=ret_prv<2'h3; 
  assign _GEN_171=insn_ret ? _GEN_159:_GEN_134; 
  assign _GEN_172=insn_ret ? {24'b0,_GEN_161}:tvec; 
  assign _GEN_181=insn_cease|io_status_cease_r; 
  assign _io_rw_rdata_T_1=_T_46 ? _T_7:64'h0; 
  assign _io_rw_rdata_T_2=_T_47 ? _T_10:64'h0; 
  assign _io_rw_rdata_T_4=_T_49 ? reg_misa:64'h0; 
  assign _io_rw_rdata_T_5=_T_50 ? read_mstatus:64'h0; 
  assign _io_rw_rdata_T_6=_T_51 ? read_mtvec:64'h0; 
  assign _io_rw_rdata_T_7=_T_52 ? read_mip:16'h0; 
  assign _io_rw_rdata_T_8=_T_53 ? reg_mie:64'h0; 
  assign _io_rw_rdata_T_9=_T_54 ? reg_mscratch:64'h0; 
  assign _io_rw_rdata_T_10=_T_55 ? _T_18:64'h0; 
  assign _io_rw_rdata_T_11=_T_56 ? _T_21:64'h0; 
  assign _io_rw_rdata_T_12=_T_57 ? reg_mcause:64'h0; 
  assign _io_rw_rdata_T_13=_T_58&io_hartid; 
  assign _io_rw_rdata_T_14=_T_59 ? _T_22:32'h0; 
  assign _io_rw_rdata_T_15=_T_60 ? _T_29:64'h0; 
  assign _io_rw_rdata_T_16=_T_61 ? reg_dscratch:64'h0; 
  assign _io_rw_rdata_T_17=_T_62 ? reg_fflags:5'h0; 
  assign _io_rw_rdata_T_18=_T_63 ? reg_frm:3'h0; 
  assign _io_rw_rdata_T_19=_T_64 ? read_fcsr:8'h0; 
  assign _io_rw_rdata_T_20=_T_65 ? reg_mcountinhibit:3'h0; 
  assign _io_rw_rdata_T_21=_T_66 ? value_1:64'h0; 
  assign _io_rw_rdata_T_22=_T_67 ? value:64'h0; 
  assign _io_rw_rdata_T_110=_T_155 ? read_mcounteren:32'h0; 
  assign _io_rw_rdata_T_111=_T_156 ? value_1:64'h0; 
  assign _io_rw_rdata_T_112=_T_157 ? value:64'h0; 
  assign _io_rw_rdata_T_113=_T_158 ? _T_30[63:0]:64'h0; 
  assign _io_rw_rdata_T_114=_T_159 ? read_sip:64'h0; 
  assign _io_rw_rdata_T_115=_T_160 ? read_sie:64'h0; 
  assign _io_rw_rdata_T_116=_T_161 ? reg_sscratch:64'h0; 
  assign _io_rw_rdata_T_117=_T_162 ? reg_scause:64'h0; 
  assign _io_rw_rdata_T_118=_T_163 ? _T_34:64'h0; 
  assign _io_rw_rdata_T_119=_T_164 ? _T_35:64'h0; 
  assign _io_rw_rdata_T_120=_T_165 ? _T_42:64'h0; 
  assign _io_rw_rdata_T_121=_T_166 ? read_stvec:64'h0; 
  assign _io_rw_rdata_T_122=_T_167 ? read_scounteren:32'h0; 
  assign _io_rw_rdata_T_123=_T_168 ? read_mideleg:64'h0; 
  assign _io_rw_rdata_T_124=_T_169 ? read_medeleg:64'h0; 
  assign _io_rw_rdata_T_125=_T_170 ? _T_43:64'h0; 
  assign _io_rw_rdata_T_127=_T_172 ? reg_pmp_0_addr:30'h0; 
  assign _io_rw_rdata_T_128=_T_173 ? reg_pmp_1_addr:30'h0; 
  assign _io_rw_rdata_T_129=_T_174 ? reg_pmp_2_addr:30'h0; 
  assign _io_rw_rdata_T_130=_T_175 ? reg_pmp_3_addr:30'h0; 
  assign _io_rw_rdata_T_131=_T_176 ? reg_pmp_4_addr:30'h0; 
  assign _io_rw_rdata_T_132=_T_177 ? reg_pmp_5_addr:30'h0; 
  assign _io_rw_rdata_T_133=_T_178 ? reg_pmp_6_addr:30'h0; 
  assign _io_rw_rdata_T_134=_T_179 ? reg_pmp_7_addr:30'h0; 
  assign _io_rw_rdata_T_143=_T_188 ? reg_custom_0:64'h0; 
  assign _io_rw_rdata_T_144=_T_189 ? 64'h1:64'h0; 
  assign _io_rw_rdata_T_146=_T_191 ? 64'h20181004:64'h0; 
  assign _io_rw_rdata_T_148=_io_rw_rdata_T_1|_io_rw_rdata_T_2; 
  assign _io_rw_rdata_T_150=_io_rw_rdata_T_148|_io_rw_rdata_T_4; 
  assign _io_rw_rdata_T_151=_io_rw_rdata_T_150|_io_rw_rdata_T_5; 
  assign _io_rw_rdata_T_152=_io_rw_rdata_T_151|_io_rw_rdata_T_6; 
  assign _GEN_565={48'b0,_io_rw_rdata_T_7}; 
  assign _io_rw_rdata_T_153=_io_rw_rdata_T_152|_GEN_565; 
  assign _io_rw_rdata_T_154=_io_rw_rdata_T_153|_io_rw_rdata_T_8; 
  assign _io_rw_rdata_T_155=_io_rw_rdata_T_154|_io_rw_rdata_T_9; 
  assign _io_rw_rdata_T_156=_io_rw_rdata_T_155|_io_rw_rdata_T_10; 
  assign _io_rw_rdata_T_157=_io_rw_rdata_T_156|_io_rw_rdata_T_11; 
  assign _io_rw_rdata_T_158=_io_rw_rdata_T_157|_io_rw_rdata_T_12; 
  assign _GEN_566={63'b0,_io_rw_rdata_T_13}; 
  assign _io_rw_rdata_T_159=_io_rw_rdata_T_158|_GEN_566; 
  assign _GEN_567={32'b0,_io_rw_rdata_T_14}; 
  assign _io_rw_rdata_T_160=_io_rw_rdata_T_159|_GEN_567; 
  assign _io_rw_rdata_T_161=_io_rw_rdata_T_160|_io_rw_rdata_T_15; 
  assign _io_rw_rdata_T_162=_io_rw_rdata_T_161|_io_rw_rdata_T_16; 
  assign _GEN_568={59'b0,_io_rw_rdata_T_17}; 
  assign _io_rw_rdata_T_163=_io_rw_rdata_T_162|_GEN_568; 
  assign _GEN_569={61'b0,_io_rw_rdata_T_18}; 
  assign _io_rw_rdata_T_164=_io_rw_rdata_T_163|_GEN_569; 
  assign _GEN_570={56'b0,_io_rw_rdata_T_19}; 
  assign _io_rw_rdata_T_165=_io_rw_rdata_T_164|_GEN_570; 
  assign _GEN_571={61'b0,_io_rw_rdata_T_20}; 
  assign _io_rw_rdata_T_166=_io_rw_rdata_T_165|_GEN_571; 
  assign _io_rw_rdata_T_167=_io_rw_rdata_T_166|_io_rw_rdata_T_21; 
  assign _io_rw_rdata_T_168=_io_rw_rdata_T_167|_io_rw_rdata_T_22; 
  assign _GEN_572={32'b0,_io_rw_rdata_T_110}; 
  assign _io_rw_rdata_T_256=_io_rw_rdata_T_168|_GEN_572; 
  assign _io_rw_rdata_T_257=_io_rw_rdata_T_256|_io_rw_rdata_T_111; 
  assign _io_rw_rdata_T_258=_io_rw_rdata_T_257|_io_rw_rdata_T_112; 
  assign _io_rw_rdata_T_259=_io_rw_rdata_T_258|_io_rw_rdata_T_113; 
  assign _io_rw_rdata_T_260=_io_rw_rdata_T_259|_io_rw_rdata_T_114; 
  assign _io_rw_rdata_T_261=_io_rw_rdata_T_260|_io_rw_rdata_T_115; 
  assign _io_rw_rdata_T_262=_io_rw_rdata_T_261|_io_rw_rdata_T_116; 
  assign _io_rw_rdata_T_263=_io_rw_rdata_T_262|_io_rw_rdata_T_117; 
  assign _io_rw_rdata_T_264=_io_rw_rdata_T_263|_io_rw_rdata_T_118; 
  assign _io_rw_rdata_T_265=_io_rw_rdata_T_264|_io_rw_rdata_T_119; 
  assign _io_rw_rdata_T_266=_io_rw_rdata_T_265|_io_rw_rdata_T_120; 
  assign _io_rw_rdata_T_267=_io_rw_rdata_T_266|_io_rw_rdata_T_121; 
  assign _GEN_573={32'b0,_io_rw_rdata_T_122}; 
  assign _io_rw_rdata_T_268=_io_rw_rdata_T_267|_GEN_573; 
  assign _io_rw_rdata_T_269=_io_rw_rdata_T_268|_io_rw_rdata_T_123; 
  assign _io_rw_rdata_T_270=_io_rw_rdata_T_269|_io_rw_rdata_T_124; 
  assign _io_rw_rdata_T_271=_io_rw_rdata_T_270|_io_rw_rdata_T_125; 
  assign _GEN_574={34'b0,_io_rw_rdata_T_127}; 
  assign _io_rw_rdata_T_273=_io_rw_rdata_T_271|_GEN_574; 
  assign _GEN_575={34'b0,_io_rw_rdata_T_128}; 
  assign _io_rw_rdata_T_274=_io_rw_rdata_T_273|_GEN_575; 
  assign _GEN_576={34'b0,_io_rw_rdata_T_129}; 
  assign _io_rw_rdata_T_275=_io_rw_rdata_T_274|_GEN_576; 
  assign _GEN_577={34'b0,_io_rw_rdata_T_130}; 
  assign _io_rw_rdata_T_276=_io_rw_rdata_T_275|_GEN_577; 
  assign _GEN_578={34'b0,_io_rw_rdata_T_131}; 
  assign _io_rw_rdata_T_277=_io_rw_rdata_T_276|_GEN_578; 
  assign _GEN_579={34'b0,_io_rw_rdata_T_132}; 
  assign _io_rw_rdata_T_278=_io_rw_rdata_T_277|_GEN_579; 
  assign _GEN_580={34'b0,_io_rw_rdata_T_133}; 
  assign _io_rw_rdata_T_279=_io_rw_rdata_T_278|_GEN_580; 
  assign _GEN_581={34'b0,_io_rw_rdata_T_134}; 
  assign _io_rw_rdata_T_280=_io_rw_rdata_T_279|_GEN_581; 
  assign _io_rw_rdata_T_289=_io_rw_rdata_T_280|_io_rw_rdata_T_143; 
  assign _io_rw_rdata_T_290=_io_rw_rdata_T_289|_io_rw_rdata_T_144; 
  assign _T_416=io_rw_cmd==3'h5; 
  assign _T_417=io_rw_cmd==3'h6; 
  assign _T_418=io_rw_cmd==3'h7; 
  assign _lo_T=reg_fflags|io_fcsr_flags_bits; 
  assign _GEN_182=io_fcsr_flags_valid ? _lo_T:reg_fflags; 
  assign _csr_wen_T_3=_T_417|_T_418; 
  assign csr_wen=_csr_wen_T_3|_T_416; 
  assign _new_mstatus_WIRE={39'b0,wdata}; 
  assign new_mstatus_sie=_new_mstatus_WIRE[1]; 
  assign new_mstatus_mie=_new_mstatus_WIRE[3]; 
  assign new_mstatus_spie=_new_mstatus_WIRE[5]; 
  assign new_mstatus_mpie=_new_mstatus_WIRE[7]; 
  assign new_mstatus_spp=_new_mstatus_WIRE[8]; 
  assign new_mstatus_mpp=_new_mstatus_WIRE[12:11]; 
  assign new_mstatus_fs=_new_mstatus_WIRE[14:13]; 
  assign new_mstatus_mprv=_new_mstatus_WIRE[17]; 
  assign new_mstatus_sum=_new_mstatus_WIRE[18]; 
  assign new_mstatus_mxr=_new_mstatus_WIRE[19]; 
  assign new_mstatus_tvm=_new_mstatus_WIRE[20]; 
  assign new_mstatus_tw=_new_mstatus_WIRE[21]; 
  assign new_mstatus_tsr=_new_mstatus_WIRE[22]; 
  assign _reg_mstatus_mpp_T_2=new_mstatus_mpp==2'h2; 
  assign _reg_mstatus_fs_T=|new_mstatus_fs; 
  assign _GEN_188=_T_50 ? {1'b0,new_mstatus_spp}:_GEN_171; 
  assign f=wdata[5]; 
  assign _T_1834=~io_pc[1]|wdata[2]; 
  assign _reg_misa_T_2={~f,3'h0}; 
  assign _GEN_582={60'b0,_reg_misa_T_2}; 
  assign _reg_misa_T_3=~wdata|_GEN_582; 
  assign _reg_misa_T_5=~_reg_misa_T_3&64'h102d; 
  assign _reg_misa_T_7=reg_misa&64'hffffffffffffefd2; 
  assign _reg_misa_T_8=_reg_misa_T_5|_reg_misa_T_7; 
  assign _new_mip_T={4'h0,2'h0,reg_mip_seip,1'h0,2'h0,reg_mip_stip,1'h0,2'h0,reg_mip_ssip,1'h0}; 
  assign _new_mip_T_2=io_rw_cmd[1] ? _new_mip_T:16'h0; 
  assign _GEN_583={48'b0,_new_mip_T_2}; 
  assign _new_mip_T_3=_GEN_583|io_rw_wdata; 
  assign _new_mip_T_8=_new_mip_T_3&~_wdata_T_5; 
  assign new_mip_ssip=_new_mip_T_8[1]; 
  assign new_mip_stip=_new_mip_T_8[5]; 
  assign new_mip_seip=_new_mip_T_8[9]; 
  assign _reg_mie_T=wdata&64'haaa; 
  assign _reg_mepc_T_1=~wdata|64'h1; 
  assign _GEN_204=_T_55 ? ~_reg_mepc_T_1:{24'b0,_GEN_136}; 
  assign _GEN_206=_T_51 ? wdata:{32'b0,reg_mtvec}; 
  assign _reg_mcause_T=wdata&64'h800000000000000f; 
  assign _reg_mcountinhibit_T_1=wdata&64'hfffffffffffffffd; 
  assign _GEN_209=_T_65 ? _reg_mcountinhibit_T_1:{61'b0,reg_mcountinhibit}; 
  assign _GEN_210=_T_66 ? wdata:{57'b0,_GEN_2}; 
  assign _GEN_212=_T_67 ? wdata:{57'b0,_GEN_0}; 
  assign _GEN_215=_T_62 ? wdata:{59'b0,_GEN_182}; 
  assign _GEN_217=_T_63 ? wdata:{61'b0,reg_frm}; 
  assign _GEN_219=_T_64 ? wdata:_GEN_215; 
  assign _GEN_220=_T_64 ? {5'b0,wdata[63:5]}:_GEN_217; 
  assign new_dcsr_prv=wdata[1:0]; 
  assign new_dcsr_step=wdata[2]; 
  assign new_dcsr_ebreaku=wdata[12]; 
  assign new_dcsr_ebreaks=wdata[13]; 
  assign new_dcsr_ebreakm=wdata[15]; 
  assign _reg_dcsr_prv_T=new_dcsr_prv==2'h2; 
  assign _GEN_226=_T_60 ? ~_reg_mepc_T_1:{24'b0,_GEN_120}; 
  assign _GEN_230=_T_158 ? {1'b0,new_mstatus_spp}:_GEN_188; 
  assign _new_sip_T_1=_GEN_45&~read_mideleg; 
  assign _new_sip_T_2=wdata&read_mideleg; 
  assign _new_sip_T_3=_new_sip_T_1|_new_sip_T_2; 
  assign new_sip_ssip=_new_sip_T_3[1]; 
  assign new_satp_ppn=wdata[43:0]; 
  assign new_satp_mode=wdata[63:60]; 
  assign _T_1837=new_satp_mode==4'h0; 
  assign _T_1838=new_satp_mode==4'h8; 
  assign _T_1839=_T_1837|_T_1838; 
  assign _reg_satp_mode_T=new_satp_mode&4'h8; 
  assign _reg_mie_T_2=reg_mie&~read_mideleg; 
  assign _reg_mie_T_4=_reg_mie_T_2|_new_sip_T_2; 
  assign _GEN_242=_T_165 ? ~_reg_mepc_T_1:{24'b0,_GEN_129}; 
  assign _GEN_243=_T_166 ? wdata:{25'b0,reg_stvec}; 
  assign _reg_scause_T=wdata&64'h800000000000001f; 
  assign _GEN_248=_T_167 ? wdata:{32'b0,reg_scounteren}; 
  assign _GEN_249=_T_155 ? wdata:{32'b0,reg_mcounteren}; 
  assign _T_1842=~reg_bp_0_control_dmode|reg_debug; 
  assign _GEN_251=_T_47 ? wdata:{25'b0,reg_bp_0_address}; 
  assign _newBPC_T_2=io_rw_cmd[1] ? _T_7:64'h0; 
  assign _newBPC_T_3=_newBPC_T_2|io_rw_wdata; 
  assign _newBPC_T_8=_newBPC_T_3&~_wdata_T_5; 
  assign newBPC_action=_newBPC_T_8[12]; 
  assign newBPC_dmode=_newBPC_T_8[59]; 
  assign dMode=newBPC_dmode&reg_debug; 
  assign _GEN_252=dMode&newBPC_action; 
  assign _GEN_268=_T_1842 ? _GEN_251:{25'b0,reg_bp_0_address}; 
  assign _T_1853=_T_170&~reg_pmp_0_cfg_l; 
  assign newCfg_r=wdata[0]; 
  assign newCfg_w=wdata[1]; 
  assign newCfg_x=wdata[2]; 
  assign newCfg_a=wdata[4:3]; 
  assign newCfg_l=wdata[7]; 
  assign _reg_pmp_0_cfg_w_T=newCfg_w&newCfg_r; 
  assign _T_1857=~reg_pmp_1_cfg_a[1]&pmp_mask_base_lo_1; 
  assign _T_1858=reg_pmp_1_cfg_l&_T_1857; 
  assign _T_1859=reg_pmp_0_cfg_l|_T_1858; 
  assign _T_1861=_T_172&~_T_1859; 
  assign _GEN_323=_T_1861 ? wdata:{34'b0,reg_pmp_0_addr}; 
  assign _T_1863=_T_170&~reg_pmp_1_cfg_l; 
  assign newCfg_1_r=wdata[8]; 
  assign newCfg_1_w=wdata[9]; 
  assign newCfg_1_x=wdata[10]; 
  assign newCfg_1_a=wdata[12:11]; 
  assign newCfg_1_l=wdata[15]; 
  assign _reg_pmp_1_cfg_w_T=newCfg_1_w&newCfg_1_r; 
  assign _T_1867=~reg_pmp_2_cfg_a[1]&pmp_mask_base_lo_2; 
  assign _T_1868=reg_pmp_2_cfg_l&_T_1867; 
  assign _T_1869=reg_pmp_1_cfg_l|_T_1868; 
  assign _T_1871=_T_173&~_T_1869; 
  assign _GEN_330=_T_1871 ? wdata:{34'b0,reg_pmp_1_addr}; 
  assign _T_1873=_T_170&~reg_pmp_2_cfg_l; 
  assign newCfg_2_r=wdata[16]; 
  assign newCfg_2_w=wdata[17]; 
  assign newCfg_2_x=wdata[18]; 
  assign newCfg_2_a=wdata[20:19]; 
  assign newCfg_2_l=wdata[23]; 
  assign _reg_pmp_2_cfg_w_T=newCfg_2_w&newCfg_2_r; 
  assign _T_1877=~reg_pmp_3_cfg_a[1]&pmp_mask_base_lo_3; 
  assign _T_1878=reg_pmp_3_cfg_l&_T_1877; 
  assign _T_1879=reg_pmp_2_cfg_l|_T_1878; 
  assign _T_1881=_T_174&~_T_1879; 
  assign _GEN_337=_T_1881 ? wdata:{34'b0,reg_pmp_2_addr}; 
  assign _T_1883=_T_170&~reg_pmp_3_cfg_l; 
  assign newCfg_3_r=wdata[24]; 
  assign newCfg_3_w=wdata[25]; 
  assign newCfg_3_x=wdata[26]; 
  assign newCfg_3_a=wdata[28:27]; 
  assign newCfg_3_l=wdata[31]; 
  assign _reg_pmp_3_cfg_w_T=newCfg_3_w&newCfg_3_r; 
  assign _T_1887=~reg_pmp_4_cfg_a[1]&pmp_mask_base_lo_4; 
  assign _T_1888=reg_pmp_4_cfg_l&_T_1887; 
  assign _T_1889=reg_pmp_3_cfg_l|_T_1888; 
  assign _T_1891=_T_175&~_T_1889; 
  assign _GEN_344=_T_1891 ? wdata:{34'b0,reg_pmp_3_addr}; 
  assign _T_1893=_T_170&~reg_pmp_4_cfg_l; 
  assign newCfg_4_r=wdata[32]; 
  assign newCfg_4_w=wdata[33]; 
  assign newCfg_4_x=wdata[34]; 
  assign newCfg_4_a=wdata[36:35]; 
  assign newCfg_4_l=wdata[39]; 
  assign _reg_pmp_4_cfg_w_T=newCfg_4_w&newCfg_4_r; 
  assign _T_1897=~reg_pmp_5_cfg_a[1]&pmp_mask_base_lo_5; 
  assign _T_1898=reg_pmp_5_cfg_l&_T_1897; 
  assign _T_1899=reg_pmp_4_cfg_l|_T_1898; 
  assign _T_1901=_T_176&~_T_1899; 
  assign _GEN_351=_T_1901 ? wdata:{34'b0,reg_pmp_4_addr}; 
  assign _T_1903=_T_170&~reg_pmp_5_cfg_l; 
  assign newCfg_5_r=wdata[40]; 
  assign newCfg_5_w=wdata[41]; 
  assign newCfg_5_x=wdata[42]; 
  assign newCfg_5_a=wdata[44:43]; 
  assign newCfg_5_l=wdata[47]; 
  assign _reg_pmp_5_cfg_w_T=newCfg_5_w&newCfg_5_r; 
  assign _T_1907=~reg_pmp_6_cfg_a[1]&pmp_mask_base_lo_6; 
  assign _T_1908=reg_pmp_6_cfg_l&_T_1907; 
  assign _T_1909=reg_pmp_5_cfg_l|_T_1908; 
  assign _T_1911=_T_177&~_T_1909; 
  assign _GEN_358=_T_1911 ? wdata:{34'b0,reg_pmp_5_addr}; 
  assign _T_1913=_T_170&~reg_pmp_6_cfg_l; 
  assign newCfg_6_r=wdata[48]; 
  assign newCfg_6_w=wdata[49]; 
  assign newCfg_6_x=wdata[50]; 
  assign newCfg_6_a=wdata[52:51]; 
  assign newCfg_6_l=wdata[55]; 
  assign _reg_pmp_6_cfg_w_T=newCfg_6_w&newCfg_6_r; 
  assign _T_1917=~reg_pmp_7_cfg_a[1]&pmp_mask_base_lo_7; 
  assign _T_1918=reg_pmp_7_cfg_l&_T_1917; 
  assign _T_1919=reg_pmp_6_cfg_l|_T_1918; 
  assign _T_1921=_T_178&~_T_1919; 
  assign _GEN_365=_T_1921 ? wdata:{34'b0,reg_pmp_6_addr}; 
  assign _T_1923=_T_170&~reg_pmp_7_cfg_l; 
  assign newCfg_7_r=wdata[56]; 
  assign newCfg_7_w=wdata[57]; 
  assign newCfg_7_x=wdata[58]; 
  assign newCfg_7_a=wdata[60:59]; 
  assign newCfg_7_l=wdata[63]; 
  assign _reg_pmp_7_cfg_w_T=newCfg_7_w&newCfg_7_r; 
  assign _T_1929=reg_pmp_7_cfg_l|_T_1918; 
  assign _T_1931=_T_179&~_T_1929; 
  assign _GEN_372=_T_1931 ? wdata:{34'b0,reg_pmp_7_addr}; 
  assign _reg_custom_0_T=wdata&64'h208; 
  assign _reg_custom_0_T_2=reg_custom_0&64'hfffffffffffffdf7; 
  assign _reg_custom_0_T_3=_reg_custom_0_T|_reg_custom_0_T_2; 
  assign _GEN_385=csr_wen ? _GEN_230:_GEN_171; 
  assign _GEN_400=csr_wen ? _GEN_204:{24'b0,_GEN_136}; 
  assign _GEN_402=csr_wen ? _GEN_206:{32'b0,reg_mtvec}; 
  assign _GEN_405=csr_wen ? _GEN_209:{61'b0,reg_mcountinhibit}; 
  assign _GEN_406=csr_wen ? _GEN_210:{57'b0,_GEN_2}; 
  assign _GEN_408=csr_wen ? _GEN_212:{57'b0,_GEN_0}; 
  assign _GEN_411=csr_wen ? _GEN_219:{59'b0,_GEN_182}; 
  assign _GEN_412=csr_wen ? _GEN_220:{61'b0,reg_frm}; 
  assign _GEN_418=csr_wen ? _GEN_226:{24'b0,_GEN_120}; 
  assign _GEN_423=csr_wen ? _GEN_242:{24'b0,_GEN_129}; 
  assign _GEN_424=csr_wen ? _GEN_243:{25'b0,reg_stvec}; 
  assign _GEN_429=csr_wen ? _GEN_248:{32'b0,reg_scounteren}; 
  assign _GEN_430=csr_wen ? _GEN_249:{32'b0,reg_mcounteren}; 
  assign _GEN_432=csr_wen ? _GEN_268:{25'b0,reg_bp_0_address}; 
  assign _GEN_470=csr_wen ? _GEN_323:{34'b0,reg_pmp_0_addr}; 
  assign _GEN_477=csr_wen ? _GEN_330:{34'b0,reg_pmp_1_addr}; 
  assign _GEN_484=csr_wen ? _GEN_337:{34'b0,reg_pmp_2_addr}; 
  assign _GEN_491=csr_wen ? _GEN_344:{34'b0,reg_pmp_3_addr}; 
  assign _GEN_498=csr_wen ? _GEN_351:{34'b0,reg_pmp_4_addr}; 
  assign _GEN_505=csr_wen ? _GEN_358:{34'b0,reg_pmp_5_addr}; 
  assign _GEN_512=csr_wen ? _GEN_365:{34'b0,reg_pmp_6_addr}; 
  assign _GEN_519=csr_wen ? _GEN_372:{34'b0,reg_pmp_7_addr}; 
  assign _io_trace_0_valid_T=io_retire>1'h0; 
  assign io_rw_rdata=_io_rw_rdata_T_290|_io_rw_rdata_T_146; 
  assign io_decode_0_fp_illegal=_io_decode_0_fp_illegal_T|~reg_misa[5]; 
  assign io_decode_0_fp_csr=_io_decode_0_fp_csr_T==12'h0; 
  assign io_decode_0_read_illegal=_io_decode_0_read_illegal_T_317|_io_decode_0_read_illegal_T_320; 
  assign io_decode_0_write_illegal=&io_decode_0_csr[11:10]; 
  assign io_decode_0_write_flush=~_io_decode_0_write_flush_T_6; 
  assign io_decode_0_system_illegal=_io_decode_0_system_illegal_T_14|_io_decode_0_system_illegal_T_16; 
  assign io_csr_stall=reg_wfi|io_status_cease; 
  assign io_eret=_exception_T|insn_ret; 
  assign io_singleStep=reg_dcsr_step&~reg_debug; 
  assign io_status_debug=reg_debug; 
  assign io_status_cease=io_status_cease_r; 
  assign io_status_wfi=reg_wfi; 
  assign io_status_isa=reg_misa[31:0]; 
  assign io_status_dprv=io_status_dprv_REG; 
  assign io_status_prv=reg_mstatus_prv; 
  assign io_status_sd=_io_status_sd_T_2|_io_status_sd_T_3; 
  assign io_status_zero2=27'h0; 
  assign io_status_sxl=2'h2; 
  assign io_status_uxl=2'h2; 
  assign io_status_sd_rv32=1'h0; 
  assign io_status_zero1=8'h0; 
  assign io_status_tsr=reg_mstatus_tsr; 
  assign io_status_tw=reg_mstatus_tw; 
  assign io_status_tvm=reg_mstatus_tvm; 
  assign io_status_mxr=reg_mstatus_mxr; 
  assign io_status_sum=reg_mstatus_sum; 
  assign io_status_mprv=reg_mstatus_mprv; 
  assign io_status_xs=2'h0; 
  assign io_status_fs=reg_mstatus_fs; 
  assign io_status_mpp=reg_mstatus_mpp; 
  assign io_status_vs=2'h0; 
  assign io_status_spp=reg_mstatus_spp; 
  assign io_status_mpie=reg_mstatus_mpie; 
  assign io_status_hpie=1'h0; 
  assign io_status_spie=reg_mstatus_spie; 
  assign io_status_upie=1'h0; 
  assign io_status_mie=reg_mstatus_mie; 
  assign io_status_hie=1'h0; 
  assign io_status_sie=reg_mstatus_sie; 
  assign io_status_uie=1'h0; 
  assign io_ptbr_mode=reg_satp_mode; 
  assign io_ptbr_ppn=reg_satp_ppn; 
  assign io_evec=_GEN_172[39:0]; 
  assign io_time={value_hi_1,value_lo_1}; 
  assign io_fcsr_rm=reg_frm; 
  assign io_interrupt=_io_interrupt_T_2&~_io_interrupt_T_3; 
  assign io_interrupt_cause=64'h8000000000000000+_GEN_556; 
  assign io_bp_0_control_action=reg_bp_0_control_action; 
  assign io_bp_0_control_tmatch=reg_bp_0_control_tmatch; 
  assign io_bp_0_control_m=reg_bp_0_control_m; 
  assign io_bp_0_control_s=reg_bp_0_control_s; 
  assign io_bp_0_control_u=reg_bp_0_control_u; 
  assign io_bp_0_control_x=reg_bp_0_control_x; 
  assign io_bp_0_control_w=reg_bp_0_control_w; 
  assign io_bp_0_control_r=reg_bp_0_control_r; 
  assign io_bp_0_address=reg_bp_0_address; 
  assign io_pmp_0_cfg_l=reg_pmp_0_cfg_l; 
  assign io_pmp_0_cfg_a=reg_pmp_0_cfg_a; 
  assign io_pmp_0_cfg_x=reg_pmp_0_cfg_x; 
  assign io_pmp_0_cfg_w=reg_pmp_0_cfg_w; 
  assign io_pmp_0_cfg_r=reg_pmp_0_cfg_r; 
  assign io_pmp_0_addr=reg_pmp_0_addr; 
  assign io_pmp_0_mask=_pmp_mask_T_3[31:0]; 
  assign io_pmp_1_cfg_l=reg_pmp_1_cfg_l; 
  assign io_pmp_1_cfg_a=reg_pmp_1_cfg_a; 
  assign io_pmp_1_cfg_x=reg_pmp_1_cfg_x; 
  assign io_pmp_1_cfg_w=reg_pmp_1_cfg_w; 
  assign io_pmp_1_cfg_r=reg_pmp_1_cfg_r; 
  assign io_pmp_1_addr=reg_pmp_1_addr; 
  assign io_pmp_1_mask=_pmp_mask_T_7[31:0]; 
  assign io_pmp_2_cfg_l=reg_pmp_2_cfg_l; 
  assign io_pmp_2_cfg_a=reg_pmp_2_cfg_a; 
  assign io_pmp_2_cfg_x=reg_pmp_2_cfg_x; 
  assign io_pmp_2_cfg_w=reg_pmp_2_cfg_w; 
  assign io_pmp_2_cfg_r=reg_pmp_2_cfg_r; 
  assign io_pmp_2_addr=reg_pmp_2_addr; 
  assign io_pmp_2_mask=_pmp_mask_T_11[31:0]; 
  assign io_pmp_3_cfg_l=reg_pmp_3_cfg_l; 
  assign io_pmp_3_cfg_a=reg_pmp_3_cfg_a; 
  assign io_pmp_3_cfg_x=reg_pmp_3_cfg_x; 
  assign io_pmp_3_cfg_w=reg_pmp_3_cfg_w; 
  assign io_pmp_3_cfg_r=reg_pmp_3_cfg_r; 
  assign io_pmp_3_addr=reg_pmp_3_addr; 
  assign io_pmp_3_mask=_pmp_mask_T_15[31:0]; 
  assign io_pmp_4_cfg_l=reg_pmp_4_cfg_l; 
  assign io_pmp_4_cfg_a=reg_pmp_4_cfg_a; 
  assign io_pmp_4_cfg_x=reg_pmp_4_cfg_x; 
  assign io_pmp_4_cfg_w=reg_pmp_4_cfg_w; 
  assign io_pmp_4_cfg_r=reg_pmp_4_cfg_r; 
  assign io_pmp_4_addr=reg_pmp_4_addr; 
  assign io_pmp_4_mask=_pmp_mask_T_19[31:0]; 
  assign io_pmp_5_cfg_l=reg_pmp_5_cfg_l; 
  assign io_pmp_5_cfg_a=reg_pmp_5_cfg_a; 
  assign io_pmp_5_cfg_x=reg_pmp_5_cfg_x; 
  assign io_pmp_5_cfg_w=reg_pmp_5_cfg_w; 
  assign io_pmp_5_cfg_r=reg_pmp_5_cfg_r; 
  assign io_pmp_5_addr=reg_pmp_5_addr; 
  assign io_pmp_5_mask=_pmp_mask_T_23[31:0]; 
  assign io_pmp_6_cfg_l=reg_pmp_6_cfg_l; 
  assign io_pmp_6_cfg_a=reg_pmp_6_cfg_a; 
  assign io_pmp_6_cfg_x=reg_pmp_6_cfg_x; 
  assign io_pmp_6_cfg_w=reg_pmp_6_cfg_w; 
  assign io_pmp_6_cfg_r=reg_pmp_6_cfg_r; 
  assign io_pmp_6_addr=reg_pmp_6_addr; 
  assign io_pmp_6_mask=_pmp_mask_T_27[31:0]; 
  assign io_pmp_7_cfg_l=reg_pmp_7_cfg_l; 
  assign io_pmp_7_cfg_a=reg_pmp_7_cfg_a; 
  assign io_pmp_7_cfg_x=reg_pmp_7_cfg_x; 
  assign io_pmp_7_cfg_w=reg_pmp_7_cfg_w; 
  assign io_pmp_7_cfg_r=reg_pmp_7_cfg_r; 
  assign io_pmp_7_addr=reg_pmp_7_addr; 
  assign io_pmp_7_mask=_pmp_mask_T_31[31:0]; 
  assign io_inhibit_cycle=reg_mcountinhibit[0]; 
  assign io_trace_0_valid=_io_trace_0_valid_T|io_trace_0_exception; 
  assign io_trace_0_iaddr=io_pc; 
  assign io_trace_0_insn=io_inst_0; 
  assign io_trace_0_priv={reg_debug,reg_mstatus_prv}; 
  assign io_trace_0_exception=_exception_T|io_exception; 
  assign io_trace_0_interrupt=cause[63]; 
  assign io_trace_0_cause=insn_call ? {60'b0,_cause_T_1}:_cause_T_2; 
  assign io_trace_0_tval=io_tval; 
  assign io_customCSRs_0_value=reg_custom_0; 
  assign CSRFile_cov_read_addr=CSRFile_state; 
  assign CSRFile_cov_read_data=CSRFile_cov[CSRFile_cov_read_addr]; 
  assign CSRFile_cov_write_data=1'h1; 
  assign CSRFile_cov_write_addr=CSRFile_state; 
  assign CSRFile_cov_write_mask=1'h1; 
  assign CSRFile_cov_write_en=1'h1; 
  assign reg_pmp_5_cfg_l_shl={reg_pmp_5_cfg_l,19'h0}; 
  assign reg_pmp_5_cfg_l_pad=reg_pmp_5_cfg_l_shl; 
  assign reg_debug_shl={reg_debug,1'h0}; 
  assign reg_debug_pad={18'h0,reg_debug_shl}; 
  assign reg_mstatus_sie_shl={reg_mstatus_sie,16'h0}; 
  assign reg_mstatus_sie_pad={3'h0,reg_mstatus_sie_shl}; 
  assign reg_dcsr_prv_shl={reg_dcsr_prv,13'h0}; 
  assign reg_dcsr_prv_pad={5'h0,reg_dcsr_prv_shl}; 
  assign reg_mcountinhibit_shl={reg_mcountinhibit,15'h0}; 
  assign reg_mcountinhibit_pad={2'h0,reg_mcountinhibit_shl}; 
  assign reg_unmie_shl={reg_unmie,2'h0}; 
  assign reg_unmie_pad={17'h0,reg_unmie_shl}; 
  assign reg_pmp_7_cfg_a_shl={reg_pmp_7_cfg_a,13'h0}; 
  assign reg_pmp_7_cfg_a_pad={5'h0,reg_pmp_7_cfg_a_shl}; 
  assign reg_mstatus_mpp_shl=reg_mstatus_mpp; 
  assign reg_mstatus_mpp_pad={18'h0,reg_mstatus_mpp_shl}; 
  assign reg_pmp_2_cfg_l_shl={reg_pmp_2_cfg_l,6'h0}; 
  assign reg_pmp_2_cfg_l_pad={13'h0,reg_pmp_2_cfg_l_shl}; 
  assign reg_pmp_1_cfg_l_shl={reg_pmp_1_cfg_l,18'h0}; 
  assign reg_pmp_1_cfg_l_pad={1'h0,reg_pmp_1_cfg_l_shl}; 
  assign reg_mip_seip_shl={reg_mip_seip,9'h0}; 
  assign reg_mip_seip_pad={10'h0,reg_mip_seip_shl}; 
  assign reg_rnmie_shl={reg_rnmie,1'h0}; 
  assign reg_rnmie_pad={18'h0,reg_rnmie_shl}; 
  assign reg_mip_ssip_shl={reg_mip_ssip,10'h0}; 
  assign reg_mip_ssip_pad={9'h0,reg_mip_ssip_shl}; 
  assign reg_bp_0_control_dmode_shl={reg_bp_0_control_dmode,2'h0}; 
  assign reg_bp_0_control_dmode_pad={17'h0,reg_bp_0_control_dmode_shl}; 
  assign reg_pmp_4_cfg_l_shl={reg_pmp_4_cfg_l,11'h0}; 
  assign reg_pmp_4_cfg_l_pad={8'h0,reg_pmp_4_cfg_l_shl}; 
  assign reg_dcsr_ebreaks_shl={reg_dcsr_ebreaks,1'h0}; 
  assign reg_dcsr_ebreaks_pad={18'h0,reg_dcsr_ebreaks_shl}; 
  assign reg_pmp_6_cfg_l_shl={reg_pmp_6_cfg_l,13'h0}; 
  assign reg_pmp_6_cfg_l_pad={6'h0,reg_pmp_6_cfg_l_shl}; 
  assign reg_mstatus_prv_shl={reg_mstatus_prv,2'h0}; 
  assign reg_mstatus_prv_pad={16'h0,reg_mstatus_prv_shl}; 
  assign reg_dcsr_ebreakm_shl={reg_dcsr_ebreakm,8'h0}; 
  assign reg_dcsr_ebreakm_pad={11'h0,reg_dcsr_ebreakm_shl}; 
  assign reg_pmp_7_cfg_l_shl=reg_pmp_7_cfg_l; 
  assign reg_pmp_7_cfg_l_pad={19'h0,reg_pmp_7_cfg_l_shl}; 
  assign reg_pmp_0_cfg_l_shl={reg_pmp_0_cfg_l,18'h0}; 
  assign reg_pmp_0_cfg_l_pad={1'h0,reg_pmp_0_cfg_l_shl}; 
  assign reg_pmp_3_cfg_l_shl={reg_pmp_3_cfg_l,1'h0}; 
  assign reg_pmp_3_cfg_l_pad={18'h0,reg_pmp_3_cfg_l_shl}; 
  assign reg_mstatus_spp_shl={reg_mstatus_spp,13'h0}; 
  assign reg_mstatus_spp_pad={6'h0,reg_mstatus_spp_shl}; 
  assign reg_mip_stip_shl={reg_mip_stip,12'h0}; 
  assign reg_mip_stip_pad={7'h0,reg_mip_stip_shl}; 
  assign reg_dcsr_ebreaku_shl={reg_dcsr_ebreaku,13'h0}; 
  assign reg_dcsr_ebreaku_pad={6'h0,reg_dcsr_ebreaku_shl}; 
  assign reg_mstatus_mprv_shl=reg_mstatus_mprv; 
  assign reg_mstatus_mprv_pad={19'h0,reg_mstatus_mprv_shl}; 
  assign reg_singleStepped_shl={reg_singleStepped,13'h0}; 
  assign reg_singleStepped_pad={6'h0,reg_singleStepped_shl}; 
  assign reg_mstatus_mie_shl={reg_mstatus_mie,11'h0}; 
  assign reg_mstatus_mie_pad={8'h0,reg_mstatus_mie_shl}; 
  assign CSRFile_xor16=reg_debug_pad^reg_mstatus_sie_pad; 
  assign CSRFile_xor7=reg_pmp_5_cfg_l_pad^CSRFile_xor16; 
  assign CSRFile_xor17=reg_dcsr_prv_pad^reg_mcountinhibit_pad; 
  assign CSRFile_xor18=reg_unmie_pad^reg_pmp_7_cfg_a_pad; 
  assign CSRFile_xor8=CSRFile_xor17^CSRFile_xor18; 
  assign CSRFile_xor3=CSRFile_xor7^CSRFile_xor8; 
  assign CSRFile_xor20=reg_pmp_2_cfg_l_pad^reg_pmp_1_cfg_l_pad; 
  assign CSRFile_xor9=reg_mstatus_mpp_pad^CSRFile_xor20; 
  assign CSRFile_xor21=reg_mip_seip_pad^reg_rnmie_pad; 
  assign CSRFile_xor22=reg_mip_ssip_pad^reg_bp_0_control_dmode_pad; 
  assign CSRFile_xor10=CSRFile_xor21^CSRFile_xor22; 
  assign CSRFile_xor4=CSRFile_xor9^CSRFile_xor10; 
  assign CSRFile_xor1=CSRFile_xor3^CSRFile_xor4; 
  assign CSRFile_xor24=reg_dcsr_ebreaks_pad^reg_pmp_6_cfg_l_pad; 
  assign CSRFile_xor11=reg_pmp_4_cfg_l_pad^CSRFile_xor24; 
  assign CSRFile_xor25=reg_mstatus_prv_pad^reg_dcsr_ebreakm_pad; 
  assign CSRFile_xor26=reg_pmp_7_cfg_l_pad^reg_pmp_0_cfg_l_pad; 
  assign CSRFile_xor12=CSRFile_xor25^CSRFile_xor26; 
  assign CSRFile_xor5=CSRFile_xor11^CSRFile_xor12; 
  assign CSRFile_xor28=reg_mstatus_spp_pad^reg_mip_stip_pad; 
  assign CSRFile_xor13=reg_pmp_3_cfg_l_pad^CSRFile_xor28; 
  assign CSRFile_xor29=reg_dcsr_ebreaku_pad^reg_mstatus_mprv_pad; 
  assign CSRFile_xor30=reg_singleStepped_pad^reg_mstatus_mie_pad; 
  assign CSRFile_xor14=CSRFile_xor29^CSRFile_xor30; 
  assign CSRFile_xor6=CSRFile_xor13^CSRFile_xor14; 
  assign CSRFile_xor2=CSRFile_xor5^CSRFile_xor6; 
  assign CSRFile_xor0=CSRFile_xor1^CSRFile_xor2; 
  assign io_covSum=CSRFile_covSum; 
  assign stopEn0=~_T_252; 
  assign stopEn1=~_T_274; 
  assign CSRFile_or0=stopEn0|stopEn1; 
  assign metaAssert=CSRFile_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              reg_mstatus_prv <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_prv <=2'h3;
               end 
             else 
               if (_reg_mstatus_prv_T)
                  begin 
                    reg_mstatus_prv <=2'h0;
                  end 
                else 
                  if (insn_ret)
                     begin 
                       if (~io_rw_addr[9])
                          begin 
                            reg_mstatus_prv <={1'b0,reg_mstatus_spp};
                          end 
                        else 
                          if (_T_406)
                             begin 
                               reg_mstatus_prv <=reg_dcsr_prv;
                             end 
                           else 
                             begin 
                               reg_mstatus_prv <=reg_mstatus_mpp;
                             end 
                     end 
                   else 
                     if (exception)
                        begin 
                          if (trapToDebug)
                             begin 
                               if (~reg_debug)
                                  begin 
                                    reg_mstatus_prv <=2'h3;
                                  end 
                             end 
                           else 
                             if (_T_279)
                                begin 
                                  reg_mstatus_prv <=2'h1;
                                end 
                              else 
                                begin 
                                  reg_mstatus_prv <=2'h3;
                                end 
                        end 
         if (metaReset)
            begin 
              reg_mstatus_tsr <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_tsr <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_50)
                       begin 
                         reg_mstatus_tsr <=new_mstatus_tsr;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_mstatus_tw <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_tw <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_50)
                       begin 
                         reg_mstatus_tw <=new_mstatus_tw;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_mstatus_tvm <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_tvm <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_50)
                       begin 
                         reg_mstatus_tvm <=new_mstatus_tvm;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_mstatus_mxr <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_mxr <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_158)
                       begin 
                         reg_mstatus_mxr <=new_mstatus_mxr;
                       end 
                     else 
                       if (_T_50)
                          begin 
                            reg_mstatus_mxr <=new_mstatus_mxr;
                          end 
                  end 
         if (metaReset)
            begin 
              reg_mstatus_sum <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_sum <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_158)
                       begin 
                         reg_mstatus_sum <=new_mstatus_sum;
                       end 
                     else 
                       if (_T_50)
                          begin 
                            reg_mstatus_sum <=new_mstatus_sum;
                          end 
                  end 
         if (metaReset)
            begin 
              reg_mstatus_mprv <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_mprv <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_50)
                       begin 
                         reg_mstatus_mprv <=new_mstatus_mprv;
                       end 
                     else 
                       if (insn_ret)
                          begin 
                            if (_T_412)
                               begin 
                                 reg_mstatus_mprv <=1'h0;
                               end 
                          end 
                  end 
                else 
                  if (insn_ret)
                     begin 
                       if (_T_412)
                          begin 
                            reg_mstatus_mprv <=1'h0;
                          end 
                     end 
         if (metaReset)
            begin 
              reg_mstatus_fs <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_fs <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_158)
                       begin 
                         if (_reg_mstatus_fs_T)
                            begin 
                              reg_mstatus_fs <=2'h3;
                            end 
                          else 
                            begin 
                              reg_mstatus_fs <=2'h0;
                            end 
                       end 
                     else 
                       if (_T_50)
                          begin 
                            if (_reg_mstatus_fs_T)
                               begin 
                                 reg_mstatus_fs <=2'h3;
                               end 
                             else 
                               begin 
                                 reg_mstatus_fs <=2'h0;
                               end 
                          end 
                  end 
         if (metaReset)
            begin 
              reg_mstatus_mpp <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_mpp <=2'h3;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_50)
                       begin 
                         if (_reg_mstatus_mpp_T_2)
                            begin 
                              reg_mstatus_mpp <=2'h0;
                            end 
                          else 
                            begin 
                              reg_mstatus_mpp <=new_mstatus_mpp;
                            end 
                       end 
                     else 
                       if (insn_ret)
                          begin 
                            if (~io_rw_addr[9])
                               begin 
                                 if (exception)
                                    begin 
                                      if (!(trapToDebug))
                                         begin 
                                           if (!(_T_279))
                                              begin 
                                                reg_mstatus_mpp <=reg_mstatus_prv;
                                              end 
                                         end 
                                    end 
                               end 
                             else 
                               if (_T_406)
                                  begin 
                                    if (exception)
                                       begin 
                                         if (!(trapToDebug))
                                            begin 
                                              if (!(_T_279))
                                                 begin 
                                                   reg_mstatus_mpp <=reg_mstatus_prv;
                                                 end 
                                            end 
                                       end 
                                  end 
                                else 
                                  begin 
                                    reg_mstatus_mpp <=2'h0;
                                  end 
                          end 
                        else 
                          if (exception)
                             begin 
                               if (!(trapToDebug))
                                  begin 
                                    if (!(_T_279))
                                       begin 
                                         reg_mstatus_mpp <=reg_mstatus_prv;
                                       end 
                                  end 
                             end 
                  end 
                else 
                  if (insn_ret)
                     begin 
                       if (~io_rw_addr[9])
                          begin 
                            if (exception)
                               begin 
                                 if (!(trapToDebug))
                                    begin 
                                      if (!(_T_279))
                                         begin 
                                           reg_mstatus_mpp <=reg_mstatus_prv;
                                         end 
                                    end 
                               end 
                          end 
                        else 
                          if (_T_406)
                             begin 
                               reg_mstatus_mpp <=_GEN_140;
                             end 
                           else 
                             begin 
                               reg_mstatus_mpp <=2'h0;
                             end 
                     end 
                   else 
                     begin 
                       reg_mstatus_mpp <=_GEN_140;
                     end 
         if (metaReset)
            begin 
              reg_mstatus_spp <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_spp <=1'h0;
               end 
             else 
               begin 
                 reg_mstatus_spp <=_GEN_385[0];
               end 
         if (metaReset)
            begin 
              reg_mstatus_mpie <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_mpie <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_50)
                       begin 
                         reg_mstatus_mpie <=new_mstatus_mpie;
                       end 
                     else 
                       if (insn_ret)
                          begin 
                            if (~io_rw_addr[9])
                               begin 
                                 if (exception)
                                    begin 
                                      if (!(trapToDebug))
                                         begin 
                                           if (!(_T_279))
                                              begin 
                                                reg_mstatus_mpie <=reg_mstatus_mie;
                                              end 
                                         end 
                                    end 
                               end 
                             else 
                               if (_T_406)
                                  begin 
                                    if (exception)
                                       begin 
                                         if (!(trapToDebug))
                                            begin 
                                              if (!(_T_279))
                                                 begin 
                                                   reg_mstatus_mpie <=reg_mstatus_mie;
                                                 end 
                                            end 
                                       end 
                                  end 
                                else 
                                  begin 
                                    reg_mstatus_mpie <=1'h1;
                                  end 
                          end 
                        else 
                          if (exception)
                             begin 
                               if (!(trapToDebug))
                                  begin 
                                    if (!(_T_279))
                                       begin 
                                         reg_mstatus_mpie <=reg_mstatus_mie;
                                       end 
                                  end 
                             end 
                  end 
                else 
                  if (insn_ret)
                     begin 
                       if (~io_rw_addr[9])
                          begin 
                            if (exception)
                               begin 
                                 if (!(trapToDebug))
                                    begin 
                                      if (!(_T_279))
                                         begin 
                                           reg_mstatus_mpie <=reg_mstatus_mie;
                                         end 
                                    end 
                               end 
                          end 
                        else 
                          if (_T_406)
                             begin 
                               reg_mstatus_mpie <=_GEN_139;
                             end 
                           else 
                             begin 
                               reg_mstatus_mpie <=1'h1;
                             end 
                     end 
                   else 
                     begin 
                       reg_mstatus_mpie <=_GEN_139;
                     end 
         if (metaReset)
            begin 
              reg_mstatus_spie <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_spie <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_158)
                       begin 
                         reg_mstatus_spie <=new_mstatus_spie;
                       end 
                     else 
                       if (_T_50)
                          begin 
                            reg_mstatus_spie <=new_mstatus_spie;
                          end 
                        else 
                          if (insn_ret)
                             begin 
                               reg_mstatus_spie <=_GEN_158;
                             end 
                           else 
                             if (exception)
                                begin 
                                  if (!(trapToDebug))
                                     begin 
                                       if (_T_279)
                                          begin 
                                            reg_mstatus_spie <=reg_mstatus_sie;
                                          end 
                                     end 
                                end 
                  end 
                else 
                  if (insn_ret)
                     begin 
                       reg_mstatus_spie <=_GEN_158;
                     end 
                   else 
                     if (exception)
                        begin 
                          if (!(trapToDebug))
                             begin 
                               if (_T_279)
                                  begin 
                                    reg_mstatus_spie <=reg_mstatus_sie;
                                  end 
                             end 
                        end 
         if (metaReset)
            begin 
              reg_mstatus_mie <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_mie <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_50)
                       begin 
                         reg_mstatus_mie <=new_mstatus_mie;
                       end 
                     else 
                       if (insn_ret)
                          begin 
                            if (~io_rw_addr[9])
                               begin 
                                 if (exception)
                                    begin 
                                      if (!(trapToDebug))
                                         begin 
                                           reg_mstatus_mie <=_GEN_76;
                                         end 
                                    end 
                               end 
                             else 
                               if (_T_406)
                                  begin 
                                    if (exception)
                                       begin 
                                         if (!(trapToDebug))
                                            begin 
                                              reg_mstatus_mie <=_GEN_76;
                                            end 
                                       end 
                                  end 
                                else 
                                  begin 
                                    reg_mstatus_mie <=reg_mstatus_mpie;
                                  end 
                          end 
                        else 
                          if (exception)
                             begin 
                               if (!(trapToDebug))
                                  begin 
                                    reg_mstatus_mie <=_GEN_76;
                                  end 
                             end 
                  end 
                else 
                  if (insn_ret)
                     begin 
                       if (~io_rw_addr[9])
                          begin 
                            if (exception)
                               begin 
                                 if (!(trapToDebug))
                                    begin 
                                      reg_mstatus_mie <=_GEN_76;
                                    end 
                               end 
                          end 
                        else 
                          if (_T_406)
                             begin 
                               reg_mstatus_mie <=_GEN_141;
                             end 
                           else 
                             begin 
                               reg_mstatus_mie <=reg_mstatus_mpie;
                             end 
                     end 
                   else 
                     begin 
                       reg_mstatus_mie <=_GEN_141;
                     end 
         if (metaReset)
            begin 
              reg_mstatus_sie <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mstatus_sie <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_158)
                       begin 
                         reg_mstatus_sie <=new_mstatus_sie;
                       end 
                     else 
                       if (_T_50)
                          begin 
                            reg_mstatus_sie <=new_mstatus_sie;
                          end 
                        else 
                          if (insn_ret)
                             begin 
                               if (~io_rw_addr[9])
                                  begin 
                                    reg_mstatus_sie <=reg_mstatus_spie;
                                  end 
                                else 
                                  if (exception)
                                     begin 
                                       if (!(trapToDebug))
                                          begin 
                                            if (_T_279)
                                               begin 
                                                 reg_mstatus_sie <=1'h0;
                                               end 
                                          end 
                                     end 
                             end 
                           else 
                             if (exception)
                                begin 
                                  if (!(trapToDebug))
                                     begin 
                                       if (_T_279)
                                          begin 
                                            reg_mstatus_sie <=1'h0;
                                          end 
                                     end 
                                end 
                  end 
                else 
                  if (insn_ret)
                     begin 
                       if (~io_rw_addr[9])
                          begin 
                            reg_mstatus_sie <=reg_mstatus_spie;
                          end 
                        else 
                          if (exception)
                             begin 
                               if (!(trapToDebug))
                                  begin 
                                    if (_T_279)
                                       begin 
                                         reg_mstatus_sie <=1'h0;
                                       end 
                                  end 
                             end 
                     end 
                   else 
                     if (exception)
                        begin 
                          if (!(trapToDebug))
                             begin 
                               if (_T_279)
                                  begin 
                                    reg_mstatus_sie <=1'h0;
                                  end 
                             end 
                        end 
         if (metaReset)
            begin 
              reg_dcsr_prv <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_dcsr_prv <=2'h3;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_59)
                       begin 
                         if (_reg_dcsr_prv_T)
                            begin 
                              reg_dcsr_prv <=2'h0;
                            end 
                          else 
                            begin 
                              reg_dcsr_prv <=new_dcsr_prv;
                            end 
                       end 
                     else 
                       if (exception)
                          begin 
                            if (trapToDebug)
                               begin 
                                 if (~reg_debug)
                                    begin 
                                      reg_dcsr_prv <=reg_mstatus_prv;
                                    end 
                               end 
                          end 
                  end 
                else 
                  if (exception)
                     begin 
                       if (trapToDebug)
                          begin 
                            if (~reg_debug)
                               begin 
                                 reg_dcsr_prv <=reg_mstatus_prv;
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              reg_singleStepped <=1'h0;
            end 
          else 
            if (~io_singleStep)
               begin 
                 reg_singleStepped <=1'h0;
               end 
             else 
               begin 
                 reg_singleStepped <=_GEN_50;
               end 
         if (metaReset)
            begin 
              reg_dcsr_ebreakm <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_dcsr_ebreakm <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_59)
                       begin 
                         reg_dcsr_ebreakm <=new_dcsr_ebreakm;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_dcsr_ebreaks <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_dcsr_ebreaks <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_59)
                       begin 
                         reg_dcsr_ebreaks <=new_dcsr_ebreaks;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_dcsr_ebreaku <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_dcsr_ebreaku <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_59)
                       begin 
                         reg_dcsr_ebreaku <=new_dcsr_ebreaku;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_debug <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_debug <=1'h0;
               end 
             else 
               if (insn_ret)
                  begin 
                    if (~io_rw_addr[9])
                       begin 
                         if (exception)
                            begin 
                              if (trapToDebug)
                                 begin 
                                   reg_debug <=_GEN_52;
                                 end 
                            end 
                       end 
                     else 
                       if (_T_406)
                          begin 
                            reg_debug <=1'h0;
                          end 
                        else 
                          if (exception)
                             begin 
                               if (trapToDebug)
                                  begin 
                                    reg_debug <=_GEN_52;
                                  end 
                             end 
                  end 
                else 
                  if (exception)
                     begin 
                       if (trapToDebug)
                          begin 
                            reg_debug <=_GEN_52;
                          end 
                     end 
         if (metaReset)
            begin 
              reg_rnmie <=1'h0;
            end 
          else 
            begin 
              reg_rnmie <=reset|reg_rnmie;
            end 
         if (metaReset)
            begin 
              reg_unmie <=1'h0;
            end 
          else 
            begin 
              reg_unmie <=reset|reg_unmie;
            end 
         if (metaReset)
            begin 
              reg_mideleg <=64'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_168)
                    begin 
                      reg_mideleg <=wdata;
                    end 
               end 
         if (metaReset)
            begin 
              reg_medeleg <=64'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_169)
                    begin 
                      reg_medeleg <=wdata;
                    end 
               end 
         if (metaReset)
            begin 
              reg_dcsr_cause <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_dcsr_cause <=3'h0;
               end 
             else 
               if (exception)
                  begin 
                    if (trapToDebug)
                       begin 
                         if (~reg_debug)
                            begin 
                              if (reg_singleStepped)
                                 begin 
                                   reg_dcsr_cause <=3'h4;
                                 end 
                               else 
                                 begin 
                                   reg_dcsr_cause <={1'b0,_reg_dcsr_cause_T_1};
                                 end 
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_dcsr_step <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_dcsr_step <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_59)
                       begin 
                         reg_dcsr_step <=new_dcsr_step;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_dpc <=40'h0;
            end 
          else 
            begin 
              reg_dpc <=_GEN_418[39:0];
            end 
         if (metaReset)
            begin 
              reg_dscratch <=64'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_61)
                    begin 
                      reg_dscratch <=wdata;
                    end 
               end 
         if (metaReset)
            begin 
              reg_bp_0_control_dmode <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_bp_0_control_dmode <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1842)
                       begin 
                         if (_T_46)
                            begin 
                              reg_bp_0_control_dmode <=dMode;
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_bp_0_control_action <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_bp_0_control_action <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1842)
                       begin 
                         if (_T_46)
                            begin 
                              reg_bp_0_control_action <=_GEN_252;
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_bp_0_control_tmatch <=2'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1842)
                    begin 
                      if (_T_46)
                         begin 
                           reg_bp_0_control_tmatch <=wdata[8:7];
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              reg_bp_0_control_m <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1842)
                    begin 
                      if (_T_46)
                         begin 
                           reg_bp_0_control_m <=wdata[6];
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              reg_bp_0_control_s <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1842)
                    begin 
                      if (_T_46)
                         begin 
                           reg_bp_0_control_s <=wdata[4];
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              reg_bp_0_control_u <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1842)
                    begin 
                      if (_T_46)
                         begin 
                           reg_bp_0_control_u <=wdata[3];
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              reg_bp_0_control_x <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_bp_0_control_x <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1842)
                       begin 
                         if (_T_46)
                            begin 
                              reg_bp_0_control_x <=wdata[2];
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_bp_0_control_w <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_bp_0_control_w <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1842)
                       begin 
                         if (_T_46)
                            begin 
                              reg_bp_0_control_w <=wdata[1];
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_bp_0_control_r <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_bp_0_control_r <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1842)
                       begin 
                         if (_T_46)
                            begin 
                              reg_bp_0_control_r <=wdata[0];
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_bp_0_address <=39'h0;
            end 
          else 
            begin 
              reg_bp_0_address <=_GEN_432[38:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_0_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_0_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1853)
                       begin 
                         reg_pmp_0_cfg_l <=newCfg_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_0_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_0_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1853)
                       begin 
                         reg_pmp_0_cfg_a <=newCfg_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_0_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1853)
                    begin 
                      reg_pmp_0_cfg_x <=newCfg_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_0_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1853)
                    begin 
                      reg_pmp_0_cfg_w <=_reg_pmp_0_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_0_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1853)
                    begin 
                      reg_pmp_0_cfg_r <=newCfg_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_0_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_0_addr <=_GEN_470[29:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_1_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_1_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1863)
                       begin 
                         reg_pmp_1_cfg_l <=newCfg_1_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_1_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_1_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1863)
                       begin 
                         reg_pmp_1_cfg_a <=newCfg_1_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_1_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1863)
                    begin 
                      reg_pmp_1_cfg_x <=newCfg_1_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_1_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1863)
                    begin 
                      reg_pmp_1_cfg_w <=_reg_pmp_1_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_1_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1863)
                    begin 
                      reg_pmp_1_cfg_r <=newCfg_1_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_1_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_1_addr <=_GEN_477[29:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_2_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_2_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1873)
                       begin 
                         reg_pmp_2_cfg_l <=newCfg_2_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_2_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_2_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1873)
                       begin 
                         reg_pmp_2_cfg_a <=newCfg_2_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_2_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1873)
                    begin 
                      reg_pmp_2_cfg_x <=newCfg_2_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_2_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1873)
                    begin 
                      reg_pmp_2_cfg_w <=_reg_pmp_2_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_2_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1873)
                    begin 
                      reg_pmp_2_cfg_r <=newCfg_2_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_2_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_2_addr <=_GEN_484[29:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_3_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_3_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1883)
                       begin 
                         reg_pmp_3_cfg_l <=newCfg_3_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_3_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_3_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1883)
                       begin 
                         reg_pmp_3_cfg_a <=newCfg_3_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_3_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1883)
                    begin 
                      reg_pmp_3_cfg_x <=newCfg_3_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_3_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1883)
                    begin 
                      reg_pmp_3_cfg_w <=_reg_pmp_3_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_3_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1883)
                    begin 
                      reg_pmp_3_cfg_r <=newCfg_3_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_3_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_3_addr <=_GEN_491[29:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_4_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_4_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1893)
                       begin 
                         reg_pmp_4_cfg_l <=newCfg_4_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_4_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_4_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1893)
                       begin 
                         reg_pmp_4_cfg_a <=newCfg_4_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_4_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1893)
                    begin 
                      reg_pmp_4_cfg_x <=newCfg_4_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_4_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1893)
                    begin 
                      reg_pmp_4_cfg_w <=_reg_pmp_4_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_4_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1893)
                    begin 
                      reg_pmp_4_cfg_r <=newCfg_4_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_4_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_4_addr <=_GEN_498[29:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_5_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_5_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1903)
                       begin 
                         reg_pmp_5_cfg_l <=newCfg_5_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_5_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_5_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1903)
                       begin 
                         reg_pmp_5_cfg_a <=newCfg_5_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_5_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1903)
                    begin 
                      reg_pmp_5_cfg_x <=newCfg_5_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_5_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1903)
                    begin 
                      reg_pmp_5_cfg_w <=_reg_pmp_5_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_5_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1903)
                    begin 
                      reg_pmp_5_cfg_r <=newCfg_5_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_5_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_5_addr <=_GEN_505[29:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_6_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_6_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1913)
                       begin 
                         reg_pmp_6_cfg_l <=newCfg_6_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_6_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_6_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1913)
                       begin 
                         reg_pmp_6_cfg_a <=newCfg_6_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_6_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1913)
                    begin 
                      reg_pmp_6_cfg_x <=newCfg_6_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_6_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1913)
                    begin 
                      reg_pmp_6_cfg_w <=_reg_pmp_6_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_6_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1913)
                    begin 
                      reg_pmp_6_cfg_r <=newCfg_6_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_6_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_6_addr <=_GEN_512[29:0];
            end 
         if (metaReset)
            begin 
              reg_pmp_7_cfg_l <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_7_cfg_l <=1'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1923)
                       begin 
                         reg_pmp_7_cfg_l <=newCfg_7_l;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_7_cfg_a <=2'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_pmp_7_cfg_a <=2'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_1923)
                       begin 
                         reg_pmp_7_cfg_a <=newCfg_7_a;
                       end 
                  end 
         if (metaReset)
            begin 
              reg_pmp_7_cfg_x <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1923)
                    begin 
                      reg_pmp_7_cfg_x <=newCfg_7_x;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_7_cfg_w <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1923)
                    begin 
                      reg_pmp_7_cfg_w <=_reg_pmp_7_cfg_w_T;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_7_cfg_r <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_1923)
                    begin 
                      reg_pmp_7_cfg_r <=newCfg_7_r;
                    end 
               end 
         if (metaReset)
            begin 
              reg_pmp_7_addr <=30'h0;
            end 
          else 
            begin 
              reg_pmp_7_addr <=_GEN_519[29:0];
            end 
         if (metaReset)
            begin 
              reg_mie <=64'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_160)
                    begin 
                      reg_mie <=_reg_mie_T_4;
                    end 
                  else 
                    if (_T_53)
                       begin 
                         reg_mie <=_reg_mie_T;
                       end 
               end 
         if (metaReset)
            begin 
              reg_mip_seip <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_52)
                    begin 
                      reg_mip_seip <=new_mip_seip;
                    end 
               end 
         if (metaReset)
            begin 
              reg_mip_stip <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_52)
                    begin 
                      reg_mip_stip <=new_mip_stip;
                    end 
               end 
         if (metaReset)
            begin 
              reg_mip_ssip <=1'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_159)
                    begin 
                      reg_mip_ssip <=new_sip_ssip;
                    end 
                  else 
                    if (_T_52)
                       begin 
                         reg_mip_ssip <=new_mip_ssip;
                       end 
               end 
         if (metaReset)
            begin 
              reg_mepc <=40'h0;
            end 
          else 
            begin 
              reg_mepc <=_GEN_400[39:0];
            end 
         if (metaReset)
            begin 
              reg_mcause <=64'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mcause <=64'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_57)
                       begin 
                         reg_mcause <=_reg_mcause_T;
                       end 
                     else 
                       if (exception)
                          begin 
                            if (!(trapToDebug))
                               begin 
                                 if (!(_T_279))
                                    begin 
                                      if (insn_call)
                                         begin 
                                           reg_mcause <={60'b0,_cause_T_1};
                                         end 
                                       else 
                                         if (insn_break)
                                            begin 
                                              reg_mcause <=64'h3;
                                            end 
                                          else 
                                            begin 
                                              reg_mcause <=io_cause;
                                            end 
                                    end 
                               end 
                          end 
                  end 
                else 
                  if (exception)
                     begin 
                       if (!(trapToDebug))
                          begin 
                            if (!(_T_279))
                               begin 
                                 if (insn_call)
                                    begin 
                                      reg_mcause <={60'b0,_cause_T_1};
                                    end 
                                  else 
                                    if (insn_break)
                                       begin 
                                         reg_mcause <=64'h3;
                                       end 
                                     else 
                                       begin 
                                         reg_mcause <=io_cause;
                                       end 
                               end 
                          end 
                     end 
         if (metaReset)
            begin 
              reg_mtval <=40'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_56)
                    begin 
                      reg_mtval <=wdata[39:0];
                    end 
                  else 
                    if (exception)
                       begin 
                         if (!(trapToDebug))
                            begin 
                              if (!(_T_279))
                                 begin 
                                   reg_mtval <=io_tval;
                                 end 
                            end 
                       end 
               end 
             else 
               if (exception)
                  begin 
                    if (!(trapToDebug))
                       begin 
                         if (!(_T_279))
                            begin 
                              reg_mtval <=io_tval;
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_mscratch <=64'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_54)
                    begin 
                      reg_mscratch <=wdata;
                    end 
               end 
         if (metaReset)
            begin 
              reg_mtvec <=32'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mtvec <=32'h0;
               end 
             else 
               begin 
                 reg_mtvec <=_GEN_402[31:0];
               end 
         if (metaReset)
            begin 
              reg_mcounteren <=32'h0;
            end 
          else 
            begin 
              reg_mcounteren <=_GEN_430[31:0];
            end 
         if (metaReset)
            begin 
              reg_scounteren <=32'h0;
            end 
          else 
            begin 
              reg_scounteren <=_GEN_429[31:0];
            end 
         if (metaReset)
            begin 
              reg_sepc <=40'h0;
            end 
          else 
            begin 
              reg_sepc <=_GEN_423[39:0];
            end 
         if (metaReset)
            begin 
              reg_scause <=64'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_162)
                    begin 
                      reg_scause <=_reg_scause_T;
                    end 
                  else 
                    if (exception)
                       begin 
                         if (!(trapToDebug))
                            begin 
                              if (_T_279)
                                 begin 
                                   if (insn_call)
                                      begin 
                                        reg_scause <={60'b0,_cause_T_1};
                                      end 
                                    else 
                                      if (insn_break)
                                         begin 
                                           reg_scause <=64'h3;
                                         end 
                                       else 
                                         begin 
                                           reg_scause <=io_cause;
                                         end 
                                 end 
                            end 
                       end 
               end 
             else 
               if (exception)
                  begin 
                    if (!(trapToDebug))
                       begin 
                         if (_T_279)
                            begin 
                              if (insn_call)
                                 begin 
                                   reg_scause <={60'b0,_cause_T_1};
                                 end 
                               else 
                                 if (insn_break)
                                    begin 
                                      reg_scause <=64'h3;
                                    end 
                                  else 
                                    begin 
                                      reg_scause <=io_cause;
                                    end 
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_stval <=40'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_163)
                    begin 
                      reg_stval <=wdata[39:0];
                    end 
                  else 
                    if (exception)
                       begin 
                         if (!(trapToDebug))
                            begin 
                              if (_T_279)
                                 begin 
                                   reg_stval <=io_tval;
                                 end 
                            end 
                       end 
               end 
             else 
               if (exception)
                  begin 
                    if (!(trapToDebug))
                       begin 
                         if (_T_279)
                            begin 
                              reg_stval <=io_tval;
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_sscratch <=64'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_161)
                    begin 
                      reg_sscratch <=wdata;
                    end 
               end 
         if (metaReset)
            begin 
              reg_stvec <=39'h0;
            end 
          else 
            begin 
              reg_stvec <=_GEN_424[38:0];
            end 
         if (metaReset)
            begin 
              reg_satp_mode <=4'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_164)
                    begin 
                      if (_T_1839)
                         begin 
                           reg_satp_mode <=_reg_satp_mode_T;
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              reg_satp_ppn <=44'h0;
            end 
          else 
            if (csr_wen)
               begin 
                 if (_T_164)
                    begin 
                      if (_T_1839)
                         begin 
                           reg_satp_ppn <={24'b0,new_satp_ppn[19:0]};
                         end 
                    end 
               end 
         if (metaReset)
            begin 
              reg_fflags <=5'h0;
            end 
          else 
            begin 
              reg_fflags <=_GEN_411[4:0];
            end 
         if (metaReset)
            begin 
              reg_frm <=3'h0;
            end 
          else 
            begin 
              reg_frm <=_GEN_412[2:0];
            end 
         if (metaReset)
            begin 
              reg_mcountinhibit <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_mcountinhibit <=3'h0;
               end 
             else 
               begin 
                 reg_mcountinhibit <=_GEN_405[2:0];
               end 
         if (metaReset)
            begin 
              value_lo <=6'h0;
            end 
          else 
            if (reset)
               begin 
                 value_lo <=6'h0;
               end 
             else 
               begin 
                 value_lo <=_GEN_408[5:0];
               end 
         if (metaReset)
            begin 
              value_hi <=58'h0;
            end 
          else 
            if (reset)
               begin 
                 value_hi <=58'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_67)
                       begin 
                         value_hi <=wdata[63:6];
                       end 
                     else 
                       if (_large_T_2)
                          begin 
                            value_hi <=_large_r_T_1;
                          end 
                  end 
                else 
                  if (_large_T_2)
                     begin 
                       value_hi <=_large_r_T_1;
                     end 
         if (metaReset)
            begin 
              value_lo_1 <=6'h0;
            end 
          else 
            if (reset)
               begin 
                 value_lo_1 <=6'h0;
               end 
             else 
               begin 
                 value_lo_1 <=_GEN_406[5:0];
               end 
         if (metaReset)
            begin 
              value_hi_1 <=58'h0;
            end 
          else 
            if (reset)
               begin 
                 value_hi_1 <=58'h0;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_66)
                       begin 
                         value_hi_1 <=wdata[63:6];
                       end 
                     else 
                       if (_large_T_5)
                          begin 
                            value_hi_1 <=_large_r_T_3;
                          end 
                  end 
                else 
                  if (_large_T_5)
                     begin 
                       value_hi_1 <=_large_r_T_3;
                     end 
         if (metaReset)
            begin 
              reg_misa <=64'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_misa <=64'h800000000094112d;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_49)
                       begin 
                         if (_T_1834)
                            begin 
                              reg_misa <=_reg_misa_T_8;
                            end 
                       end 
                  end 
         if (metaReset)
            begin 
              reg_custom_0 <=64'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_custom_0 <=64'h208;
               end 
             else 
               if (csr_wen)
                  begin 
                    if (_T_188)
                       begin 
                         reg_custom_0 <=_reg_custom_0_T_3;
                       end 
                  end 
         if (metaReset)
            begin 
              io_status_dprv_REG <=2'h0;
            end 
          else 
            if (_io_status_dprv_x87_T_1)
               begin 
                 io_status_dprv_REG <=reg_mstatus_mpp;
               end 
             else 
               begin 
                 io_status_dprv_REG <=reg_mstatus_prv;
               end 
         if (metaReset)
            begin 
              io_status_cease_r <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 io_status_cease_r <=1'h0;
               end 
             else 
               begin 
                 io_status_cease_r <=_GEN_181;
               end 
         if (~_T_252)
            begin $display("Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:739 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n");
            end 
         if (~_T_252)
            begin $display("fatal");
            end 
         if (~_T_274)
            begin $display("Assertion failed\n    at CSR.scala:748 assert(!reg_singleStepped || io.retire === UInt(0))\n");
            end 
         if (~_T_274)
            begin $display("fatal");
            end 
         CSRFile_state <=CSRFile_xor0;
         if (!(CSRFile_cov_read_data))
            begin 
              CSRFile_covSum <=CSRFile_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              CSRFile_metaAssert <=1'h0;
            end 
          else 
            begin 
              CSRFile_metaAssert <=CSRFile_metaAssert|CSRFile_or0;
            end 
       end
  
  always @( posedge io_ungated_clock)
       begin 
         if (metaReset)
            begin 
              reg_wfi <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 reg_wfi <=1'h0;
               end 
             else 
               if (_T_260)
                  begin 
                    reg_wfi <=1'h0;
                  end 
                else 
                  begin 
                    reg_wfi <=_GEN_48;
                  end 
       end
  
  always @( posedge clock)
       begin 
         if (CSRFile_cov_write_en&CSRFile_cov_write_mask)
            begin 
              CSRFile_cov [CSRFile_cov_write_addr]<=CSRFile_cov_write_data;
            end 
       end
  
endmodule
 
module BreakpointUnit (
  input io_status_debug,
  input [1:0] io_status_prv,
  input io_bp_0_control_action,
  input [1:0] io_bp_0_control_tmatch,
  input io_bp_0_control_m,
  input io_bp_0_control_s,
  input io_bp_0_control_u,
  input io_bp_0_control_x,
  input io_bp_0_control_w,
  input io_bp_0_control_r,
  input [38:0] io_bp_0_address,
  input [38:0] io_pc,
  input [38:0] io_ea,
  output io_xcpt_if,
  output io_xcpt_ld,
  output io_xcpt_st,
  output io_debug_if,
  output io_debug_ld,
  output io_debug_st,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [3:0] _en_T_1 ;  
   wire [3:0] _en_T_2 ;  
   wire en ;  
   wire _r_T ;  
   wire _r_T_2 ;  
   wire _r_T_4 ;  
   wire r_lo_hi ;  
   wire r_hi_lo ;  
   wire r_hi_hi ;  
   wire [3:0] _r_T_9 ;  
   wire [38:0] _GEN_11 ;  
   wire [38:0] _r_T_10 ;  
   wire [38:0] _r_T_16 ;  
   wire _r_T_17 ;  
   wire _r_T_18 ;  
   wire r ;  
   wire _w_T ;  
   wire w ;  
   wire _x_T ;  
   wire _x_T_2 ;  
   wire _x_T_4 ;  
   wire [38:0] _x_T_10 ;  
   wire _x_T_17 ;  
   wire _x_T_18 ;  
   wire x ;  
   wire [29:0] BreakpointUnit_covSum ;  
  assign _en_T_1={io_bp_0_control_m,1'h0,io_bp_0_control_s,io_bp_0_control_u}; 
  assign _en_T_2=_en_T_1>>io_status_prv; 
  assign en=~io_status_debug&_en_T_2[0]; 
  assign _r_T=en&io_bp_0_control_r; 
  assign _r_T_2=io_ea>=io_bp_0_address; 
  assign _r_T_4=_r_T_2^io_bp_0_control_tmatch[0]; 
  assign r_lo_hi=io_bp_0_control_tmatch[0]&io_bp_0_address[0]; 
  assign r_hi_lo=r_lo_hi&io_bp_0_address[1]; 
  assign r_hi_hi=r_hi_lo&io_bp_0_address[2]; 
  assign _r_T_9={r_hi_hi,r_hi_lo,r_lo_hi,io_bp_0_control_tmatch[0]}; 
  assign _GEN_11={35'b0,_r_T_9}; 
  assign _r_T_10=~io_ea|_GEN_11; 
  assign _r_T_16=~io_bp_0_address|_GEN_11; 
  assign _r_T_17=_r_T_10==_r_T_16; 
  assign _r_T_18=io_bp_0_control_tmatch[1] ? _r_T_4:_r_T_17; 
  assign r=_r_T&_r_T_18; 
  assign _w_T=en&io_bp_0_control_w; 
  assign w=_w_T&_r_T_18; 
  assign _x_T=en&io_bp_0_control_x; 
  assign _x_T_2=io_pc>=io_bp_0_address; 
  assign _x_T_4=_x_T_2^io_bp_0_control_tmatch[0]; 
  assign _x_T_10=~io_pc|_GEN_11; 
  assign _x_T_17=_x_T_10==_r_T_16; 
  assign _x_T_18=io_bp_0_control_tmatch[1] ? _x_T_4:_x_T_17; 
  assign x=_x_T&_x_T_18; 
  assign io_xcpt_if=x&~io_bp_0_control_action; 
  assign io_xcpt_ld=r&~io_bp_0_control_action; 
  assign io_xcpt_st=w&~io_bp_0_control_action; 
  assign io_debug_if=x&io_bp_0_control_action; 
  assign io_debug_ld=r&io_bp_0_control_action; 
  assign io_debug_st=w&io_bp_0_control_action; 
  assign BreakpointUnit_covSum=30'h0; 
  assign io_covSum=BreakpointUnit_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module ALU (
  input io_dw,
  input [3:0] io_fn,
  input [63:0] io_in2,
  input [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output io_cmp_out,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [63:0] in2_inv ;  
   wire [63:0] in1_xor_in2 ;  
   wire [63:0] _io_adder_out_T_1 ;  
   wire [63:0] _GEN_1 ;  
   wire _slt_T_2 ;  
   wire _slt_T_7 ;  
   wire slt ;  
   wire _io_cmp_out_T_3 ;  
   wire _io_cmp_out_T_4 ;  
   wire _T_2 ;  
   wire [31:0] _T_4 ;  
   wire [31:0] hi ;  
   wire hi_1 ;  
   wire [4:0] lo ;  
   wire [5:0] shamt ;  
   wire [31:0] lo_1 ;  
   wire [63:0] shin_r ;  
   wire _shin_T ;  
   wire _shin_T_1 ;  
   wire _shin_T_2 ;  
   wire [63:0] _shin_T_6 ;  
   wire [63:0] _shin_T_8 ;  
   wire [63:0] _shin_T_10 ;  
   wire [63:0] _shin_T_11 ;  
   wire [63:0] _GEN_2 ;  
   wire [63:0] _shin_T_16 ;  
   wire [63:0] _shin_T_18 ;  
   wire [63:0] _shin_T_20 ;  
   wire [63:0] _shin_T_21 ;  
   wire [63:0] _GEN_3 ;  
   wire [63:0] _shin_T_26 ;  
   wire [63:0] _shin_T_28 ;  
   wire [63:0] _shin_T_30 ;  
   wire [63:0] _shin_T_31 ;  
   wire [63:0] _GEN_4 ;  
   wire [63:0] _shin_T_36 ;  
   wire [63:0] _shin_T_38 ;  
   wire [63:0] _shin_T_40 ;  
   wire [63:0] _shin_T_41 ;  
   wire [63:0] _GEN_5 ;  
   wire [63:0] _shin_T_46 ;  
   wire [63:0] _shin_T_48 ;  
   wire [63:0] _shin_T_50 ;  
   wire [63:0] _shin_T_51 ;  
   wire [63:0] _GEN_6 ;  
   wire [63:0] _shin_T_56 ;  
   wire [63:0] _shin_T_58 ;  
   wire [63:0] _shin_T_60 ;  
   wire [63:0] _shin_T_61 ;  
   wire [63:0] shin ;  
   wire shout_r_hi ;  
   wire [64:0] _shout_r_T_3 ;  
   wire [64:0] _shout_r_T_4 ;  
   wire [63:0] shout_r ;  
   wire [63:0] _shout_l_T_3 ;  
   wire [63:0] _shout_l_T_5 ;  
   wire [63:0] _shout_l_T_7 ;  
   wire [63:0] _shout_l_T_8 ;  
   wire [63:0] _GEN_7 ;  
   wire [63:0] _shout_l_T_13 ;  
   wire [63:0] _shout_l_T_15 ;  
   wire [63:0] _shout_l_T_17 ;  
   wire [63:0] _shout_l_T_18 ;  
   wire [63:0] _GEN_8 ;  
   wire [63:0] _shout_l_T_23 ;  
   wire [63:0] _shout_l_T_25 ;  
   wire [63:0] _shout_l_T_27 ;  
   wire [63:0] _shout_l_T_28 ;  
   wire [63:0] _GEN_9 ;  
   wire [63:0] _shout_l_T_33 ;  
   wire [63:0] _shout_l_T_35 ;  
   wire [63:0] _shout_l_T_37 ;  
   wire [63:0] _shout_l_T_38 ;  
   wire [63:0] _GEN_10 ;  
   wire [63:0] _shout_l_T_43 ;  
   wire [63:0] _shout_l_T_45 ;  
   wire [63:0] _shout_l_T_47 ;  
   wire [63:0] _shout_l_T_48 ;  
   wire [63:0] _GEN_11 ;  
   wire [63:0] _shout_l_T_53 ;  
   wire [63:0] _shout_l_T_55 ;  
   wire [63:0] _shout_l_T_57 ;  
   wire [63:0] shout_l ;  
   wire [63:0] _shout_T_3 ;  
   wire _shout_T_4 ;  
   wire [63:0] _shout_T_5 ;  
   wire [63:0] shout ;  
   wire _logic_T ;  
   wire _logic_T_1 ;  
   wire _logic_T_2 ;  
   wire [63:0] _logic_T_3 ;  
   wire _logic_T_5 ;  
   wire _logic_T_6 ;  
   wire [63:0] _logic_T_7 ;  
   wire [63:0] _logic_T_8 ;  
   wire [63:0] logic_ ;  
   wire _shift_logic_T ;  
   wire _shift_logic_T_1 ;  
   wire [63:0] _GEN_12 ;  
   wire [63:0] _shift_logic_T_2 ;  
   wire [63:0] shift_logic ;  
   wire _out_T ;  
   wire _out_T_1 ;  
   wire _out_T_2 ;  
   wire [63:0] out ;  
   wire [31:0] io_out_hi ;  
   wire [31:0] io_out_lo ;  
   wire [63:0] _io_out_T_2 ;  
   wire [29:0] ALU_covSum ;  
  assign in2_inv=io_fn[3] ? ~io_in2:io_in2; 
  assign in1_xor_in2=io_in1^in2_inv; 
  assign _io_adder_out_T_1=io_in1+in2_inv; 
  assign _GEN_1={63'b0,io_fn[3]}; 
  assign _slt_T_2=io_in1[63]==io_in2[63]; 
  assign _slt_T_7=io_fn[1] ? io_in2[63]:io_in1[63]; 
  assign slt=_slt_T_2 ? io_adder_out[63]:_slt_T_7; 
  assign _io_cmp_out_T_3=in1_xor_in2==64'h0; 
  assign _io_cmp_out_T_4=io_fn[3] ? slt:_io_cmp_out_T_3; 
  assign _T_2=io_fn[3]&io_in1[31]; 
  assign _T_4=_T_2 ? 32'hffffffff:32'h0; 
  assign hi=io_dw ? io_in1[63:32]:_T_4; 
  assign hi_1=io_in2[5]&io_dw; 
  assign lo=io_in2[4:0]; 
  assign shamt={hi_1,lo}; 
  assign lo_1=io_in1[31:0]; 
  assign shin_r={hi,lo_1}; 
  assign _shin_T=io_fn==4'h5; 
  assign _shin_T_1=io_fn==4'hb; 
  assign _shin_T_2=_shin_T|_shin_T_1; 
  assign _shin_T_6={32'b0,shin_r[63:32]}; 
  assign _shin_T_8={shin_r[31:0],32'h0}; 
  assign _shin_T_10=_shin_T_8&64'hffffffff00000000; 
  assign _shin_T_11=_shin_T_6|_shin_T_10; 
  assign _GEN_2={16'b0,_shin_T_11[63:16]}; 
  assign _shin_T_16=_GEN_2&64'hffff0000ffff; 
  assign _shin_T_18={_shin_T_11[47:0],16'h0}; 
  assign _shin_T_20=_shin_T_18&64'hffff0000ffff0000; 
  assign _shin_T_21=_shin_T_16|_shin_T_20; 
  assign _GEN_3={8'b0,_shin_T_21[63:8]}; 
  assign _shin_T_26=_GEN_3&64'hff00ff00ff00ff; 
  assign _shin_T_28={_shin_T_21[55:0],8'h0}; 
  assign _shin_T_30=_shin_T_28&64'hff00ff00ff00ff00; 
  assign _shin_T_31=_shin_T_26|_shin_T_30; 
  assign _GEN_4={4'b0,_shin_T_31[63:4]}; 
  assign _shin_T_36=_GEN_4&64'hf0f0f0f0f0f0f0f; 
  assign _shin_T_38={_shin_T_31[59:0],4'h0}; 
  assign _shin_T_40=_shin_T_38&64'hf0f0f0f0f0f0f0f0; 
  assign _shin_T_41=_shin_T_36|_shin_T_40; 
  assign _GEN_5={2'b0,_shin_T_41[63:2]}; 
  assign _shin_T_46=_GEN_5&64'h3333333333333333; 
  assign _shin_T_48={_shin_T_41[61:0],2'h0}; 
  assign _shin_T_50=_shin_T_48&64'hcccccccccccccccc; 
  assign _shin_T_51=_shin_T_46|_shin_T_50; 
  assign _GEN_6={1'b0,_shin_T_51[63:1]}; 
  assign _shin_T_56=_GEN_6&64'h5555555555555555; 
  assign _shin_T_58={_shin_T_51[62:0],1'h0}; 
  assign _shin_T_60=_shin_T_58&64'haaaaaaaaaaaaaaaa; 
  assign _shin_T_61=_shin_T_56|_shin_T_60; 
  assign shin=_shin_T_2 ? shin_r:_shin_T_61; 
  assign shout_r_hi=io_fn[3]&shin[63]; 
  assign _shout_r_T_3={shout_r_hi,shin}; 
  assign _shout_r_T_4=$signed(_shout_r_T_3)>>>shamt; 
  assign shout_r=_shout_r_T_4[63:0]; 
  assign _shout_l_T_3={32'b0,shout_r[63:32]}; 
  assign _shout_l_T_5={shout_r[31:0],32'h0}; 
  assign _shout_l_T_7=_shout_l_T_5&64'hffffffff00000000; 
  assign _shout_l_T_8=_shout_l_T_3|_shout_l_T_7; 
  assign _GEN_7={16'b0,_shout_l_T_8[63:16]}; 
  assign _shout_l_T_13=_GEN_7&64'hffff0000ffff; 
  assign _shout_l_T_15={_shout_l_T_8[47:0],16'h0}; 
  assign _shout_l_T_17=_shout_l_T_15&64'hffff0000ffff0000; 
  assign _shout_l_T_18=_shout_l_T_13|_shout_l_T_17; 
  assign _GEN_8={8'b0,_shout_l_T_18[63:8]}; 
  assign _shout_l_T_23=_GEN_8&64'hff00ff00ff00ff; 
  assign _shout_l_T_25={_shout_l_T_18[55:0],8'h0}; 
  assign _shout_l_T_27=_shout_l_T_25&64'hff00ff00ff00ff00; 
  assign _shout_l_T_28=_shout_l_T_23|_shout_l_T_27; 
  assign _GEN_9={4'b0,_shout_l_T_28[63:4]}; 
  assign _shout_l_T_33=_GEN_9&64'hf0f0f0f0f0f0f0f; 
  assign _shout_l_T_35={_shout_l_T_28[59:0],4'h0}; 
  assign _shout_l_T_37=_shout_l_T_35&64'hf0f0f0f0f0f0f0f0; 
  assign _shout_l_T_38=_shout_l_T_33|_shout_l_T_37; 
  assign _GEN_10={2'b0,_shout_l_T_38[63:2]}; 
  assign _shout_l_T_43=_GEN_10&64'h3333333333333333; 
  assign _shout_l_T_45={_shout_l_T_38[61:0],2'h0}; 
  assign _shout_l_T_47=_shout_l_T_45&64'hcccccccccccccccc; 
  assign _shout_l_T_48=_shout_l_T_43|_shout_l_T_47; 
  assign _GEN_11={1'b0,_shout_l_T_48[63:1]}; 
  assign _shout_l_T_53=_GEN_11&64'h5555555555555555; 
  assign _shout_l_T_55={_shout_l_T_48[62:0],1'h0}; 
  assign _shout_l_T_57=_shout_l_T_55&64'haaaaaaaaaaaaaaaa; 
  assign shout_l=_shout_l_T_53|_shout_l_T_57; 
  assign _shout_T_3=_shin_T_2 ? shout_r:64'h0; 
  assign _shout_T_4=io_fn==4'h1; 
  assign _shout_T_5=_shout_T_4 ? shout_l:64'h0; 
  assign shout=_shout_T_3|_shout_T_5; 
  assign _logic_T=io_fn==4'h4; 
  assign _logic_T_1=io_fn==4'h6; 
  assign _logic_T_2=_logic_T|_logic_T_1; 
  assign _logic_T_3=_logic_T_2 ? in1_xor_in2:64'h0; 
  assign _logic_T_5=io_fn==4'h7; 
  assign _logic_T_6=_logic_T_1|_logic_T_5; 
  assign _logic_T_7=io_in1&io_in2; 
  assign _logic_T_8=_logic_T_6 ? _logic_T_7:64'h0; 
  assign logic_=_logic_T_3|_logic_T_8; 
  assign _shift_logic_T=io_fn>=4'hc; 
  assign _shift_logic_T_1=_shift_logic_T&slt; 
  assign _GEN_12={63'b0,_shift_logic_T_1}; 
  assign _shift_logic_T_2=_GEN_12|logic_; 
  assign shift_logic=_shift_logic_T_2|shout; 
  assign _out_T=io_fn==4'h0; 
  assign _out_T_1=io_fn==4'ha; 
  assign _out_T_2=_out_T|_out_T_1; 
  assign out=_out_T_2 ? io_adder_out:shift_logic; 
  assign io_out_hi=out[31] ? 32'hffffffff:32'h0; 
  assign io_out_lo=out[31:0]; 
  assign _io_out_T_2={io_out_hi,io_out_lo}; 
  assign io_out=io_dw ? out:_io_out_T_2; 
  assign io_adder_out=_io_adder_out_T_1+_GEN_1; 
  assign io_cmp_out=io_fn[0]^_io_cmp_out_T_4; 
  assign ALU_covSum=30'h0; 
  assign io_covSum=ALU_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module MulDiv (
  input clock,
  input reset,
  output io_req_ready,
  input io_req_valid,
  input [3:0] io_req_bits_fn,
  input io_req_bits_dw,
  input [63:0] io_req_bits_in1,
  input [63:0] io_req_bits_in2,
  input [4:0] io_req_bits_tag,
  input io_kill,
  input io_resp_ready,
  output io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0] io_resp_bits_tag,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg [2:0] state ;  
   reg [31:0] _RAND_0 ;  
   reg req_dw ;  
   reg [31:0] _RAND_1 ;  
   reg [4:0] req_tag ;  
   reg [31:0] _RAND_2 ;  
   reg [6:0] count ;  
   reg [31:0] _RAND_3 ;  
   reg neg_out ;  
   reg [31:0] _RAND_4 ;  
   reg isHi ;  
   reg [31:0] _RAND_5 ;  
   reg resHi ;  
   reg [31:0] _RAND_6 ;  
   reg [64:0] divisor ;  
   reg [95:0] _RAND_7 ;  
   reg [129:0] remainder ;  
   reg [159:0] _RAND_8 ;  
   wire [3:0] _T ;  
   wire cmdMul ;  
   wire [3:0] _T_3 ;  
   wire _T_4 ;  
   wire [3:0] _T_5 ;  
   wire _T_6 ;  
   wire cmdHi ;  
   wire [3:0] _T_9 ;  
   wire _T_10 ;  
   wire [3:0] _T_11 ;  
   wire _T_12 ;  
   wire lhsSigned ;  
   wire _T_16 ;  
   wire rhsSigned ;  
   wire _sign_T_2 ;  
   wire lhs_sign ;  
   wire [31:0] _hi_T_1 ;  
   wire [31:0] hi ;  
   wire [31:0] lo ;  
   wire [63:0] lhs_in ;  
   wire _sign_T_5 ;  
   wire rhs_sign ;  
   wire [31:0] _hi_T_4 ;  
   wire [31:0] hi_1 ;  
   wire [31:0] lo_1 ;  
   wire [64:0] subtractor ;  
   wire [63:0] result ;  
   wire [63:0] negated_remainder ;  
   wire _T_23 ;  
   wire _T_26 ;  
   wire _T_27 ;  
   wire [64:0] mulReg_hi ;  
   wire [128:0] mulReg ;  
   wire prod_hi ;  
   wire [63:0] mplier ;  
   wire [64:0] accum ;  
   wire [7:0] prod_lo ;  
   wire [8:0] _prod_T_1 ;  
   wire [64:0] _GEN_37 ;  
   wire [73:0] _prod_T_2 ;  
   wire [73:0] _GEN_38 ;  
   wire [55:0] nextMulReg_lo ;  
   wire [73:0] nextMulReg_hi ;  
   wire [129:0] nextMulReg ;  
   wire _nextMplierSign_T ;  
   wire remainder_hi_lo ;  
   wire [10:0] _eOutMask_T ;  
   wire [64:0] _eOutMask_T_2 ;  
   wire [63:0] eOutMask ;  
   wire _eOut_T ;  
   wire _eOut_T_2 ;  
   wire _eOut_T_3 ;  
   wire _eOut_T_5 ;  
   wire [63:0] _eOut_T_7 ;  
   wire _eOut_T_8 ;  
   wire eOut ;  
   wire [10:0] _eOutRes_T_2 ;  
   wire [128:0] eOutRes ;  
   wire [64:0] nextMulReg1_hi ;  
   wire [129:0] _nextMulReg1_T ;  
   wire [63:0] nextMulReg1_lo ;  
   wire [128:0] nextMulReg1 ;  
   wire [64:0] remainder_hi_hi ;  
   wire [63:0] remainder_lo ;  
   wire [129:0] _remainder_T ;  
   wire [6:0] _count_T_1 ;  
   wire _T_28 ;  
   wire _T_29 ;  
   wire _T_30 ;  
   wire unrolls_less ;  
   wire [63:0] unrolls_hi_hi ;  
   wire unrolls_lo ;  
   wire [128:0] unrolls_0 ;  
   wire _T_31 ;  
   wire _divby0_T ;  
   wire divby0 ;  
   wire [31:0] divisorMSB_hi ;  
   wire [31:0] divisorMSB_lo ;  
   wire divisorMSB_hi_1 ;  
   wire [15:0] divisorMSB_hi_2 ;  
   wire [15:0] divisorMSB_lo_1 ;  
   wire divisorMSB_hi_3 ;  
   wire [7:0] divisorMSB_hi_4 ;  
   wire [7:0] divisorMSB_lo_2 ;  
   wire divisorMSB_hi_5 ;  
   wire [3:0] divisorMSB_hi_6 ;  
   wire [3:0] divisorMSB_lo_3 ;  
   wire divisorMSB_hi_7 ;  
   wire [1:0] _divisorMSB_T_4 ;  
   wire [1:0] _divisorMSB_T_5 ;  
   wire [1:0] _divisorMSB_T_9 ;  
   wire [1:0] _divisorMSB_T_10 ;  
   wire [1:0] divisorMSB_lo_4 ;  
   wire [2:0] _divisorMSB_T_11 ;  
   wire [3:0] divisorMSB_hi_8 ;  
   wire [3:0] divisorMSB_lo_5 ;  
   wire divisorMSB_hi_9 ;  
   wire [1:0] _divisorMSB_T_15 ;  
   wire [1:0] _divisorMSB_T_16 ;  
   wire [1:0] _divisorMSB_T_20 ;  
   wire [1:0] _divisorMSB_T_21 ;  
   wire [1:0] divisorMSB_lo_6 ;  
   wire [2:0] _divisorMSB_T_22 ;  
   wire [2:0] divisorMSB_lo_7 ;  
   wire [3:0] _divisorMSB_T_23 ;  
   wire [7:0] divisorMSB_hi_10 ;  
   wire [7:0] divisorMSB_lo_8 ;  
   wire divisorMSB_hi_11 ;  
   wire [3:0] divisorMSB_hi_12 ;  
   wire [3:0] divisorMSB_lo_9 ;  
   wire divisorMSB_hi_13 ;  
   wire [1:0] _divisorMSB_T_27 ;  
   wire [1:0] _divisorMSB_T_28 ;  
   wire [1:0] _divisorMSB_T_32 ;  
   wire [1:0] _divisorMSB_T_33 ;  
   wire [1:0] divisorMSB_lo_10 ;  
   wire [2:0] _divisorMSB_T_34 ;  
   wire [3:0] divisorMSB_hi_14 ;  
   wire [3:0] divisorMSB_lo_11 ;  
   wire divisorMSB_hi_15 ;  
   wire [1:0] _divisorMSB_T_38 ;  
   wire [1:0] _divisorMSB_T_39 ;  
   wire [1:0] _divisorMSB_T_43 ;  
   wire [1:0] _divisorMSB_T_44 ;  
   wire [1:0] divisorMSB_lo_12 ;  
   wire [2:0] _divisorMSB_T_45 ;  
   wire [2:0] divisorMSB_lo_13 ;  
   wire [3:0] _divisorMSB_T_46 ;  
   wire [3:0] divisorMSB_lo_14 ;  
   wire [4:0] _divisorMSB_T_47 ;  
   wire [15:0] divisorMSB_hi_16 ;  
   wire [15:0] divisorMSB_lo_15 ;  
   wire divisorMSB_hi_17 ;  
   wire [7:0] divisorMSB_hi_18 ;  
   wire [7:0] divisorMSB_lo_16 ;  
   wire divisorMSB_hi_19 ;  
   wire [3:0] divisorMSB_hi_20 ;  
   wire [3:0] divisorMSB_lo_17 ;  
   wire divisorMSB_hi_21 ;  
   wire [1:0] _divisorMSB_T_51 ;  
   wire [1:0] _divisorMSB_T_52 ;  
   wire [1:0] _divisorMSB_T_56 ;  
   wire [1:0] _divisorMSB_T_57 ;  
   wire [1:0] divisorMSB_lo_18 ;  
   wire [2:0] _divisorMSB_T_58 ;  
   wire [3:0] divisorMSB_hi_22 ;  
   wire [3:0] divisorMSB_lo_19 ;  
   wire divisorMSB_hi_23 ;  
   wire [1:0] _divisorMSB_T_62 ;  
   wire [1:0] _divisorMSB_T_63 ;  
   wire [1:0] _divisorMSB_T_67 ;  
   wire [1:0] _divisorMSB_T_68 ;  
   wire [1:0] divisorMSB_lo_20 ;  
   wire [2:0] _divisorMSB_T_69 ;  
   wire [2:0] divisorMSB_lo_21 ;  
   wire [3:0] _divisorMSB_T_70 ;  
   wire [7:0] divisorMSB_hi_24 ;  
   wire [7:0] divisorMSB_lo_22 ;  
   wire divisorMSB_hi_25 ;  
   wire [3:0] divisorMSB_hi_26 ;  
   wire [3:0] divisorMSB_lo_23 ;  
   wire divisorMSB_hi_27 ;  
   wire [1:0] _divisorMSB_T_74 ;  
   wire [1:0] _divisorMSB_T_75 ;  
   wire [1:0] _divisorMSB_T_79 ;  
   wire [1:0] _divisorMSB_T_80 ;  
   wire [1:0] divisorMSB_lo_24 ;  
   wire [2:0] _divisorMSB_T_81 ;  
   wire [3:0] divisorMSB_hi_28 ;  
   wire [3:0] divisorMSB_lo_25 ;  
   wire divisorMSB_hi_29 ;  
   wire [1:0] _divisorMSB_T_85 ;  
   wire [1:0] _divisorMSB_T_86 ;  
   wire [1:0] _divisorMSB_T_90 ;  
   wire [1:0] _divisorMSB_T_91 ;  
   wire [1:0] divisorMSB_lo_26 ;  
   wire [2:0] _divisorMSB_T_92 ;  
   wire [2:0] divisorMSB_lo_27 ;  
   wire [3:0] _divisorMSB_T_93 ;  
   wire [3:0] divisorMSB_lo_28 ;  
   wire [4:0] _divisorMSB_T_94 ;  
   wire [4:0] divisorMSB_lo_29 ;  
   wire [5:0] divisorMSB ;  
   wire [31:0] dividendMSB_hi ;  
   wire [31:0] dividendMSB_lo ;  
   wire dividendMSB_hi_1 ;  
   wire [15:0] dividendMSB_hi_2 ;  
   wire [15:0] dividendMSB_lo_1 ;  
   wire dividendMSB_hi_3 ;  
   wire [7:0] dividendMSB_hi_4 ;  
   wire [7:0] dividendMSB_lo_2 ;  
   wire dividendMSB_hi_5 ;  
   wire [3:0] dividendMSB_hi_6 ;  
   wire [3:0] dividendMSB_lo_3 ;  
   wire dividendMSB_hi_7 ;  
   wire [1:0] _dividendMSB_T_4 ;  
   wire [1:0] _dividendMSB_T_5 ;  
   wire [1:0] _dividendMSB_T_9 ;  
   wire [1:0] _dividendMSB_T_10 ;  
   wire [1:0] dividendMSB_lo_4 ;  
   wire [2:0] _dividendMSB_T_11 ;  
   wire [3:0] dividendMSB_hi_8 ;  
   wire [3:0] dividendMSB_lo_5 ;  
   wire dividendMSB_hi_9 ;  
   wire [1:0] _dividendMSB_T_15 ;  
   wire [1:0] _dividendMSB_T_16 ;  
   wire [1:0] _dividendMSB_T_20 ;  
   wire [1:0] _dividendMSB_T_21 ;  
   wire [1:0] dividendMSB_lo_6 ;  
   wire [2:0] _dividendMSB_T_22 ;  
   wire [2:0] dividendMSB_lo_7 ;  
   wire [3:0] _dividendMSB_T_23 ;  
   wire [7:0] dividendMSB_hi_10 ;  
   wire [7:0] dividendMSB_lo_8 ;  
   wire dividendMSB_hi_11 ;  
   wire [3:0] dividendMSB_hi_12 ;  
   wire [3:0] dividendMSB_lo_9 ;  
   wire dividendMSB_hi_13 ;  
   wire [1:0] _dividendMSB_T_27 ;  
   wire [1:0] _dividendMSB_T_28 ;  
   wire [1:0] _dividendMSB_T_32 ;  
   wire [1:0] _dividendMSB_T_33 ;  
   wire [1:0] dividendMSB_lo_10 ;  
   wire [2:0] _dividendMSB_T_34 ;  
   wire [3:0] dividendMSB_hi_14 ;  
   wire [3:0] dividendMSB_lo_11 ;  
   wire dividendMSB_hi_15 ;  
   wire [1:0] _dividendMSB_T_38 ;  
   wire [1:0] _dividendMSB_T_39 ;  
   wire [1:0] _dividendMSB_T_43 ;  
   wire [1:0] _dividendMSB_T_44 ;  
   wire [1:0] dividendMSB_lo_12 ;  
   wire [2:0] _dividendMSB_T_45 ;  
   wire [2:0] dividendMSB_lo_13 ;  
   wire [3:0] _dividendMSB_T_46 ;  
   wire [3:0] dividendMSB_lo_14 ;  
   wire [4:0] _dividendMSB_T_47 ;  
   wire [15:0] dividendMSB_hi_16 ;  
   wire [15:0] dividendMSB_lo_15 ;  
   wire dividendMSB_hi_17 ;  
   wire [7:0] dividendMSB_hi_18 ;  
   wire [7:0] dividendMSB_lo_16 ;  
   wire dividendMSB_hi_19 ;  
   wire [3:0] dividendMSB_hi_20 ;  
   wire [3:0] dividendMSB_lo_17 ;  
   wire dividendMSB_hi_21 ;  
   wire [1:0] _dividendMSB_T_51 ;  
   wire [1:0] _dividendMSB_T_52 ;  
   wire [1:0] _dividendMSB_T_56 ;  
   wire [1:0] _dividendMSB_T_57 ;  
   wire [1:0] dividendMSB_lo_18 ;  
   wire [2:0] _dividendMSB_T_58 ;  
   wire [3:0] dividendMSB_hi_22 ;  
   wire [3:0] dividendMSB_lo_19 ;  
   wire dividendMSB_hi_23 ;  
   wire [1:0] _dividendMSB_T_62 ;  
   wire [1:0] _dividendMSB_T_63 ;  
   wire [1:0] _dividendMSB_T_67 ;  
   wire [1:0] _dividendMSB_T_68 ;  
   wire [1:0] dividendMSB_lo_20 ;  
   wire [2:0] _dividendMSB_T_69 ;  
   wire [2:0] dividendMSB_lo_21 ;  
   wire [3:0] _dividendMSB_T_70 ;  
   wire [7:0] dividendMSB_hi_24 ;  
   wire [7:0] dividendMSB_lo_22 ;  
   wire dividendMSB_hi_25 ;  
   wire [3:0] dividendMSB_hi_26 ;  
   wire [3:0] dividendMSB_lo_23 ;  
   wire dividendMSB_hi_27 ;  
   wire [1:0] _dividendMSB_T_74 ;  
   wire [1:0] _dividendMSB_T_75 ;  
   wire [1:0] _dividendMSB_T_79 ;  
   wire [1:0] _dividendMSB_T_80 ;  
   wire [1:0] dividendMSB_lo_24 ;  
   wire [2:0] _dividendMSB_T_81 ;  
   wire [3:0] dividendMSB_hi_28 ;  
   wire [3:0] dividendMSB_lo_25 ;  
   wire dividendMSB_hi_29 ;  
   wire [1:0] _dividendMSB_T_85 ;  
   wire [1:0] _dividendMSB_T_86 ;  
   wire [1:0] _dividendMSB_T_90 ;  
   wire [1:0] _dividendMSB_T_91 ;  
   wire [1:0] dividendMSB_lo_26 ;  
   wire [2:0] _dividendMSB_T_92 ;  
   wire [2:0] dividendMSB_lo_27 ;  
   wire [3:0] _dividendMSB_T_93 ;  
   wire [3:0] dividendMSB_lo_28 ;  
   wire [4:0] _dividendMSB_T_94 ;  
   wire [4:0] dividendMSB_lo_29 ;  
   wire [5:0] dividendMSB ;  
   wire [5:0] _eOutPos_T_1 ;  
   wire [5:0] eOutPos ;  
   wire _eOut_T_11 ;  
   wire _eOut_T_12 ;  
   wire eOut_1 ;  
   wire [126:0] _GEN_39 ;  
   wire [126:0] _remainder_T_2 ;  
   wire [128:0] _GEN_16 ;  
   wire _T_33 ;  
   wire _T_34 ;  
   wire _T_35 ;  
   wire _T_36 ;  
   wire _state_T_1 ;  
   wire _count_T_7 ;  
   wire [2:0] _count_T_8 ;  
   wire _neg_out_T ;  
   wire [64:0] _divisor_T ;  
   wire [2:0] _outMul_T_1 ;  
   wire outMul ;  
   wire _loOut_T_3 ;  
   wire [31:0] loOut ;  
   wire [31:0] _hiOut_T_4 ;  
   wire [31:0] hiOut ;  
   wire _io_resp_valid_T ;  
   wire _io_resp_valid_T_1 ;  
   reg [19:0] MulDiv_state ;  
   reg [31:0] _RAND_9 ;  
   reg MulDiv_cov[0:1048575] ;  
   reg [31:0] _RAND_10 ;  
   wire MulDiv_cov_read_data ;  
   wire [19:0] MulDiv_cov_read_addr ;  
   wire MulDiv_cov_write_data ;  
   wire [19:0] MulDiv_cov_write_addr ;  
   wire MulDiv_cov_write_mask ;  
   wire MulDiv_cov_write_en ;  
   reg [29:0] MulDiv_covSum ;  
   reg [31:0] _RAND_11 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire mux_cond_4 ;  
   wire mux_cond_5 ;  
   wire mux_cond_6 ;  
   wire mux_cond_7 ;  
   wire mux_cond_8 ;  
   wire mux_cond_9 ;  
   wire mux_cond_10 ;  
   wire mux_cond_11 ;  
   wire mux_cond_12 ;  
   wire mux_cond_13 ;  
   wire mux_cond_14 ;  
   wire mux_cond_15 ;  
   wire mux_cond_16 ;  
   wire mux_cond_17 ;  
   wire mux_cond_18 ;  
   wire mux_cond_19 ;  
   wire mux_cond_20 ;  
   wire mux_cond_21 ;  
   wire mux_cond_22 ;  
   wire mux_cond_23 ;  
   wire mux_cond_24 ;  
   wire mux_cond_25 ;  
   wire mux_cond_26 ;  
   wire mux_cond_27 ;  
   wire mux_cond_28 ;  
   wire mux_cond_29 ;  
   wire mux_cond_30 ;  
   wire mux_cond_31 ;  
   wire mux_cond_32 ;  
   wire mux_cond_33 ;  
   wire mux_cond_34 ;  
   wire mux_cond_35 ;  
   wire mux_cond_36 ;  
   wire mux_cond_37 ;  
   wire mux_cond_38 ;  
   wire mux_cond_39 ;  
   wire mux_cond_40 ;  
   wire mux_cond_41 ;  
   wire mux_cond_42 ;  
   wire mux_cond_43 ;  
   wire mux_cond_44 ;  
   wire mux_cond_45 ;  
   wire mux_cond_46 ;  
   wire mux_cond_47 ;  
   wire mux_cond_48 ;  
   wire mux_cond_49 ;  
   wire mux_cond_50 ;  
   wire mux_cond_51 ;  
   wire mux_cond_52 ;  
   wire mux_cond_53 ;  
   wire mux_cond_54 ;  
   wire mux_cond_55 ;  
   wire mux_cond_56 ;  
   wire mux_cond_57 ;  
   wire mux_cond_58 ;  
   wire mux_cond_59 ;  
   wire mux_cond_60 ;  
   wire mux_cond_61 ;  
   wire mux_cond_62 ;  
   wire mux_cond_63 ;  
   wire mux_cond_64 ;  
   wire mux_cond_65 ;  
   wire mux_cond_66 ;  
   wire mux_cond_67 ;  
   wire mux_cond_68 ;  
   wire mux_cond_69 ;  
   wire mux_cond_70 ;  
   wire mux_cond_71 ;  
   wire mux_cond_72 ;  
   wire mux_cond_73 ;  
   wire mux_cond_74 ;  
   wire mux_cond_75 ;  
   wire mux_cond_76 ;  
   wire mux_cond_77 ;  
   wire mux_cond_78 ;  
   wire mux_cond_79 ;  
   wire mux_cond_80 ;  
   wire mux_cond_81 ;  
   wire mux_cond_82 ;  
   wire mux_cond_83 ;  
   wire mux_cond_84 ;  
   wire mux_cond_85 ;  
   wire mux_cond_86 ;  
   wire mux_cond_87 ;  
   wire mux_cond_88 ;  
   wire mux_cond_89 ;  
   wire mux_cond_90 ;  
   wire mux_cond_91 ;  
   wire mux_cond_92 ;  
   wire mux_cond_93 ;  
   wire mux_cond_94 ;  
   wire mux_cond_95 ;  
   wire mux_cond_96 ;  
   wire mux_cond_97 ;  
   wire [4:0] isHi_shl ;  
   wire [19:0] isHi_pad ;  
   wire [12:0] neg_out_shl ;  
   wire [19:0] neg_out_pad ;  
   wire [4:0] req_dw_shl ;  
   wire [19:0] req_dw_pad ;  
   wire [10:0] state_shl ;  
   wire [19:0] state_pad ;  
   wire [1:0] resHi_shl ;  
   wire [19:0] resHi_pad ;  
   wire [12:0] mux_cond_0_shl ;  
   wire [19:0] mux_cond_0_pad ;  
   wire [1:0] mux_cond_1_shl ;  
   wire [19:0] mux_cond_1_pad ;  
   wire mux_cond_2_shl ;  
   wire [19:0] mux_cond_2_pad ;  
   wire [12:0] mux_cond_3_shl ;  
   wire [19:0] mux_cond_3_pad ;  
   wire [15:0] mux_cond_4_shl ;  
   wire [19:0] mux_cond_4_pad ;  
   wire [11:0] mux_cond_5_shl ;  
   wire [19:0] mux_cond_5_pad ;  
   wire [7:0] mux_cond_6_shl ;  
   wire [19:0] mux_cond_6_pad ;  
   wire [17:0] mux_cond_7_shl ;  
   wire [19:0] mux_cond_7_pad ;  
   wire [11:0] mux_cond_8_shl ;  
   wire [19:0] mux_cond_8_pad ;  
   wire [15:0] mux_cond_9_shl ;  
   wire [19:0] mux_cond_9_pad ;  
   wire [13:0] mux_cond_10_shl ;  
   wire [19:0] mux_cond_10_pad ;  
   wire mux_cond_11_shl ;  
   wire [19:0] mux_cond_11_pad ;  
   wire [7:0] mux_cond_12_shl ;  
   wire [19:0] mux_cond_12_pad ;  
   wire [13:0] mux_cond_13_shl ;  
   wire [19:0] mux_cond_13_pad ;  
   wire mux_cond_14_shl ;  
   wire [19:0] mux_cond_14_pad ;  
   wire [9:0] mux_cond_15_shl ;  
   wire [19:0] mux_cond_15_pad ;  
   wire [8:0] mux_cond_16_shl ;  
   wire [19:0] mux_cond_16_pad ;  
   wire [8:0] mux_cond_17_shl ;  
   wire [19:0] mux_cond_17_pad ;  
   wire [8:0] mux_cond_18_shl ;  
   wire [19:0] mux_cond_18_pad ;  
   wire [2:0] mux_cond_19_shl ;  
   wire [19:0] mux_cond_19_pad ;  
   wire [16:0] mux_cond_20_shl ;  
   wire [19:0] mux_cond_20_pad ;  
   wire [6:0] mux_cond_21_shl ;  
   wire [19:0] mux_cond_21_pad ;  
   wire [11:0] mux_cond_22_shl ;  
   wire [19:0] mux_cond_22_pad ;  
   wire mux_cond_23_shl ;  
   wire [19:0] mux_cond_23_pad ;  
   wire [6:0] mux_cond_24_shl ;  
   wire [19:0] mux_cond_24_pad ;  
   wire [12:0] mux_cond_25_shl ;  
   wire [19:0] mux_cond_25_pad ;  
   wire [4:0] mux_cond_26_shl ;  
   wire [19:0] mux_cond_26_pad ;  
   wire [11:0] mux_cond_27_shl ;  
   wire [19:0] mux_cond_27_pad ;  
   wire [6:0] mux_cond_28_shl ;  
   wire [19:0] mux_cond_28_pad ;  
   wire [12:0] mux_cond_29_shl ;  
   wire [19:0] mux_cond_29_pad ;  
   wire [1:0] mux_cond_30_shl ;  
   wire [19:0] mux_cond_30_pad ;  
   wire [11:0] mux_cond_31_shl ;  
   wire [19:0] mux_cond_31_pad ;  
   wire [6:0] mux_cond_32_shl ;  
   wire [19:0] mux_cond_32_pad ;  
   wire [5:0] mux_cond_33_shl ;  
   wire [19:0] mux_cond_33_pad ;  
   wire [18:0] mux_cond_34_shl ;  
   wire [19:0] mux_cond_34_pad ;  
   wire [12:0] mux_cond_35_shl ;  
   wire [19:0] mux_cond_35_pad ;  
   wire mux_cond_36_shl ;  
   wire [19:0] mux_cond_36_pad ;  
   wire [8:0] mux_cond_37_shl ;  
   wire [19:0] mux_cond_37_pad ;  
   wire [5:0] mux_cond_38_shl ;  
   wire [19:0] mux_cond_38_pad ;  
   wire [16:0] mux_cond_39_shl ;  
   wire [19:0] mux_cond_39_pad ;  
   wire [3:0] mux_cond_40_shl ;  
   wire [19:0] mux_cond_40_pad ;  
   wire [9:0] mux_cond_41_shl ;  
   wire [19:0] mux_cond_41_pad ;  
   wire [15:0] mux_cond_42_shl ;  
   wire [19:0] mux_cond_42_pad ;  
   wire [13:0] mux_cond_43_shl ;  
   wire [19:0] mux_cond_43_pad ;  
   wire [12:0] mux_cond_44_shl ;  
   wire [19:0] mux_cond_44_pad ;  
   wire mux_cond_45_shl ;  
   wire [19:0] mux_cond_45_pad ;  
   wire [3:0] mux_cond_46_shl ;  
   wire [19:0] mux_cond_46_pad ;  
   wire [14:0] mux_cond_47_shl ;  
   wire [19:0] mux_cond_47_pad ;  
   wire [16:0] mux_cond_48_shl ;  
   wire [19:0] mux_cond_48_pad ;  
   wire [18:0] mux_cond_49_shl ;  
   wire [19:0] mux_cond_49_pad ;  
   wire mux_cond_50_shl ;  
   wire [19:0] mux_cond_50_pad ;  
   wire [7:0] mux_cond_51_shl ;  
   wire [19:0] mux_cond_51_pad ;  
   wire mux_cond_52_shl ;  
   wire [19:0] mux_cond_52_pad ;  
   wire [19:0] mux_cond_53_shl ;  
   wire [19:0] mux_cond_53_pad ;  
   wire [10:0] mux_cond_54_shl ;  
   wire [19:0] mux_cond_54_pad ;  
   wire [13:0] mux_cond_55_shl ;  
   wire [19:0] mux_cond_55_pad ;  
   wire [9:0] mux_cond_56_shl ;  
   wire [19:0] mux_cond_56_pad ;  
   wire [6:0] mux_cond_57_shl ;  
   wire [19:0] mux_cond_57_pad ;  
   wire [17:0] mux_cond_58_shl ;  
   wire [19:0] mux_cond_58_pad ;  
   wire [19:0] mux_cond_59_shl ;  
   wire [19:0] mux_cond_59_pad ;  
   wire [3:0] mux_cond_60_shl ;  
   wire [19:0] mux_cond_60_pad ;  
   wire [14:0] mux_cond_61_shl ;  
   wire [19:0] mux_cond_61_pad ;  
   wire [4:0] mux_cond_62_shl ;  
   wire [19:0] mux_cond_62_pad ;  
   wire mux_cond_63_shl ;  
   wire [19:0] mux_cond_63_pad ;  
   wire [10:0] mux_cond_64_shl ;  
   wire [19:0] mux_cond_64_pad ;  
   wire [17:0] mux_cond_65_shl ;  
   wire [19:0] mux_cond_65_pad ;  
   wire [9:0] mux_cond_66_shl ;  
   wire [19:0] mux_cond_66_pad ;  
   wire [6:0] mux_cond_67_shl ;  
   wire [19:0] mux_cond_67_pad ;  
   wire [19:0] mux_cond_68_shl ;  
   wire [19:0] mux_cond_68_pad ;  
   wire [10:0] mux_cond_69_shl ;  
   wire [19:0] mux_cond_69_pad ;  
   wire [10:0] mux_cond_70_shl ;  
   wire [19:0] mux_cond_70_pad ;  
   wire [13:0] mux_cond_71_shl ;  
   wire [19:0] mux_cond_71_pad ;  
   wire [18:0] mux_cond_72_shl ;  
   wire [19:0] mux_cond_72_pad ;  
   wire [12:0] mux_cond_73_shl ;  
   wire [19:0] mux_cond_73_pad ;  
   wire [13:0] mux_cond_74_shl ;  
   wire [19:0] mux_cond_74_pad ;  
   wire [13:0] mux_cond_75_shl ;  
   wire [19:0] mux_cond_75_pad ;  
   wire [13:0] mux_cond_76_shl ;  
   wire [19:0] mux_cond_76_pad ;  
   wire [13:0] mux_cond_77_shl ;  
   wire [19:0] mux_cond_77_pad ;  
   wire [17:0] mux_cond_78_shl ;  
   wire [19:0] mux_cond_78_pad ;  
   wire [12:0] mux_cond_79_shl ;  
   wire [19:0] mux_cond_79_pad ;  
   wire [17:0] mux_cond_80_shl ;  
   wire [19:0] mux_cond_80_pad ;  
   wire [13:0] mux_cond_81_shl ;  
   wire [19:0] mux_cond_81_pad ;  
   wire [12:0] mux_cond_82_shl ;  
   wire [19:0] mux_cond_82_pad ;  
   wire [4:0] mux_cond_83_shl ;  
   wire [19:0] mux_cond_83_pad ;  
   wire [16:0] mux_cond_84_shl ;  
   wire [19:0] mux_cond_84_pad ;  
   wire [9:0] mux_cond_85_shl ;  
   wire [19:0] mux_cond_85_pad ;  
   wire [10:0] mux_cond_86_shl ;  
   wire [19:0] mux_cond_86_pad ;  
   wire [2:0] mux_cond_87_shl ;  
   wire [19:0] mux_cond_87_pad ;  
   wire [6:0] mux_cond_88_shl ;  
   wire [19:0] mux_cond_88_pad ;  
   wire [11:0] mux_cond_89_shl ;  
   wire [19:0] mux_cond_89_pad ;  
   wire [7:0] mux_cond_90_shl ;  
   wire [19:0] mux_cond_90_pad ;  
   wire [16:0] mux_cond_91_shl ;  
   wire [19:0] mux_cond_91_pad ;  
   wire [17:0] mux_cond_92_shl ;  
   wire [19:0] mux_cond_92_pad ;  
   wire [5:0] mux_cond_93_shl ;  
   wire [19:0] mux_cond_93_pad ;  
   wire [18:0] mux_cond_94_shl ;  
   wire [19:0] mux_cond_94_pad ;  
   wire [1:0] mux_cond_95_shl ;  
   wire [19:0] mux_cond_95_pad ;  
   wire [17:0] mux_cond_96_shl ;  
   wire [19:0] mux_cond_96_pad ;  
   wire [1:0] mux_cond_97_shl ;  
   wire [19:0] mux_cond_97_pad ;  
   wire [19:0] MulDiv_xor64 ;  
   wire [19:0] MulDiv_xor31 ;  
   wire [19:0] MulDiv_xor66 ;  
   wire [19:0] MulDiv_xor32 ;  
   wire [19:0] MulDiv_xor15 ;  
   wire [19:0] MulDiv_xor68 ;  
   wire [19:0] MulDiv_xor33 ;  
   wire [19:0] MulDiv_xor70 ;  
   wire [19:0] MulDiv_xor34 ;  
   wire [19:0] MulDiv_xor16 ;  
   wire [19:0] MulDiv_xor7 ;  
   wire [19:0] MulDiv_xor72 ;  
   wire [19:0] MulDiv_xor35 ;  
   wire [19:0] MulDiv_xor74 ;  
   wire [19:0] MulDiv_xor36 ;  
   wire [19:0] MulDiv_xor17 ;  
   wire [19:0] MulDiv_xor76 ;  
   wire [19:0] MulDiv_xor37 ;  
   wire [19:0] MulDiv_xor77 ;  
   wire [19:0] MulDiv_xor78 ;  
   wire [19:0] MulDiv_xor38 ;  
   wire [19:0] MulDiv_xor18 ;  
   wire [19:0] MulDiv_xor8 ;  
   wire [19:0] MulDiv_xor3 ;  
   wire [19:0] MulDiv_xor80 ;  
   wire [19:0] MulDiv_xor39 ;  
   wire [19:0] MulDiv_xor82 ;  
   wire [19:0] MulDiv_xor40 ;  
   wire [19:0] MulDiv_xor19 ;  
   wire [19:0] MulDiv_xor84 ;  
   wire [19:0] MulDiv_xor41 ;  
   wire [19:0] MulDiv_xor85 ;  
   wire [19:0] MulDiv_xor86 ;  
   wire [19:0] MulDiv_xor42 ;  
   wire [19:0] MulDiv_xor20 ;  
   wire [19:0] MulDiv_xor9 ;  
   wire [19:0] MulDiv_xor88 ;  
   wire [19:0] MulDiv_xor43 ;  
   wire [19:0] MulDiv_xor90 ;  
   wire [19:0] MulDiv_xor44 ;  
   wire [19:0] MulDiv_xor21 ;  
   wire [19:0] MulDiv_xor92 ;  
   wire [19:0] MulDiv_xor45 ;  
   wire [19:0] MulDiv_xor93 ;  
   wire [19:0] MulDiv_xor94 ;  
   wire [19:0] MulDiv_xor46 ;  
   wire [19:0] MulDiv_xor22 ;  
   wire [19:0] MulDiv_xor10 ;  
   wire [19:0] MulDiv_xor4 ;  
   wire [19:0] MulDiv_xor1 ;  
   wire [19:0] MulDiv_xor96 ;  
   wire [19:0] MulDiv_xor47 ;  
   wire [19:0] MulDiv_xor98 ;  
   wire [19:0] MulDiv_xor48 ;  
   wire [19:0] MulDiv_xor23 ;  
   wire [19:0] MulDiv_xor100 ;  
   wire [19:0] MulDiv_xor49 ;  
   wire [19:0] MulDiv_xor101 ;  
   wire [19:0] MulDiv_xor102 ;  
   wire [19:0] MulDiv_xor50 ;  
   wire [19:0] MulDiv_xor24 ;  
   wire [19:0] MulDiv_xor11 ;  
   wire [19:0] MulDiv_xor104 ;  
   wire [19:0] MulDiv_xor51 ;  
   wire [19:0] MulDiv_xor106 ;  
   wire [19:0] MulDiv_xor52 ;  
   wire [19:0] MulDiv_xor25 ;  
   wire [19:0] MulDiv_xor108 ;  
   wire [19:0] MulDiv_xor53 ;  
   wire [19:0] MulDiv_xor109 ;  
   wire [19:0] MulDiv_xor110 ;  
   wire [19:0] MulDiv_xor54 ;  
   wire [19:0] MulDiv_xor26 ;  
   wire [19:0] MulDiv_xor12 ;  
   wire [19:0] MulDiv_xor5 ;  
   wire [19:0] MulDiv_xor112 ;  
   wire [19:0] MulDiv_xor55 ;  
   wire [19:0] MulDiv_xor114 ;  
   wire [19:0] MulDiv_xor56 ;  
   wire [19:0] MulDiv_xor27 ;  
   wire [19:0] MulDiv_xor116 ;  
   wire [19:0] MulDiv_xor57 ;  
   wire [19:0] MulDiv_xor117 ;  
   wire [19:0] MulDiv_xor118 ;  
   wire [19:0] MulDiv_xor58 ;  
   wire [19:0] MulDiv_xor28 ;  
   wire [19:0] MulDiv_xor13 ;  
   wire [19:0] MulDiv_xor120 ;  
   wire [19:0] MulDiv_xor59 ;  
   wire [19:0] MulDiv_xor122 ;  
   wire [19:0] MulDiv_xor60 ;  
   wire [19:0] MulDiv_xor29 ;  
   wire [19:0] MulDiv_xor124 ;  
   wire [19:0] MulDiv_xor61 ;  
   wire [19:0] MulDiv_xor125 ;  
   wire [19:0] MulDiv_xor126 ;  
   wire [19:0] MulDiv_xor62 ;  
   wire [19:0] MulDiv_xor30 ;  
   wire [19:0] MulDiv_xor14 ;  
   wire [19:0] MulDiv_xor6 ;  
   wire [19:0] MulDiv_xor2 ;  
   wire [19:0] MulDiv_xor0 ;  
  assign _T=io_req_bits_fn&4'h4; 
  assign cmdMul=_T==4'h0; 
  assign _T_3=io_req_bits_fn&4'h5; 
  assign _T_4=_T_3==4'h1; 
  assign _T_5=io_req_bits_fn&4'h2; 
  assign _T_6=_T_5==4'h2; 
  assign cmdHi=_T_4|_T_6; 
  assign _T_9=io_req_bits_fn&4'h6; 
  assign _T_10=_T_9==4'h0; 
  assign _T_11=io_req_bits_fn&4'h1; 
  assign _T_12=_T_11==4'h0; 
  assign lhsSigned=_T_10|_T_12; 
  assign _T_16=_T_3==4'h4; 
  assign rhsSigned=_T_10|_T_16; 
  assign _sign_T_2=io_req_bits_dw ? io_req_bits_in1[63]:io_req_bits_in1[31]; 
  assign lhs_sign=lhsSigned&_sign_T_2; 
  assign _hi_T_1=lhs_sign ? 32'hffffffff:32'h0; 
  assign hi=io_req_bits_dw ? io_req_bits_in1[63:32]:_hi_T_1; 
  assign lo=io_req_bits_in1[31:0]; 
  assign lhs_in={hi,lo}; 
  assign _sign_T_5=io_req_bits_dw ? io_req_bits_in2[63]:io_req_bits_in2[31]; 
  assign rhs_sign=rhsSigned&_sign_T_5; 
  assign _hi_T_4=rhs_sign ? 32'hffffffff:32'h0; 
  assign hi_1=io_req_bits_dw ? io_req_bits_in2[63:32]:_hi_T_4; 
  assign lo_1=io_req_bits_in2[31:0]; 
  assign subtractor=remainder[128:64]-divisor; 
  assign result=resHi ? remainder[128:65]:remainder[63:0]; 
  assign negated_remainder=64'h0-result; 
  assign _T_23=state==3'h1; 
  assign _T_26=state==3'h5; 
  assign _T_27=state==3'h2; 
  assign mulReg_hi=remainder[129:65]; 
  assign mulReg={mulReg_hi,remainder[63:0]}; 
  assign prod_hi=remainder[64]; 
  assign mplier=mulReg[63:0]; 
  assign accum=mulReg[128:64]; 
  assign prod_lo=mplier[7:0]; 
  assign _prod_T_1={prod_hi,prod_lo}; 
  assign _GEN_37={{56{_prod_T_1[8]}},_prod_T_1}; 
  assign _prod_T_2=$signed(_GEN_37)*$signed(divisor); 
  assign _GEN_38={{9{accum[64]}},accum}; 
  assign nextMulReg_lo=mplier[63:8]; 
  assign nextMulReg_hi=$signed(_prod_T_2)+$signed(_GEN_38); 
  assign nextMulReg={nextMulReg_hi,nextMulReg_lo}; 
  assign _nextMplierSign_T=count==7'h6; 
  assign remainder_hi_lo=_nextMplierSign_T&neg_out; 
  assign _eOutMask_T=count*7'h8; 
  assign _eOutMask_T_2=-65'sh10000000000000000>>>_eOutMask_T[5:0]; 
  assign eOutMask=_eOutMask_T_2[63:0]; 
  assign _eOut_T=count!=7'h7; 
  assign _eOut_T_2=count!=7'h0; 
  assign _eOut_T_3=_eOut_T&_eOut_T_2; 
  assign _eOut_T_5=_eOut_T_3&~isHi; 
  assign _eOut_T_7=mplier&~eOutMask; 
  assign _eOut_T_8=_eOut_T_7==64'h0; 
  assign eOut=_eOut_T_5&_eOut_T_8; 
  assign _eOutRes_T_2=11'h40-_eOutMask_T; 
  assign eOutRes=mulReg>>_eOutRes_T_2[5:0]; 
  assign nextMulReg1_hi=nextMulReg[128:64]; 
  assign _nextMulReg1_T=eOut ? {1'b0,eOutRes}:nextMulReg; 
  assign nextMulReg1_lo=_nextMulReg1_T[63:0]; 
  assign nextMulReg1={nextMulReg1_hi,nextMulReg1_lo}; 
  assign remainder_hi_hi=nextMulReg1[128:64]; 
  assign remainder_lo=nextMulReg1[63:0]; 
  assign _remainder_T={remainder_hi_hi,remainder_hi_lo,remainder_lo}; 
  assign _count_T_1=count+7'h1; 
  assign _T_28=count==7'h7; 
  assign _T_29=eOut|_T_28; 
  assign _T_30=state==3'h3; 
  assign unrolls_less=subtractor[64]; 
  assign unrolls_hi_hi=unrolls_less ? remainder[127:64]:subtractor[63:0]; 
  assign unrolls_lo=~unrolls_less; 
  assign unrolls_0={unrolls_hi_hi,remainder[63:0],unrolls_lo}; 
  assign _T_31=count==7'h40; 
  assign _divby0_T=count==7'h0; 
  assign divby0=_divby0_T&unrolls_lo; 
  assign divisorMSB_hi=divisor[63:32]; 
  assign divisorMSB_lo=divisor[31:0]; 
  assign divisorMSB_hi_1=|divisorMSB_hi; 
  assign divisorMSB_hi_2=divisorMSB_hi[31:16]; 
  assign divisorMSB_lo_1=divisorMSB_hi[15:0]; 
  assign divisorMSB_hi_3=|divisorMSB_hi_2; 
  assign divisorMSB_hi_4=divisorMSB_hi_2[15:8]; 
  assign divisorMSB_lo_2=divisorMSB_hi_2[7:0]; 
  assign divisorMSB_hi_5=|divisorMSB_hi_4; 
  assign divisorMSB_hi_6=divisorMSB_hi_4[7:4]; 
  assign divisorMSB_lo_3=divisorMSB_hi_4[3:0]; 
  assign divisorMSB_hi_7=|divisorMSB_hi_6; 
  assign _divisorMSB_T_4=divisorMSB_hi_6[2] ? 2'h2:{1'b0,divisorMSB_hi_6[1]}; 
  assign _divisorMSB_T_5=divisorMSB_hi_6[3] ? 2'h3:_divisorMSB_T_4; 
  assign _divisorMSB_T_9=divisorMSB_lo_3[2] ? 2'h2:{1'b0,divisorMSB_lo_3[1]}; 
  assign _divisorMSB_T_10=divisorMSB_lo_3[3] ? 2'h3:_divisorMSB_T_9; 
  assign divisorMSB_lo_4=divisorMSB_hi_7 ? _divisorMSB_T_5:_divisorMSB_T_10; 
  assign _divisorMSB_T_11={divisorMSB_hi_7,divisorMSB_lo_4}; 
  assign divisorMSB_hi_8=divisorMSB_lo_2[7:4]; 
  assign divisorMSB_lo_5=divisorMSB_lo_2[3:0]; 
  assign divisorMSB_hi_9=|divisorMSB_hi_8; 
  assign _divisorMSB_T_15=divisorMSB_hi_8[2] ? 2'h2:{1'b0,divisorMSB_hi_8[1]}; 
  assign _divisorMSB_T_16=divisorMSB_hi_8[3] ? 2'h3:_divisorMSB_T_15; 
  assign _divisorMSB_T_20=divisorMSB_lo_5[2] ? 2'h2:{1'b0,divisorMSB_lo_5[1]}; 
  assign _divisorMSB_T_21=divisorMSB_lo_5[3] ? 2'h3:_divisorMSB_T_20; 
  assign divisorMSB_lo_6=divisorMSB_hi_9 ? _divisorMSB_T_16:_divisorMSB_T_21; 
  assign _divisorMSB_T_22={divisorMSB_hi_9,divisorMSB_lo_6}; 
  assign divisorMSB_lo_7=divisorMSB_hi_5 ? _divisorMSB_T_11:_divisorMSB_T_22; 
  assign _divisorMSB_T_23={divisorMSB_hi_5,divisorMSB_lo_7}; 
  assign divisorMSB_hi_10=divisorMSB_lo_1[15:8]; 
  assign divisorMSB_lo_8=divisorMSB_lo_1[7:0]; 
  assign divisorMSB_hi_11=|divisorMSB_hi_10; 
  assign divisorMSB_hi_12=divisorMSB_hi_10[7:4]; 
  assign divisorMSB_lo_9=divisorMSB_hi_10[3:0]; 
  assign divisorMSB_hi_13=|divisorMSB_hi_12; 
  assign _divisorMSB_T_27=divisorMSB_hi_12[2] ? 2'h2:{1'b0,divisorMSB_hi_12[1]}; 
  assign _divisorMSB_T_28=divisorMSB_hi_12[3] ? 2'h3:_divisorMSB_T_27; 
  assign _divisorMSB_T_32=divisorMSB_lo_9[2] ? 2'h2:{1'b0,divisorMSB_lo_9[1]}; 
  assign _divisorMSB_T_33=divisorMSB_lo_9[3] ? 2'h3:_divisorMSB_T_32; 
  assign divisorMSB_lo_10=divisorMSB_hi_13 ? _divisorMSB_T_28:_divisorMSB_T_33; 
  assign _divisorMSB_T_34={divisorMSB_hi_13,divisorMSB_lo_10}; 
  assign divisorMSB_hi_14=divisorMSB_lo_8[7:4]; 
  assign divisorMSB_lo_11=divisorMSB_lo_8[3:0]; 
  assign divisorMSB_hi_15=|divisorMSB_hi_14; 
  assign _divisorMSB_T_38=divisorMSB_hi_14[2] ? 2'h2:{1'b0,divisorMSB_hi_14[1]}; 
  assign _divisorMSB_T_39=divisorMSB_hi_14[3] ? 2'h3:_divisorMSB_T_38; 
  assign _divisorMSB_T_43=divisorMSB_lo_11[2] ? 2'h2:{1'b0,divisorMSB_lo_11[1]}; 
  assign _divisorMSB_T_44=divisorMSB_lo_11[3] ? 2'h3:_divisorMSB_T_43; 
  assign divisorMSB_lo_12=divisorMSB_hi_15 ? _divisorMSB_T_39:_divisorMSB_T_44; 
  assign _divisorMSB_T_45={divisorMSB_hi_15,divisorMSB_lo_12}; 
  assign divisorMSB_lo_13=divisorMSB_hi_11 ? _divisorMSB_T_34:_divisorMSB_T_45; 
  assign _divisorMSB_T_46={divisorMSB_hi_11,divisorMSB_lo_13}; 
  assign divisorMSB_lo_14=divisorMSB_hi_3 ? _divisorMSB_T_23:_divisorMSB_T_46; 
  assign _divisorMSB_T_47={divisorMSB_hi_3,divisorMSB_lo_14}; 
  assign divisorMSB_hi_16=divisorMSB_lo[31:16]; 
  assign divisorMSB_lo_15=divisorMSB_lo[15:0]; 
  assign divisorMSB_hi_17=|divisorMSB_hi_16; 
  assign divisorMSB_hi_18=divisorMSB_hi_16[15:8]; 
  assign divisorMSB_lo_16=divisorMSB_hi_16[7:0]; 
  assign divisorMSB_hi_19=|divisorMSB_hi_18; 
  assign divisorMSB_hi_20=divisorMSB_hi_18[7:4]; 
  assign divisorMSB_lo_17=divisorMSB_hi_18[3:0]; 
  assign divisorMSB_hi_21=|divisorMSB_hi_20; 
  assign _divisorMSB_T_51=divisorMSB_hi_20[2] ? 2'h2:{1'b0,divisorMSB_hi_20[1]}; 
  assign _divisorMSB_T_52=divisorMSB_hi_20[3] ? 2'h3:_divisorMSB_T_51; 
  assign _divisorMSB_T_56=divisorMSB_lo_17[2] ? 2'h2:{1'b0,divisorMSB_lo_17[1]}; 
  assign _divisorMSB_T_57=divisorMSB_lo_17[3] ? 2'h3:_divisorMSB_T_56; 
  assign divisorMSB_lo_18=divisorMSB_hi_21 ? _divisorMSB_T_52:_divisorMSB_T_57; 
  assign _divisorMSB_T_58={divisorMSB_hi_21,divisorMSB_lo_18}; 
  assign divisorMSB_hi_22=divisorMSB_lo_16[7:4]; 
  assign divisorMSB_lo_19=divisorMSB_lo_16[3:0]; 
  assign divisorMSB_hi_23=|divisorMSB_hi_22; 
  assign _divisorMSB_T_62=divisorMSB_hi_22[2] ? 2'h2:{1'b0,divisorMSB_hi_22[1]}; 
  assign _divisorMSB_T_63=divisorMSB_hi_22[3] ? 2'h3:_divisorMSB_T_62; 
  assign _divisorMSB_T_67=divisorMSB_lo_19[2] ? 2'h2:{1'b0,divisorMSB_lo_19[1]}; 
  assign _divisorMSB_T_68=divisorMSB_lo_19[3] ? 2'h3:_divisorMSB_T_67; 
  assign divisorMSB_lo_20=divisorMSB_hi_23 ? _divisorMSB_T_63:_divisorMSB_T_68; 
  assign _divisorMSB_T_69={divisorMSB_hi_23,divisorMSB_lo_20}; 
  assign divisorMSB_lo_21=divisorMSB_hi_19 ? _divisorMSB_T_58:_divisorMSB_T_69; 
  assign _divisorMSB_T_70={divisorMSB_hi_19,divisorMSB_lo_21}; 
  assign divisorMSB_hi_24=divisorMSB_lo_15[15:8]; 
  assign divisorMSB_lo_22=divisorMSB_lo_15[7:0]; 
  assign divisorMSB_hi_25=|divisorMSB_hi_24; 
  assign divisorMSB_hi_26=divisorMSB_hi_24[7:4]; 
  assign divisorMSB_lo_23=divisorMSB_hi_24[3:0]; 
  assign divisorMSB_hi_27=|divisorMSB_hi_26; 
  assign _divisorMSB_T_74=divisorMSB_hi_26[2] ? 2'h2:{1'b0,divisorMSB_hi_26[1]}; 
  assign _divisorMSB_T_75=divisorMSB_hi_26[3] ? 2'h3:_divisorMSB_T_74; 
  assign _divisorMSB_T_79=divisorMSB_lo_23[2] ? 2'h2:{1'b0,divisorMSB_lo_23[1]}; 
  assign _divisorMSB_T_80=divisorMSB_lo_23[3] ? 2'h3:_divisorMSB_T_79; 
  assign divisorMSB_lo_24=divisorMSB_hi_27 ? _divisorMSB_T_75:_divisorMSB_T_80; 
  assign _divisorMSB_T_81={divisorMSB_hi_27,divisorMSB_lo_24}; 
  assign divisorMSB_hi_28=divisorMSB_lo_22[7:4]; 
  assign divisorMSB_lo_25=divisorMSB_lo_22[3:0]; 
  assign divisorMSB_hi_29=|divisorMSB_hi_28; 
  assign _divisorMSB_T_85=divisorMSB_hi_28[2] ? 2'h2:{1'b0,divisorMSB_hi_28[1]}; 
  assign _divisorMSB_T_86=divisorMSB_hi_28[3] ? 2'h3:_divisorMSB_T_85; 
  assign _divisorMSB_T_90=divisorMSB_lo_25[2] ? 2'h2:{1'b0,divisorMSB_lo_25[1]}; 
  assign _divisorMSB_T_91=divisorMSB_lo_25[3] ? 2'h3:_divisorMSB_T_90; 
  assign divisorMSB_lo_26=divisorMSB_hi_29 ? _divisorMSB_T_86:_divisorMSB_T_91; 
  assign _divisorMSB_T_92={divisorMSB_hi_29,divisorMSB_lo_26}; 
  assign divisorMSB_lo_27=divisorMSB_hi_25 ? _divisorMSB_T_81:_divisorMSB_T_92; 
  assign _divisorMSB_T_93={divisorMSB_hi_25,divisorMSB_lo_27}; 
  assign divisorMSB_lo_28=divisorMSB_hi_17 ? _divisorMSB_T_70:_divisorMSB_T_93; 
  assign _divisorMSB_T_94={divisorMSB_hi_17,divisorMSB_lo_28}; 
  assign divisorMSB_lo_29=divisorMSB_hi_1 ? _divisorMSB_T_47:_divisorMSB_T_94; 
  assign divisorMSB={divisorMSB_hi_1,divisorMSB_lo_29}; 
  assign dividendMSB_hi=remainder[63:32]; 
  assign dividendMSB_lo=remainder[31:0]; 
  assign dividendMSB_hi_1=|dividendMSB_hi; 
  assign dividendMSB_hi_2=dividendMSB_hi[31:16]; 
  assign dividendMSB_lo_1=dividendMSB_hi[15:0]; 
  assign dividendMSB_hi_3=|dividendMSB_hi_2; 
  assign dividendMSB_hi_4=dividendMSB_hi_2[15:8]; 
  assign dividendMSB_lo_2=dividendMSB_hi_2[7:0]; 
  assign dividendMSB_hi_5=|dividendMSB_hi_4; 
  assign dividendMSB_hi_6=dividendMSB_hi_4[7:4]; 
  assign dividendMSB_lo_3=dividendMSB_hi_4[3:0]; 
  assign dividendMSB_hi_7=|dividendMSB_hi_6; 
  assign _dividendMSB_T_4=dividendMSB_hi_6[2] ? 2'h2:{1'b0,dividendMSB_hi_6[1]}; 
  assign _dividendMSB_T_5=dividendMSB_hi_6[3] ? 2'h3:_dividendMSB_T_4; 
  assign _dividendMSB_T_9=dividendMSB_lo_3[2] ? 2'h2:{1'b0,dividendMSB_lo_3[1]}; 
  assign _dividendMSB_T_10=dividendMSB_lo_3[3] ? 2'h3:_dividendMSB_T_9; 
  assign dividendMSB_lo_4=dividendMSB_hi_7 ? _dividendMSB_T_5:_dividendMSB_T_10; 
  assign _dividendMSB_T_11={dividendMSB_hi_7,dividendMSB_lo_4}; 
  assign dividendMSB_hi_8=dividendMSB_lo_2[7:4]; 
  assign dividendMSB_lo_5=dividendMSB_lo_2[3:0]; 
  assign dividendMSB_hi_9=|dividendMSB_hi_8; 
  assign _dividendMSB_T_15=dividendMSB_hi_8[2] ? 2'h2:{1'b0,dividendMSB_hi_8[1]}; 
  assign _dividendMSB_T_16=dividendMSB_hi_8[3] ? 2'h3:_dividendMSB_T_15; 
  assign _dividendMSB_T_20=dividendMSB_lo_5[2] ? 2'h2:{1'b0,dividendMSB_lo_5[1]}; 
  assign _dividendMSB_T_21=dividendMSB_lo_5[3] ? 2'h3:_dividendMSB_T_20; 
  assign dividendMSB_lo_6=dividendMSB_hi_9 ? _dividendMSB_T_16:_dividendMSB_T_21; 
  assign _dividendMSB_T_22={dividendMSB_hi_9,dividendMSB_lo_6}; 
  assign dividendMSB_lo_7=dividendMSB_hi_5 ? _dividendMSB_T_11:_dividendMSB_T_22; 
  assign _dividendMSB_T_23={dividendMSB_hi_5,dividendMSB_lo_7}; 
  assign dividendMSB_hi_10=dividendMSB_lo_1[15:8]; 
  assign dividendMSB_lo_8=dividendMSB_lo_1[7:0]; 
  assign dividendMSB_hi_11=|dividendMSB_hi_10; 
  assign dividendMSB_hi_12=dividendMSB_hi_10[7:4]; 
  assign dividendMSB_lo_9=dividendMSB_hi_10[3:0]; 
  assign dividendMSB_hi_13=|dividendMSB_hi_12; 
  assign _dividendMSB_T_27=dividendMSB_hi_12[2] ? 2'h2:{1'b0,dividendMSB_hi_12[1]}; 
  assign _dividendMSB_T_28=dividendMSB_hi_12[3] ? 2'h3:_dividendMSB_T_27; 
  assign _dividendMSB_T_32=dividendMSB_lo_9[2] ? 2'h2:{1'b0,dividendMSB_lo_9[1]}; 
  assign _dividendMSB_T_33=dividendMSB_lo_9[3] ? 2'h3:_dividendMSB_T_32; 
  assign dividendMSB_lo_10=dividendMSB_hi_13 ? _dividendMSB_T_28:_dividendMSB_T_33; 
  assign _dividendMSB_T_34={dividendMSB_hi_13,dividendMSB_lo_10}; 
  assign dividendMSB_hi_14=dividendMSB_lo_8[7:4]; 
  assign dividendMSB_lo_11=dividendMSB_lo_8[3:0]; 
  assign dividendMSB_hi_15=|dividendMSB_hi_14; 
  assign _dividendMSB_T_38=dividendMSB_hi_14[2] ? 2'h2:{1'b0,dividendMSB_hi_14[1]}; 
  assign _dividendMSB_T_39=dividendMSB_hi_14[3] ? 2'h3:_dividendMSB_T_38; 
  assign _dividendMSB_T_43=dividendMSB_lo_11[2] ? 2'h2:{1'b0,dividendMSB_lo_11[1]}; 
  assign _dividendMSB_T_44=dividendMSB_lo_11[3] ? 2'h3:_dividendMSB_T_43; 
  assign dividendMSB_lo_12=dividendMSB_hi_15 ? _dividendMSB_T_39:_dividendMSB_T_44; 
  assign _dividendMSB_T_45={dividendMSB_hi_15,dividendMSB_lo_12}; 
  assign dividendMSB_lo_13=dividendMSB_hi_11 ? _dividendMSB_T_34:_dividendMSB_T_45; 
  assign _dividendMSB_T_46={dividendMSB_hi_11,dividendMSB_lo_13}; 
  assign dividendMSB_lo_14=dividendMSB_hi_3 ? _dividendMSB_T_23:_dividendMSB_T_46; 
  assign _dividendMSB_T_47={dividendMSB_hi_3,dividendMSB_lo_14}; 
  assign dividendMSB_hi_16=dividendMSB_lo[31:16]; 
  assign dividendMSB_lo_15=dividendMSB_lo[15:0]; 
  assign dividendMSB_hi_17=|dividendMSB_hi_16; 
  assign dividendMSB_hi_18=dividendMSB_hi_16[15:8]; 
  assign dividendMSB_lo_16=dividendMSB_hi_16[7:0]; 
  assign dividendMSB_hi_19=|dividendMSB_hi_18; 
  assign dividendMSB_hi_20=dividendMSB_hi_18[7:4]; 
  assign dividendMSB_lo_17=dividendMSB_hi_18[3:0]; 
  assign dividendMSB_hi_21=|dividendMSB_hi_20; 
  assign _dividendMSB_T_51=dividendMSB_hi_20[2] ? 2'h2:{1'b0,dividendMSB_hi_20[1]}; 
  assign _dividendMSB_T_52=dividendMSB_hi_20[3] ? 2'h3:_dividendMSB_T_51; 
  assign _dividendMSB_T_56=dividendMSB_lo_17[2] ? 2'h2:{1'b0,dividendMSB_lo_17[1]}; 
  assign _dividendMSB_T_57=dividendMSB_lo_17[3] ? 2'h3:_dividendMSB_T_56; 
  assign dividendMSB_lo_18=dividendMSB_hi_21 ? _dividendMSB_T_52:_dividendMSB_T_57; 
  assign _dividendMSB_T_58={dividendMSB_hi_21,dividendMSB_lo_18}; 
  assign dividendMSB_hi_22=dividendMSB_lo_16[7:4]; 
  assign dividendMSB_lo_19=dividendMSB_lo_16[3:0]; 
  assign dividendMSB_hi_23=|dividendMSB_hi_22; 
  assign _dividendMSB_T_62=dividendMSB_hi_22[2] ? 2'h2:{1'b0,dividendMSB_hi_22[1]}; 
  assign _dividendMSB_T_63=dividendMSB_hi_22[3] ? 2'h3:_dividendMSB_T_62; 
  assign _dividendMSB_T_67=dividendMSB_lo_19[2] ? 2'h2:{1'b0,dividendMSB_lo_19[1]}; 
  assign _dividendMSB_T_68=dividendMSB_lo_19[3] ? 2'h3:_dividendMSB_T_67; 
  assign dividendMSB_lo_20=dividendMSB_hi_23 ? _dividendMSB_T_63:_dividendMSB_T_68; 
  assign _dividendMSB_T_69={dividendMSB_hi_23,dividendMSB_lo_20}; 
  assign dividendMSB_lo_21=dividendMSB_hi_19 ? _dividendMSB_T_58:_dividendMSB_T_69; 
  assign _dividendMSB_T_70={dividendMSB_hi_19,dividendMSB_lo_21}; 
  assign dividendMSB_hi_24=dividendMSB_lo_15[15:8]; 
  assign dividendMSB_lo_22=dividendMSB_lo_15[7:0]; 
  assign dividendMSB_hi_25=|dividendMSB_hi_24; 
  assign dividendMSB_hi_26=dividendMSB_hi_24[7:4]; 
  assign dividendMSB_lo_23=dividendMSB_hi_24[3:0]; 
  assign dividendMSB_hi_27=|dividendMSB_hi_26; 
  assign _dividendMSB_T_74=dividendMSB_hi_26[2] ? 2'h2:{1'b0,dividendMSB_hi_26[1]}; 
  assign _dividendMSB_T_75=dividendMSB_hi_26[3] ? 2'h3:_dividendMSB_T_74; 
  assign _dividendMSB_T_79=dividendMSB_lo_23[2] ? 2'h2:{1'b0,dividendMSB_lo_23[1]}; 
  assign _dividendMSB_T_80=dividendMSB_lo_23[3] ? 2'h3:_dividendMSB_T_79; 
  assign dividendMSB_lo_24=dividendMSB_hi_27 ? _dividendMSB_T_75:_dividendMSB_T_80; 
  assign _dividendMSB_T_81={dividendMSB_hi_27,dividendMSB_lo_24}; 
  assign dividendMSB_hi_28=dividendMSB_lo_22[7:4]; 
  assign dividendMSB_lo_25=dividendMSB_lo_22[3:0]; 
  assign dividendMSB_hi_29=|dividendMSB_hi_28; 
  assign _dividendMSB_T_85=dividendMSB_hi_28[2] ? 2'h2:{1'b0,dividendMSB_hi_28[1]}; 
  assign _dividendMSB_T_86=dividendMSB_hi_28[3] ? 2'h3:_dividendMSB_T_85; 
  assign _dividendMSB_T_90=dividendMSB_lo_25[2] ? 2'h2:{1'b0,dividendMSB_lo_25[1]}; 
  assign _dividendMSB_T_91=dividendMSB_lo_25[3] ? 2'h3:_dividendMSB_T_90; 
  assign dividendMSB_lo_26=dividendMSB_hi_29 ? _dividendMSB_T_86:_dividendMSB_T_91; 
  assign _dividendMSB_T_92={dividendMSB_hi_29,dividendMSB_lo_26}; 
  assign dividendMSB_lo_27=dividendMSB_hi_25 ? _dividendMSB_T_81:_dividendMSB_T_92; 
  assign _dividendMSB_T_93={dividendMSB_hi_25,dividendMSB_lo_27}; 
  assign dividendMSB_lo_28=dividendMSB_hi_17 ? _dividendMSB_T_70:_dividendMSB_T_93; 
  assign _dividendMSB_T_94={dividendMSB_hi_17,dividendMSB_lo_28}; 
  assign dividendMSB_lo_29=dividendMSB_hi_1 ? _dividendMSB_T_47:_dividendMSB_T_94; 
  assign dividendMSB={dividendMSB_hi_1,dividendMSB_lo_29}; 
  assign _eOutPos_T_1=dividendMSB-divisorMSB; 
  assign eOutPos=~_eOutPos_T_1; 
  assign _eOut_T_11=_divby0_T&~divby0; 
  assign _eOut_T_12=eOutPos>=6'h1; 
  assign eOut_1=_eOut_T_11&_eOut_T_12; 
  assign _GEN_39={63'b0,remainder[63:0]}; 
  assign _remainder_T_2=_GEN_39<<eOutPos; 
  assign _GEN_16=eOut_1 ? {2'b0,_remainder_T_2}:unrolls_0; 
  assign _T_33=divby0&~isHi; 
  assign _T_34=io_resp_ready&io_resp_valid; 
  assign _T_35=_T_34|io_kill; 
  assign _T_36=io_req_ready&io_req_valid; 
  assign _state_T_1=lhs_sign|rhs_sign; 
  assign _count_T_7=cmdMul&~io_req_bits_dw; 
  assign _count_T_8=_count_T_7 ? 3'h4:3'h0; 
  assign _neg_out_T=lhs_sign!=rhs_sign; 
  assign _divisor_T={rhs_sign,hi_1,lo_1}; 
  assign _outMul_T_1=state&3'h1; 
  assign outMul=_outMul_T_1==3'h0; 
  assign _loOut_T_3=~req_dw&outMul; 
  assign loOut=_loOut_T_3 ? result[63:32]:result[31:0]; 
  assign _hiOut_T_4=loOut[31] ? 32'hffffffff:32'h0; 
  assign hiOut=req_dw ? result[63:32]:_hiOut_T_4; 
  assign _io_resp_valid_T=state==3'h6; 
  assign _io_resp_valid_T_1=state==3'h7; 
  assign io_req_ready=state==3'h0; 
  assign io_resp_valid=_io_resp_valid_T|_io_resp_valid_T_1; 
  assign io_resp_bits_data={hiOut,loOut}; 
  assign io_resp_bits_tag=req_tag; 
  assign MulDiv_cov_read_addr=MulDiv_state; 
  assign MulDiv_cov_read_data=MulDiv_cov[MulDiv_cov_read_addr]; 
  assign MulDiv_cov_write_data=1'h1; 
  assign MulDiv_cov_write_addr=MulDiv_state; 
  assign MulDiv_cov_write_mask=1'h1; 
  assign MulDiv_cov_write_en=1'h1; 
  assign mux_cond_0=dividendMSB_hi_13; 
  assign mux_cond_1=dividendMSB_lo_19[3]; 
  assign mux_cond_2=divisorMSB_hi_21; 
  assign mux_cond_3=dividendMSB_hi_28[3]; 
  assign mux_cond_4=divisorMSB_hi_3; 
  assign mux_cond_5=divisorMSB_lo_5[2]; 
  assign mux_cond_6=dividendMSB_lo_19[2]; 
  assign mux_cond_7=divisorMSB_hi_14[2]; 
  assign mux_cond_8=divisorMSB_hi_26[3]; 
  assign mux_cond_9=dividendMSB_hi_7; 
  assign mux_cond_10=divisorMSB_hi_28[3]; 
  assign mux_cond_11=dividendMSB_hi_20[2]; 
  assign mux_cond_12=dividendMSB_hi_8[3]; 
  assign mux_cond_13=dividendMSB_hi_27; 
  assign mux_cond_14=divisorMSB_lo_19[2]; 
  assign mux_cond_15=divisorMSB_lo_9[3]; 
  assign mux_cond_16=dividendMSB_lo_3[3]; 
  assign mux_cond_17=dividendMSB_hi_22[2]; 
  assign mux_cond_18=divisorMSB_hi_6[3]; 
  assign mux_cond_19=dividendMSB_lo_23[2]; 
  assign mux_cond_20=divisorMSB_hi_26[2]; 
  assign mux_cond_21=dividendMSB_hi_6[3]; 
  assign mux_cond_22=divisorMSB_lo_19[3]; 
  assign mux_cond_23=divisorMSB_lo_17[2]; 
  assign mux_cond_24=dividendMSB_lo_3[2]; 
  assign mux_cond_25=divisorMSB_hi_29; 
  assign mux_cond_26=dividendMSB_lo_17[2]; 
  assign mux_cond_27=dividendMSB_lo_25[3]; 
  assign mux_cond_28=divisorMSB_hi_7; 
  assign mux_cond_29=dividendMSB_hi_29; 
  assign mux_cond_30=divisorMSB_lo_9[2]; 
  assign mux_cond_31=dividendMSB_hi_9; 
  assign mux_cond_32=divisorMSB_hi_28[2]; 
  assign mux_cond_33=divisorMSB_hi_25; 
  assign mux_cond_34=divisorMSB_lo_25[2]; 
  assign mux_cond_35=divisorMSB_hi_11; 
  assign mux_cond_36=divisorMSB_lo_23[2]; 
  assign mux_cond_37=dividendMSB_hi_1; 
  assign mux_cond_38=dividendMSB_lo_9[2]; 
  assign mux_cond_39=divisorMSB_hi_17; 
  assign mux_cond_40=dividendMSB_lo_17[3]; 
  assign mux_cond_41=divisorMSB_lo_11[2]; 
  assign mux_cond_42=divisorMSB_hi_15; 
  assign mux_cond_43=divisorMSB_hi_14[3]; 
  assign mux_cond_44=divisor[63]; 
  assign mux_cond_45=divisorMSB_hi_6[2]; 
  assign mux_cond_46=divisorMSB_hi_8[3]; 
  assign mux_cond_47=divisorMSB_hi_20[3]; 
  assign mux_cond_48=dividendMSB_hi_28[2]; 
  assign mux_cond_49=unrolls_less; 
  assign mux_cond_50=divisorMSB_hi_8[2]; 
  assign mux_cond_51=divisorMSB_hi_23; 
  assign mux_cond_52=dividendMSB_lo_23[3]; 
  assign mux_cond_53=divisorMSB_hi_22[3]; 
  assign mux_cond_54=divisorMSB_lo_3[2]; 
  assign mux_cond_55=divisorMSB_lo_25[3]; 
  assign mux_cond_56=divisorMSB_lo_23[3]; 
  assign mux_cond_57=divisorMSB_hi_27; 
  assign mux_cond_58=divisorMSB_hi_12[2]; 
  assign mux_cond_59=dividendMSB_lo_11[3]; 
  assign mux_cond_60=divisorMSB_lo_3[3]; 
  assign mux_cond_61=dividendMSB_hi_21; 
  assign mux_cond_62=dividendMSB_hi_12[3]; 
  assign mux_cond_63=dividendMSB_hi_14[3]; 
  assign mux_cond_64=divisorMSB_hi_20[2]; 
  assign mux_cond_65=dividendMSB_lo_5[2]; 
  assign mux_cond_66=dividendMSB_hi_17; 
  assign mux_cond_67=dividendMSB_hi_8[2]; 
  assign mux_cond_68=remainder[63]; 
  assign mux_cond_69=dividendMSB_hi_12[2]; 
  assign mux_cond_70=divisorMSB_hi_22[2]; 
  assign mux_cond_71=dividendMSB_hi_19; 
  assign mux_cond_72=dividendMSB_hi_5; 
  assign mux_cond_73=loOut[31]; 
  assign mux_cond_74=dividendMSB_hi_14[2]; 
  assign mux_cond_75=divisorMSB_hi_12[3]; 
  assign mux_cond_76=divisorMSB_hi_5; 
  assign mux_cond_77=divisorMSB_lo_11[3]; 
  assign mux_cond_78=divisorMSB_lo_5[3]; 
  assign mux_cond_79=dividendMSB_lo_5[3]; 
  assign mux_cond_80=dividendMSB_hi_26[3]; 
  assign mux_cond_81=dividendMSB_hi_15; 
  assign mux_cond_82=dividendMSB_hi_25; 
  assign mux_cond_83=divisorMSB_hi_13; 
  assign mux_cond_84=dividendMSB_hi_3; 
  assign mux_cond_85=dividendMSB_hi_23; 
  assign mux_cond_86=dividendMSB_lo_9[3]; 
  assign mux_cond_87=divisorMSB_lo_17[3]; 
  assign mux_cond_88=dividendMSB_hi_22[3]; 
  assign mux_cond_89=dividendMSB_hi_6[2]; 
  assign mux_cond_90=dividendMSB_hi_11; 
  assign mux_cond_91=divisorMSB_hi_19; 
  assign mux_cond_92=dividendMSB_lo_11[2]; 
  assign mux_cond_93=divisorMSB_hi_9; 
  assign mux_cond_94=dividendMSB_lo_25[2]; 
  assign mux_cond_95=divisorMSB_hi_1; 
  assign mux_cond_96=dividendMSB_hi_20[3]; 
  assign mux_cond_97=dividendMSB_hi_26[2]; 
  assign isHi_shl={isHi,4'h0}; 
  assign isHi_pad={15'h0,isHi_shl}; 
  assign neg_out_shl={neg_out,12'h0}; 
  assign neg_out_pad={7'h0,neg_out_shl}; 
  assign req_dw_shl={req_dw,4'h0}; 
  assign req_dw_pad={15'h0,req_dw_shl}; 
  assign state_shl={state,8'h0}; 
  assign state_pad={9'h0,state_shl}; 
  assign resHi_shl={resHi,1'h0}; 
  assign resHi_pad={18'h0,resHi_shl}; 
  assign mux_cond_0_shl={mux_cond_0,12'h0}; 
  assign mux_cond_0_pad={7'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,1'h0}; 
  assign mux_cond_1_pad={18'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl=mux_cond_2; 
  assign mux_cond_2_pad={19'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,12'h0}; 
  assign mux_cond_3_pad={7'h0,mux_cond_3_shl}; 
  assign mux_cond_4_shl={mux_cond_4,15'h0}; 
  assign mux_cond_4_pad={4'h0,mux_cond_4_shl}; 
  assign mux_cond_5_shl={mux_cond_5,11'h0}; 
  assign mux_cond_5_pad={8'h0,mux_cond_5_shl}; 
  assign mux_cond_6_shl={mux_cond_6,7'h0}; 
  assign mux_cond_6_pad={12'h0,mux_cond_6_shl}; 
  assign mux_cond_7_shl={mux_cond_7,17'h0}; 
  assign mux_cond_7_pad={2'h0,mux_cond_7_shl}; 
  assign mux_cond_8_shl={mux_cond_8,11'h0}; 
  assign mux_cond_8_pad={8'h0,mux_cond_8_shl}; 
  assign mux_cond_9_shl={mux_cond_9,15'h0}; 
  assign mux_cond_9_pad={4'h0,mux_cond_9_shl}; 
  assign mux_cond_10_shl={mux_cond_10,13'h0}; 
  assign mux_cond_10_pad={6'h0,mux_cond_10_shl}; 
  assign mux_cond_11_shl=mux_cond_11; 
  assign mux_cond_11_pad={19'h0,mux_cond_11_shl}; 
  assign mux_cond_12_shl={mux_cond_12,7'h0}; 
  assign mux_cond_12_pad={12'h0,mux_cond_12_shl}; 
  assign mux_cond_13_shl={mux_cond_13,13'h0}; 
  assign mux_cond_13_pad={6'h0,mux_cond_13_shl}; 
  assign mux_cond_14_shl=mux_cond_14; 
  assign mux_cond_14_pad={19'h0,mux_cond_14_shl}; 
  assign mux_cond_15_shl={mux_cond_15,9'h0}; 
  assign mux_cond_15_pad={10'h0,mux_cond_15_shl}; 
  assign mux_cond_16_shl={mux_cond_16,8'h0}; 
  assign mux_cond_16_pad={11'h0,mux_cond_16_shl}; 
  assign mux_cond_17_shl={mux_cond_17,8'h0}; 
  assign mux_cond_17_pad={11'h0,mux_cond_17_shl}; 
  assign mux_cond_18_shl={mux_cond_18,8'h0}; 
  assign mux_cond_18_pad={11'h0,mux_cond_18_shl}; 
  assign mux_cond_19_shl={mux_cond_19,2'h0}; 
  assign mux_cond_19_pad={17'h0,mux_cond_19_shl}; 
  assign mux_cond_20_shl={mux_cond_20,16'h0}; 
  assign mux_cond_20_pad={3'h0,mux_cond_20_shl}; 
  assign mux_cond_21_shl={mux_cond_21,6'h0}; 
  assign mux_cond_21_pad={13'h0,mux_cond_21_shl}; 
  assign mux_cond_22_shl={mux_cond_22,11'h0}; 
  assign mux_cond_22_pad={8'h0,mux_cond_22_shl}; 
  assign mux_cond_23_shl=mux_cond_23; 
  assign mux_cond_23_pad={19'h0,mux_cond_23_shl}; 
  assign mux_cond_24_shl={mux_cond_24,6'h0}; 
  assign mux_cond_24_pad={13'h0,mux_cond_24_shl}; 
  assign mux_cond_25_shl={mux_cond_25,12'h0}; 
  assign mux_cond_25_pad={7'h0,mux_cond_25_shl}; 
  assign mux_cond_26_shl={mux_cond_26,4'h0}; 
  assign mux_cond_26_pad={15'h0,mux_cond_26_shl}; 
  assign mux_cond_27_shl={mux_cond_27,11'h0}; 
  assign mux_cond_27_pad={8'h0,mux_cond_27_shl}; 
  assign mux_cond_28_shl={mux_cond_28,6'h0}; 
  assign mux_cond_28_pad={13'h0,mux_cond_28_shl}; 
  assign mux_cond_29_shl={mux_cond_29,12'h0}; 
  assign mux_cond_29_pad={7'h0,mux_cond_29_shl}; 
  assign mux_cond_30_shl={mux_cond_30,1'h0}; 
  assign mux_cond_30_pad={18'h0,mux_cond_30_shl}; 
  assign mux_cond_31_shl={mux_cond_31,11'h0}; 
  assign mux_cond_31_pad={8'h0,mux_cond_31_shl}; 
  assign mux_cond_32_shl={mux_cond_32,6'h0}; 
  assign mux_cond_32_pad={13'h0,mux_cond_32_shl}; 
  assign mux_cond_33_shl={mux_cond_33,5'h0}; 
  assign mux_cond_33_pad={14'h0,mux_cond_33_shl}; 
  assign mux_cond_34_shl={mux_cond_34,18'h0}; 
  assign mux_cond_34_pad={1'h0,mux_cond_34_shl}; 
  assign mux_cond_35_shl={mux_cond_35,12'h0}; 
  assign mux_cond_35_pad={7'h0,mux_cond_35_shl}; 
  assign mux_cond_36_shl=mux_cond_36; 
  assign mux_cond_36_pad={19'h0,mux_cond_36_shl}; 
  assign mux_cond_37_shl={mux_cond_37,8'h0}; 
  assign mux_cond_37_pad={11'h0,mux_cond_37_shl}; 
  assign mux_cond_38_shl={mux_cond_38,5'h0}; 
  assign mux_cond_38_pad={14'h0,mux_cond_38_shl}; 
  assign mux_cond_39_shl={mux_cond_39,16'h0}; 
  assign mux_cond_39_pad={3'h0,mux_cond_39_shl}; 
  assign mux_cond_40_shl={mux_cond_40,3'h0}; 
  assign mux_cond_40_pad={16'h0,mux_cond_40_shl}; 
  assign mux_cond_41_shl={mux_cond_41,9'h0}; 
  assign mux_cond_41_pad={10'h0,mux_cond_41_shl}; 
  assign mux_cond_42_shl={mux_cond_42,15'h0}; 
  assign mux_cond_42_pad={4'h0,mux_cond_42_shl}; 
  assign mux_cond_43_shl={mux_cond_43,13'h0}; 
  assign mux_cond_43_pad={6'h0,mux_cond_43_shl}; 
  assign mux_cond_44_shl={mux_cond_44,12'h0}; 
  assign mux_cond_44_pad={7'h0,mux_cond_44_shl}; 
  assign mux_cond_45_shl=mux_cond_45; 
  assign mux_cond_45_pad={19'h0,mux_cond_45_shl}; 
  assign mux_cond_46_shl={mux_cond_46,3'h0}; 
  assign mux_cond_46_pad={16'h0,mux_cond_46_shl}; 
  assign mux_cond_47_shl={mux_cond_47,14'h0}; 
  assign mux_cond_47_pad={5'h0,mux_cond_47_shl}; 
  assign mux_cond_48_shl={mux_cond_48,16'h0}; 
  assign mux_cond_48_pad={3'h0,mux_cond_48_shl}; 
  assign mux_cond_49_shl={mux_cond_49,18'h0}; 
  assign mux_cond_49_pad={1'h0,mux_cond_49_shl}; 
  assign mux_cond_50_shl=mux_cond_50; 
  assign mux_cond_50_pad={19'h0,mux_cond_50_shl}; 
  assign mux_cond_51_shl={mux_cond_51,7'h0}; 
  assign mux_cond_51_pad={12'h0,mux_cond_51_shl}; 
  assign mux_cond_52_shl=mux_cond_52; 
  assign mux_cond_52_pad={19'h0,mux_cond_52_shl}; 
  assign mux_cond_53_shl={mux_cond_53,19'h0}; 
  assign mux_cond_53_pad=mux_cond_53_shl; 
  assign mux_cond_54_shl={mux_cond_54,10'h0}; 
  assign mux_cond_54_pad={9'h0,mux_cond_54_shl}; 
  assign mux_cond_55_shl={mux_cond_55,13'h0}; 
  assign mux_cond_55_pad={6'h0,mux_cond_55_shl}; 
  assign mux_cond_56_shl={mux_cond_56,9'h0}; 
  assign mux_cond_56_pad={10'h0,mux_cond_56_shl}; 
  assign mux_cond_57_shl={mux_cond_57,6'h0}; 
  assign mux_cond_57_pad={13'h0,mux_cond_57_shl}; 
  assign mux_cond_58_shl={mux_cond_58,17'h0}; 
  assign mux_cond_58_pad={2'h0,mux_cond_58_shl}; 
  assign mux_cond_59_shl={mux_cond_59,19'h0}; 
  assign mux_cond_59_pad=mux_cond_59_shl; 
  assign mux_cond_60_shl={mux_cond_60,3'h0}; 
  assign mux_cond_60_pad={16'h0,mux_cond_60_shl}; 
  assign mux_cond_61_shl={mux_cond_61,14'h0}; 
  assign mux_cond_61_pad={5'h0,mux_cond_61_shl}; 
  assign mux_cond_62_shl={mux_cond_62,4'h0}; 
  assign mux_cond_62_pad={15'h0,mux_cond_62_shl}; 
  assign mux_cond_63_shl=mux_cond_63; 
  assign mux_cond_63_pad={19'h0,mux_cond_63_shl}; 
  assign mux_cond_64_shl={mux_cond_64,10'h0}; 
  assign mux_cond_64_pad={9'h0,mux_cond_64_shl}; 
  assign mux_cond_65_shl={mux_cond_65,17'h0}; 
  assign mux_cond_65_pad={2'h0,mux_cond_65_shl}; 
  assign mux_cond_66_shl={mux_cond_66,9'h0}; 
  assign mux_cond_66_pad={10'h0,mux_cond_66_shl}; 
  assign mux_cond_67_shl={mux_cond_67,6'h0}; 
  assign mux_cond_67_pad={13'h0,mux_cond_67_shl}; 
  assign mux_cond_68_shl={mux_cond_68,19'h0}; 
  assign mux_cond_68_pad=mux_cond_68_shl; 
  assign mux_cond_69_shl={mux_cond_69,10'h0}; 
  assign mux_cond_69_pad={9'h0,mux_cond_69_shl}; 
  assign mux_cond_70_shl={mux_cond_70,10'h0}; 
  assign mux_cond_70_pad={9'h0,mux_cond_70_shl}; 
  assign mux_cond_71_shl={mux_cond_71,13'h0}; 
  assign mux_cond_71_pad={6'h0,mux_cond_71_shl}; 
  assign mux_cond_72_shl={mux_cond_72,18'h0}; 
  assign mux_cond_72_pad={1'h0,mux_cond_72_shl}; 
  assign mux_cond_73_shl={mux_cond_73,12'h0}; 
  assign mux_cond_73_pad={7'h0,mux_cond_73_shl}; 
  assign mux_cond_74_shl={mux_cond_74,13'h0}; 
  assign mux_cond_74_pad={6'h0,mux_cond_74_shl}; 
  assign mux_cond_75_shl={mux_cond_75,13'h0}; 
  assign mux_cond_75_pad={6'h0,mux_cond_75_shl}; 
  assign mux_cond_76_shl={mux_cond_76,13'h0}; 
  assign mux_cond_76_pad={6'h0,mux_cond_76_shl}; 
  assign mux_cond_77_shl={mux_cond_77,13'h0}; 
  assign mux_cond_77_pad={6'h0,mux_cond_77_shl}; 
  assign mux_cond_78_shl={mux_cond_78,17'h0}; 
  assign mux_cond_78_pad={2'h0,mux_cond_78_shl}; 
  assign mux_cond_79_shl={mux_cond_79,12'h0}; 
  assign mux_cond_79_pad={7'h0,mux_cond_79_shl}; 
  assign mux_cond_80_shl={mux_cond_80,17'h0}; 
  assign mux_cond_80_pad={2'h0,mux_cond_80_shl}; 
  assign mux_cond_81_shl={mux_cond_81,13'h0}; 
  assign mux_cond_81_pad={6'h0,mux_cond_81_shl}; 
  assign mux_cond_82_shl={mux_cond_82,12'h0}; 
  assign mux_cond_82_pad={7'h0,mux_cond_82_shl}; 
  assign mux_cond_83_shl={mux_cond_83,4'h0}; 
  assign mux_cond_83_pad={15'h0,mux_cond_83_shl}; 
  assign mux_cond_84_shl={mux_cond_84,16'h0}; 
  assign mux_cond_84_pad={3'h0,mux_cond_84_shl}; 
  assign mux_cond_85_shl={mux_cond_85,9'h0}; 
  assign mux_cond_85_pad={10'h0,mux_cond_85_shl}; 
  assign mux_cond_86_shl={mux_cond_86,10'h0}; 
  assign mux_cond_86_pad={9'h0,mux_cond_86_shl}; 
  assign mux_cond_87_shl={mux_cond_87,2'h0}; 
  assign mux_cond_87_pad={17'h0,mux_cond_87_shl}; 
  assign mux_cond_88_shl={mux_cond_88,6'h0}; 
  assign mux_cond_88_pad={13'h0,mux_cond_88_shl}; 
  assign mux_cond_89_shl={mux_cond_89,11'h0}; 
  assign mux_cond_89_pad={8'h0,mux_cond_89_shl}; 
  assign mux_cond_90_shl={mux_cond_90,7'h0}; 
  assign mux_cond_90_pad={12'h0,mux_cond_90_shl}; 
  assign mux_cond_91_shl={mux_cond_91,16'h0}; 
  assign mux_cond_91_pad={3'h0,mux_cond_91_shl}; 
  assign mux_cond_92_shl={mux_cond_92,17'h0}; 
  assign mux_cond_92_pad={2'h0,mux_cond_92_shl}; 
  assign mux_cond_93_shl={mux_cond_93,5'h0}; 
  assign mux_cond_93_pad={14'h0,mux_cond_93_shl}; 
  assign mux_cond_94_shl={mux_cond_94,18'h0}; 
  assign mux_cond_94_pad={1'h0,mux_cond_94_shl}; 
  assign mux_cond_95_shl={mux_cond_95,1'h0}; 
  assign mux_cond_95_pad={18'h0,mux_cond_95_shl}; 
  assign mux_cond_96_shl={mux_cond_96,17'h0}; 
  assign mux_cond_96_pad={2'h0,mux_cond_96_shl}; 
  assign mux_cond_97_shl={mux_cond_97,1'h0}; 
  assign mux_cond_97_pad={18'h0,mux_cond_97_shl}; 
  assign MulDiv_xor64=neg_out_pad^req_dw_pad; 
  assign MulDiv_xor31=isHi_pad^MulDiv_xor64; 
  assign MulDiv_xor66=resHi_pad^mux_cond_0_pad; 
  assign MulDiv_xor32=state_pad^MulDiv_xor66; 
  assign MulDiv_xor15=MulDiv_xor31^MulDiv_xor32; 
  assign MulDiv_xor68=mux_cond_2_pad^mux_cond_3_pad; 
  assign MulDiv_xor33=mux_cond_1_pad^MulDiv_xor68; 
  assign MulDiv_xor70=mux_cond_5_pad^mux_cond_6_pad; 
  assign MulDiv_xor34=mux_cond_4_pad^MulDiv_xor70; 
  assign MulDiv_xor16=MulDiv_xor33^MulDiv_xor34; 
  assign MulDiv_xor7=MulDiv_xor15^MulDiv_xor16; 
  assign MulDiv_xor72=mux_cond_8_pad^mux_cond_9_pad; 
  assign MulDiv_xor35=mux_cond_7_pad^MulDiv_xor72; 
  assign MulDiv_xor74=mux_cond_11_pad^mux_cond_12_pad; 
  assign MulDiv_xor36=mux_cond_10_pad^MulDiv_xor74; 
  assign MulDiv_xor17=MulDiv_xor35^MulDiv_xor36; 
  assign MulDiv_xor76=mux_cond_14_pad^mux_cond_15_pad; 
  assign MulDiv_xor37=mux_cond_13_pad^MulDiv_xor76; 
  assign MulDiv_xor77=mux_cond_16_pad^mux_cond_17_pad; 
  assign MulDiv_xor78=mux_cond_18_pad^mux_cond_19_pad; 
  assign MulDiv_xor38=MulDiv_xor77^MulDiv_xor78; 
  assign MulDiv_xor18=MulDiv_xor37^MulDiv_xor38; 
  assign MulDiv_xor8=MulDiv_xor17^MulDiv_xor18; 
  assign MulDiv_xor3=MulDiv_xor7^MulDiv_xor8; 
  assign MulDiv_xor80=mux_cond_21_pad^mux_cond_22_pad; 
  assign MulDiv_xor39=mux_cond_20_pad^MulDiv_xor80; 
  assign MulDiv_xor82=mux_cond_24_pad^mux_cond_25_pad; 
  assign MulDiv_xor40=mux_cond_23_pad^MulDiv_xor82; 
  assign MulDiv_xor19=MulDiv_xor39^MulDiv_xor40; 
  assign MulDiv_xor84=mux_cond_27_pad^mux_cond_28_pad; 
  assign MulDiv_xor41=mux_cond_26_pad^MulDiv_xor84; 
  assign MulDiv_xor85=mux_cond_29_pad^mux_cond_30_pad; 
  assign MulDiv_xor86=mux_cond_31_pad^mux_cond_32_pad; 
  assign MulDiv_xor42=MulDiv_xor85^MulDiv_xor86; 
  assign MulDiv_xor20=MulDiv_xor41^MulDiv_xor42; 
  assign MulDiv_xor9=MulDiv_xor19^MulDiv_xor20; 
  assign MulDiv_xor88=mux_cond_34_pad^mux_cond_35_pad; 
  assign MulDiv_xor43=mux_cond_33_pad^MulDiv_xor88; 
  assign MulDiv_xor90=mux_cond_37_pad^mux_cond_38_pad; 
  assign MulDiv_xor44=mux_cond_36_pad^MulDiv_xor90; 
  assign MulDiv_xor21=MulDiv_xor43^MulDiv_xor44; 
  assign MulDiv_xor92=mux_cond_40_pad^mux_cond_41_pad; 
  assign MulDiv_xor45=mux_cond_39_pad^MulDiv_xor92; 
  assign MulDiv_xor93=mux_cond_42_pad^mux_cond_43_pad; 
  assign MulDiv_xor94=mux_cond_44_pad^mux_cond_45_pad; 
  assign MulDiv_xor46=MulDiv_xor93^MulDiv_xor94; 
  assign MulDiv_xor22=MulDiv_xor45^MulDiv_xor46; 
  assign MulDiv_xor10=MulDiv_xor21^MulDiv_xor22; 
  assign MulDiv_xor4=MulDiv_xor9^MulDiv_xor10; 
  assign MulDiv_xor1=MulDiv_xor3^MulDiv_xor4; 
  assign MulDiv_xor96=mux_cond_47_pad^mux_cond_48_pad; 
  assign MulDiv_xor47=mux_cond_46_pad^MulDiv_xor96; 
  assign MulDiv_xor98=mux_cond_50_pad^mux_cond_51_pad; 
  assign MulDiv_xor48=mux_cond_49_pad^MulDiv_xor98; 
  assign MulDiv_xor23=MulDiv_xor47^MulDiv_xor48; 
  assign MulDiv_xor100=mux_cond_53_pad^mux_cond_54_pad; 
  assign MulDiv_xor49=mux_cond_52_pad^MulDiv_xor100; 
  assign MulDiv_xor101=mux_cond_55_pad^mux_cond_56_pad; 
  assign MulDiv_xor102=mux_cond_57_pad^mux_cond_58_pad; 
  assign MulDiv_xor50=MulDiv_xor101^MulDiv_xor102; 
  assign MulDiv_xor24=MulDiv_xor49^MulDiv_xor50; 
  assign MulDiv_xor11=MulDiv_xor23^MulDiv_xor24; 
  assign MulDiv_xor104=mux_cond_60_pad^mux_cond_61_pad; 
  assign MulDiv_xor51=mux_cond_59_pad^MulDiv_xor104; 
  assign MulDiv_xor106=mux_cond_63_pad^mux_cond_64_pad; 
  assign MulDiv_xor52=mux_cond_62_pad^MulDiv_xor106; 
  assign MulDiv_xor25=MulDiv_xor51^MulDiv_xor52; 
  assign MulDiv_xor108=mux_cond_66_pad^mux_cond_67_pad; 
  assign MulDiv_xor53=mux_cond_65_pad^MulDiv_xor108; 
  assign MulDiv_xor109=mux_cond_68_pad^mux_cond_69_pad; 
  assign MulDiv_xor110=mux_cond_70_pad^mux_cond_71_pad; 
  assign MulDiv_xor54=MulDiv_xor109^MulDiv_xor110; 
  assign MulDiv_xor26=MulDiv_xor53^MulDiv_xor54; 
  assign MulDiv_xor12=MulDiv_xor25^MulDiv_xor26; 
  assign MulDiv_xor5=MulDiv_xor11^MulDiv_xor12; 
  assign MulDiv_xor112=mux_cond_73_pad^mux_cond_74_pad; 
  assign MulDiv_xor55=mux_cond_72_pad^MulDiv_xor112; 
  assign MulDiv_xor114=mux_cond_76_pad^mux_cond_77_pad; 
  assign MulDiv_xor56=mux_cond_75_pad^MulDiv_xor114; 
  assign MulDiv_xor27=MulDiv_xor55^MulDiv_xor56; 
  assign MulDiv_xor116=mux_cond_79_pad^mux_cond_80_pad; 
  assign MulDiv_xor57=mux_cond_78_pad^MulDiv_xor116; 
  assign MulDiv_xor117=mux_cond_81_pad^mux_cond_82_pad; 
  assign MulDiv_xor118=mux_cond_83_pad^mux_cond_84_pad; 
  assign MulDiv_xor58=MulDiv_xor117^MulDiv_xor118; 
  assign MulDiv_xor28=MulDiv_xor57^MulDiv_xor58; 
  assign MulDiv_xor13=MulDiv_xor27^MulDiv_xor28; 
  assign MulDiv_xor120=mux_cond_86_pad^mux_cond_87_pad; 
  assign MulDiv_xor59=mux_cond_85_pad^MulDiv_xor120; 
  assign MulDiv_xor122=mux_cond_89_pad^mux_cond_90_pad; 
  assign MulDiv_xor60=mux_cond_88_pad^MulDiv_xor122; 
  assign MulDiv_xor29=MulDiv_xor59^MulDiv_xor60; 
  assign MulDiv_xor124=mux_cond_92_pad^mux_cond_93_pad; 
  assign MulDiv_xor61=mux_cond_91_pad^MulDiv_xor124; 
  assign MulDiv_xor125=mux_cond_94_pad^mux_cond_95_pad; 
  assign MulDiv_xor126=mux_cond_96_pad^mux_cond_97_pad; 
  assign MulDiv_xor62=MulDiv_xor125^MulDiv_xor126; 
  assign MulDiv_xor30=MulDiv_xor61^MulDiv_xor62; 
  assign MulDiv_xor14=MulDiv_xor29^MulDiv_xor30; 
  assign MulDiv_xor6=MulDiv_xor13^MulDiv_xor14; 
  assign MulDiv_xor2=MulDiv_xor5^MulDiv_xor6; 
  assign MulDiv_xor0=MulDiv_xor1^MulDiv_xor2; 
  assign io_covSum=MulDiv_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              state <=3'h0;
            end 
          else 
            if (reset)
               begin 
                 state <=3'h0;
               end 
             else 
               if (_T_36)
                  begin 
                    if (cmdMul)
                       begin 
                         state <=3'h2;
                       end 
                     else 
                       if (_state_T_1)
                          begin 
                            state <=3'h1;
                          end 
                        else 
                          begin 
                            state <=3'h3;
                          end 
                  end 
                else 
                  if (_T_35)
                     begin 
                       state <=3'h0;
                     end 
                   else 
                     if (_T_30)
                        begin 
                          if (_T_31)
                             begin 
                               if (neg_out)
                                  begin 
                                    state <=3'h5;
                                  end 
                                else 
                                  begin 
                                    state <=3'h7;
                                  end 
                             end 
                           else 
                             if (_T_27)
                                begin 
                                  if (_T_29)
                                     begin 
                                       state <=3'h6;
                                     end 
                                   else 
                                     if (_T_26)
                                        begin 
                                          state <=3'h7;
                                        end 
                                      else 
                                        if (_T_23)
                                           begin 
                                             state <=3'h3;
                                           end 
                                end 
                              else 
                                if (_T_26)
                                   begin 
                                     state <=3'h7;
                                   end 
                                 else 
                                   if (_T_23)
                                      begin 
                                        state <=3'h3;
                                      end 
                        end 
                      else 
                        if (_T_27)
                           begin 
                             if (_T_29)
                                begin 
                                  state <=3'h6;
                                end 
                              else 
                                if (_T_26)
                                   begin 
                                     state <=3'h7;
                                   end 
                                 else 
                                   if (_T_23)
                                      begin 
                                        state <=3'h3;
                                      end 
                           end 
                         else 
                           if (_T_26)
                              begin 
                                state <=3'h7;
                              end 
                            else 
                              if (_T_23)
                                 begin 
                                   state <=3'h3;
                                 end 
         if (metaReset)
            begin 
              req_dw <=1'h0;
            end 
          else 
            if (_T_36)
               begin 
                 req_dw <=io_req_bits_dw;
               end 
         if (metaReset)
            begin 
              req_tag <=5'h0;
            end 
          else 
            if (_T_36)
               begin 
                 req_tag <=io_req_bits_tag;
               end 
         if (metaReset)
            begin 
              count <=7'h0;
            end 
          else 
            if (_T_36)
               begin 
                 count <={4'b0,_count_T_8};
               end 
             else 
               if (_T_30)
                  begin 
                    if (eOut_1)
                       begin 
                         count <={1'b0,eOutPos};
                       end 
                     else 
                       begin 
                         count <=_count_T_1;
                       end 
                  end 
                else 
                  if (_T_27)
                     begin 
                       count <=_count_T_1;
                     end 
         if (metaReset)
            begin 
              neg_out <=1'h0;
            end 
          else 
            if (_T_36)
               begin 
                 if (cmdHi)
                    begin 
                      neg_out <=lhs_sign;
                    end 
                  else 
                    begin 
                      neg_out <=_neg_out_T;
                    end 
               end 
             else 
               if (_T_30)
                  begin 
                    if (_T_33)
                       begin 
                         neg_out <=1'h0;
                       end 
                  end 
         if (metaReset)
            begin 
              isHi <=1'h0;
            end 
          else 
            if (_T_36)
               begin 
                 isHi <=cmdHi;
               end 
         if (metaReset)
            begin 
              resHi <=1'h0;
            end 
          else 
            if (_T_36)
               begin 
                 resHi <=1'h0;
               end 
             else 
               if (_T_30)
                  begin 
                    if (_T_31)
                       begin 
                         resHi <=isHi;
                       end 
                     else 
                       if (_T_27)
                          begin 
                            if (_T_29)
                               begin 
                                 resHi <=isHi;
                               end 
                             else 
                               if (_T_26)
                                  begin 
                                    resHi <=1'h0;
                                  end 
                          end 
                        else 
                          if (_T_26)
                             begin 
                               resHi <=1'h0;
                             end 
                  end 
                else 
                  if (_T_27)
                     begin 
                       if (_T_29)
                          begin 
                            resHi <=isHi;
                          end 
                        else 
                          if (_T_26)
                             begin 
                               resHi <=1'h0;
                             end 
                     end 
                   else 
                     if (_T_26)
                        begin 
                          resHi <=1'h0;
                        end 
         if (metaReset)
            begin 
              divisor <=65'h0;
            end 
          else 
            if (_T_36)
               begin 
                 divisor <=_divisor_T;
               end 
             else 
               if (_T_23)
                  begin 
                    if (divisor[63])
                       begin 
                         divisor <=subtractor;
                       end 
                  end 
         if (metaReset)
            begin 
              remainder <=130'h0;
            end 
          else 
            if (_T_36)
               begin 
                 remainder <={66'b0,lhs_in};
               end 
             else 
               if (_T_30)
                  begin 
                    remainder <={1'b0,_GEN_16};
                  end 
                else 
                  if (_T_27)
                     begin 
                       remainder <=_remainder_T;
                     end 
                   else 
                     if (_T_26)
                        begin 
                          remainder <={66'b0,negated_remainder};
                        end 
                      else 
                        if (_T_23)
                           begin 
                             if (remainder[63])
                                begin 
                                  remainder <={66'b0,negated_remainder};
                                end 
                           end 
         MulDiv_state <=MulDiv_xor0;
         if (!(MulDiv_cov_read_data))
            begin 
              MulDiv_covSum <=MulDiv_covSum+1'h1;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (MulDiv_cov_write_en&MulDiv_cov_write_mask)
            begin 
              MulDiv_cov [MulDiv_cov_write_addr]<=MulDiv_cov_write_data;
            end 
       end
  
endmodule
 
module PlusArgTimeout (
  input clock,
  input reset,
  input [31:0] io_count,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [31:0] plusarg_reader_out ;  
   wire _T ;  
   wire _T_1 ;  
   wire _T_3 ;  
   wire [29:0] PlusArgTimeout_covSum ;  
   wire stopEn0 ;  
   wire plusarg_reader_metaAssert_wire ;  
   wire PlusArgTimeout_or0 ;  
   reg PlusArgTimeout_metaAssert ;  
   reg [31:0] _RAND_0 ;  
  assign _T=plusarg_reader_out>32'h0; 
  assign _T_1=io_count<plusarg_reader_out; 
  assign _T_3=_T_1|reset; 
  assign PlusArgTimeout_covSum=30'h0; 
  assign io_covSum=PlusArgTimeout_covSum; 
  assign stopEn0=_T&~_T_3; 
  assign PlusArgTimeout_or0=stopEn0|plusarg_reader_metaAssert_wire; 
  assign metaAssert=PlusArgTimeout_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (_T&~_T_3)
            begin $display("Assertion failed: Timeout exceeded: Kill the emulation after INT rdtime cycles. Off if 0.\n    at PlusArg.scala:64 assert (io.count < max, s\"Timeout exceeded: $docstring\")\n");
            end 
         if (_T&~_T_3)
            begin $display("fatal");
            end 
         if (metaReset)
            begin 
              PlusArgTimeout_metaAssert <=1'h0;
            end 
          else 
            begin 
              PlusArgTimeout_metaAssert <=PlusArgTimeout_metaAssert|PlusArgTimeout_or0;
            end 
       end
  
endmodule
 
module OptimizationBarrier (
  input [19:0] io_x_ppn,
  input io_x_u,
  input io_x_ae,
  input io_x_sw,
  input io_x_sx,
  input io_x_sr,
  input io_x_pw,
  input io_x_px,
  input io_x_pr,
  input io_x_ppp,
  input io_x_pal,
  input io_x_paa,
  input io_x_eff,
  input io_x_c,
  output [19:0] io_y_ppn,
  output io_y_u,
  output io_y_ae,
  output io_y_sw,
  output io_y_sx,
  output io_y_sr,
  output io_y_pw,
  output io_y_px,
  output io_y_pr,
  output io_y_ppp,
  output io_y_pal,
  output io_y_paa,
  output io_y_eff,
  output io_y_c,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [29:0] OptimizationBarrier_covSum ;  
  assign io_y_ppn=io_x_ppn; 
  assign io_y_u=io_x_u; 
  assign io_y_ae=io_x_ae; 
  assign io_y_sw=io_x_sw; 
  assign io_y_sx=io_x_sx; 
  assign io_y_sr=io_x_sr; 
  assign io_y_pw=io_x_pw; 
  assign io_y_px=io_x_px; 
  assign io_y_pr=io_x_pr; 
  assign io_y_ppp=io_x_ppp; 
  assign io_y_pal=io_x_pal; 
  assign io_y_paa=io_x_paa; 
  assign io_y_eff=io_x_eff; 
  assign io_y_c=io_x_c; 
  assign OptimizationBarrier_covSum=30'h0; 
  assign io_covSum=OptimizationBarrier_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module PMPChecker (
  input [1:0] io_prv,
  input io_pmp_0_cfg_l,
  input [1:0] io_pmp_0_cfg_a,
  input io_pmp_0_cfg_x,
  input io_pmp_0_cfg_w,
  input io_pmp_0_cfg_r,
  input [29:0] io_pmp_0_addr,
  input [31:0] io_pmp_0_mask,
  input io_pmp_1_cfg_l,
  input [1:0] io_pmp_1_cfg_a,
  input io_pmp_1_cfg_x,
  input io_pmp_1_cfg_w,
  input io_pmp_1_cfg_r,
  input [29:0] io_pmp_1_addr,
  input [31:0] io_pmp_1_mask,
  input io_pmp_2_cfg_l,
  input [1:0] io_pmp_2_cfg_a,
  input io_pmp_2_cfg_x,
  input io_pmp_2_cfg_w,
  input io_pmp_2_cfg_r,
  input [29:0] io_pmp_2_addr,
  input [31:0] io_pmp_2_mask,
  input io_pmp_3_cfg_l,
  input [1:0] io_pmp_3_cfg_a,
  input io_pmp_3_cfg_x,
  input io_pmp_3_cfg_w,
  input io_pmp_3_cfg_r,
  input [29:0] io_pmp_3_addr,
  input [31:0] io_pmp_3_mask,
  input io_pmp_4_cfg_l,
  input [1:0] io_pmp_4_cfg_a,
  input io_pmp_4_cfg_x,
  input io_pmp_4_cfg_w,
  input io_pmp_4_cfg_r,
  input [29:0] io_pmp_4_addr,
  input [31:0] io_pmp_4_mask,
  input io_pmp_5_cfg_l,
  input [1:0] io_pmp_5_cfg_a,
  input io_pmp_5_cfg_x,
  input io_pmp_5_cfg_w,
  input io_pmp_5_cfg_r,
  input [29:0] io_pmp_5_addr,
  input [31:0] io_pmp_5_mask,
  input io_pmp_6_cfg_l,
  input [1:0] io_pmp_6_cfg_a,
  input io_pmp_6_cfg_x,
  input io_pmp_6_cfg_w,
  input io_pmp_6_cfg_r,
  input [29:0] io_pmp_6_addr,
  input [31:0] io_pmp_6_mask,
  input io_pmp_7_cfg_l,
  input [1:0] io_pmp_7_cfg_a,
  input io_pmp_7_cfg_x,
  input io_pmp_7_cfg_w,
  input io_pmp_7_cfg_r,
  input [29:0] io_pmp_7_addr,
  input [31:0] io_pmp_7_mask,
  input [31:0] io_addr,
  input [1:0] io_size,
  output io_r,
  output io_w,
  output io_x,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire default_ ;  
   wire [5:0] _res_hit_lsbMask_T_1 ;  
   wire [31:0] _GEN_0 ;  
   wire [31:0] res_hit_lsbMask ;  
   wire [31:0] _res_hit_msbMatch_T_1 ;  
   wire [31:0] _res_hit_msbMatch_T_3 ;  
   wire [28:0] _res_hit_msbMatch_T_5 ;  
   wire [28:0] _res_hit_msbMatch_T_7 ;  
   wire [28:0] _res_hit_msbMatch_T_9 ;  
   wire res_hit_msbMatch ;  
   wire [2:0] _res_hit_lsbMatch_T_5 ;  
   wire [2:0] _res_hit_lsbMatch_T_7 ;  
   wire [2:0] _res_hit_lsbMatch_T_9 ;  
   wire res_hit_lsbMatch ;  
   wire _res_hit_T_1 ;  
   wire [31:0] _res_hit_msbsLess_T_1 ;  
   wire [31:0] _res_hit_msbsLess_T_3 ;  
   wire [28:0] _res_hit_msbsLess_T_5 ;  
   wire res_hit_msbsLess ;  
   wire [28:0] _res_hit_msbsEqual_T_6 ;  
   wire res_hit_msbsEqual ;  
   wire [2:0] _res_hit_lsbsLess_T_1 ;  
   wire [2:0] _res_hit_lsbsLess_T_6 ;  
   wire res_hit_lsbsLess ;  
   wire _res_hit_T_7 ;  
   wire _res_hit_T_8 ;  
   wire res_hit_msbsLess_1 ;  
   wire res_hit_msbsEqual_1 ;  
   wire res_hit_lsbsLess_1 ;  
   wire _res_hit_T_10 ;  
   wire _res_hit_T_11 ;  
   wire _res_hit_T_12 ;  
   wire _res_hit_T_13 ;  
   wire res_hit ;  
   wire res_ignore ;  
   wire [2:0] _res_aligned_straddlesLowerBound_T_15 ;  
   wire _res_aligned_straddlesLowerBound_T_16 ;  
   wire res_aligned_straddlesLowerBound ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_15 ;  
   wire _res_aligned_straddlesUpperBound_T_16 ;  
   wire res_aligned_straddlesUpperBound ;  
   wire _res_aligned_rangeAligned_T ;  
   wire res_aligned_rangeAligned ;  
   wire [2:0] _res_aligned_pow2Aligned_T_2 ;  
   wire res_aligned_pow2Aligned ;  
   wire res_aligned ;  
   wire _res_cur_cfg_r_T ;  
   wire res_cur_cfg_r ;  
   wire _res_cur_cfg_w_T ;  
   wire res_cur_cfg_w ;  
   wire _res_cur_cfg_x_T ;  
   wire res_cur_cfg_x ;  
   wire _res_T_44_cfg_x ;  
   wire _res_T_44_cfg_w ;  
   wire _res_T_44_cfg_r ;  
   wire [31:0] res_hit_lsbMask_1 ;  
   wire [28:0] _res_hit_msbMatch_T_19 ;  
   wire res_hit_msbMatch_1 ;  
   wire [2:0] _res_hit_lsbMatch_T_17 ;  
   wire [2:0] _res_hit_lsbMatch_T_19 ;  
   wire res_hit_lsbMatch_1 ;  
   wire _res_hit_T_15 ;  
   wire [31:0] _res_hit_msbsLess_T_13 ;  
   wire [31:0] _res_hit_msbsLess_T_15 ;  
   wire [28:0] _res_hit_msbsLess_T_17 ;  
   wire res_hit_msbsLess_2 ;  
   wire [28:0] _res_hit_msbsEqual_T_20 ;  
   wire res_hit_msbsEqual_2 ;  
   wire [2:0] _res_hit_lsbsLess_T_20 ;  
   wire res_hit_lsbsLess_2 ;  
   wire _res_hit_T_21 ;  
   wire _res_hit_T_22 ;  
   wire res_hit_lsbsLess_3 ;  
   wire _res_hit_T_24 ;  
   wire _res_hit_T_25 ;  
   wire _res_hit_T_26 ;  
   wire _res_hit_T_27 ;  
   wire res_hit_1 ;  
   wire res_ignore_1 ;  
   wire [2:0] _res_aligned_straddlesLowerBound_T_32 ;  
   wire _res_aligned_straddlesLowerBound_T_33 ;  
   wire res_aligned_straddlesLowerBound_1 ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_32 ;  
   wire _res_aligned_straddlesUpperBound_T_33 ;  
   wire res_aligned_straddlesUpperBound_1 ;  
   wire _res_aligned_rangeAligned_T_1 ;  
   wire res_aligned_rangeAligned_1 ;  
   wire [2:0] _res_aligned_pow2Aligned_T_5 ;  
   wire res_aligned_pow2Aligned_1 ;  
   wire res_aligned_1 ;  
   wire _res_cur_cfg_r_T_2 ;  
   wire res_cur_1_cfg_r ;  
   wire _res_cur_cfg_w_T_2 ;  
   wire res_cur_1_cfg_w ;  
   wire _res_cur_cfg_x_T_2 ;  
   wire res_cur_1_cfg_x ;  
   wire _res_T_89_cfg_x ;  
   wire _res_T_89_cfg_w ;  
   wire _res_T_89_cfg_r ;  
   wire [31:0] res_hit_lsbMask_2 ;  
   wire [28:0] _res_hit_msbMatch_T_29 ;  
   wire res_hit_msbMatch_2 ;  
   wire [2:0] _res_hit_lsbMatch_T_27 ;  
   wire [2:0] _res_hit_lsbMatch_T_29 ;  
   wire res_hit_lsbMatch_2 ;  
   wire _res_hit_T_29 ;  
   wire [31:0] _res_hit_msbsLess_T_25 ;  
   wire [31:0] _res_hit_msbsLess_T_27 ;  
   wire [28:0] _res_hit_msbsLess_T_29 ;  
   wire res_hit_msbsLess_4 ;  
   wire [28:0] _res_hit_msbsEqual_T_34 ;  
   wire res_hit_msbsEqual_4 ;  
   wire [2:0] _res_hit_lsbsLess_T_34 ;  
   wire res_hit_lsbsLess_4 ;  
   wire _res_hit_T_35 ;  
   wire _res_hit_T_36 ;  
   wire res_hit_lsbsLess_5 ;  
   wire _res_hit_T_38 ;  
   wire _res_hit_T_39 ;  
   wire _res_hit_T_40 ;  
   wire _res_hit_T_41 ;  
   wire res_hit_2 ;  
   wire res_ignore_2 ;  
   wire [2:0] _res_aligned_straddlesLowerBound_T_49 ;  
   wire _res_aligned_straddlesLowerBound_T_50 ;  
   wire res_aligned_straddlesLowerBound_2 ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_49 ;  
   wire _res_aligned_straddlesUpperBound_T_50 ;  
   wire res_aligned_straddlesUpperBound_2 ;  
   wire _res_aligned_rangeAligned_T_2 ;  
   wire res_aligned_rangeAligned_2 ;  
   wire [2:0] _res_aligned_pow2Aligned_T_8 ;  
   wire res_aligned_pow2Aligned_2 ;  
   wire res_aligned_2 ;  
   wire _res_cur_cfg_r_T_4 ;  
   wire res_cur_2_cfg_r ;  
   wire _res_cur_cfg_w_T_4 ;  
   wire res_cur_2_cfg_w ;  
   wire _res_cur_cfg_x_T_4 ;  
   wire res_cur_2_cfg_x ;  
   wire _res_T_134_cfg_x ;  
   wire _res_T_134_cfg_w ;  
   wire _res_T_134_cfg_r ;  
   wire [31:0] res_hit_lsbMask_3 ;  
   wire [28:0] _res_hit_msbMatch_T_39 ;  
   wire res_hit_msbMatch_3 ;  
   wire [2:0] _res_hit_lsbMatch_T_37 ;  
   wire [2:0] _res_hit_lsbMatch_T_39 ;  
   wire res_hit_lsbMatch_3 ;  
   wire _res_hit_T_43 ;  
   wire [31:0] _res_hit_msbsLess_T_37 ;  
   wire [31:0] _res_hit_msbsLess_T_39 ;  
   wire [28:0] _res_hit_msbsLess_T_41 ;  
   wire res_hit_msbsLess_6 ;  
   wire [28:0] _res_hit_msbsEqual_T_48 ;  
   wire res_hit_msbsEqual_6 ;  
   wire [2:0] _res_hit_lsbsLess_T_48 ;  
   wire res_hit_lsbsLess_6 ;  
   wire _res_hit_T_49 ;  
   wire _res_hit_T_50 ;  
   wire res_hit_lsbsLess_7 ;  
   wire _res_hit_T_52 ;  
   wire _res_hit_T_53 ;  
   wire _res_hit_T_54 ;  
   wire _res_hit_T_55 ;  
   wire res_hit_3 ;  
   wire res_ignore_3 ;  
   wire [2:0] _res_aligned_straddlesLowerBound_T_66 ;  
   wire _res_aligned_straddlesLowerBound_T_67 ;  
   wire res_aligned_straddlesLowerBound_3 ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_66 ;  
   wire _res_aligned_straddlesUpperBound_T_67 ;  
   wire res_aligned_straddlesUpperBound_3 ;  
   wire _res_aligned_rangeAligned_T_3 ;  
   wire res_aligned_rangeAligned_3 ;  
   wire [2:0] _res_aligned_pow2Aligned_T_11 ;  
   wire res_aligned_pow2Aligned_3 ;  
   wire res_aligned_3 ;  
   wire _res_cur_cfg_r_T_6 ;  
   wire res_cur_3_cfg_r ;  
   wire _res_cur_cfg_w_T_6 ;  
   wire res_cur_3_cfg_w ;  
   wire _res_cur_cfg_x_T_6 ;  
   wire res_cur_3_cfg_x ;  
   wire _res_T_179_cfg_x ;  
   wire _res_T_179_cfg_w ;  
   wire _res_T_179_cfg_r ;  
   wire [31:0] res_hit_lsbMask_4 ;  
   wire [28:0] _res_hit_msbMatch_T_49 ;  
   wire res_hit_msbMatch_4 ;  
   wire [2:0] _res_hit_lsbMatch_T_47 ;  
   wire [2:0] _res_hit_lsbMatch_T_49 ;  
   wire res_hit_lsbMatch_4 ;  
   wire _res_hit_T_57 ;  
   wire [31:0] _res_hit_msbsLess_T_49 ;  
   wire [31:0] _res_hit_msbsLess_T_51 ;  
   wire [28:0] _res_hit_msbsLess_T_53 ;  
   wire res_hit_msbsLess_8 ;  
   wire [28:0] _res_hit_msbsEqual_T_62 ;  
   wire res_hit_msbsEqual_8 ;  
   wire [2:0] _res_hit_lsbsLess_T_62 ;  
   wire res_hit_lsbsLess_8 ;  
   wire _res_hit_T_63 ;  
   wire _res_hit_T_64 ;  
   wire res_hit_lsbsLess_9 ;  
   wire _res_hit_T_66 ;  
   wire _res_hit_T_67 ;  
   wire _res_hit_T_68 ;  
   wire _res_hit_T_69 ;  
   wire res_hit_4 ;  
   wire res_ignore_4 ;  
   wire [2:0] _res_aligned_straddlesLowerBound_T_83 ;  
   wire _res_aligned_straddlesLowerBound_T_84 ;  
   wire res_aligned_straddlesLowerBound_4 ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_83 ;  
   wire _res_aligned_straddlesUpperBound_T_84 ;  
   wire res_aligned_straddlesUpperBound_4 ;  
   wire _res_aligned_rangeAligned_T_4 ;  
   wire res_aligned_rangeAligned_4 ;  
   wire [2:0] _res_aligned_pow2Aligned_T_14 ;  
   wire res_aligned_pow2Aligned_4 ;  
   wire res_aligned_4 ;  
   wire _res_cur_cfg_r_T_8 ;  
   wire res_cur_4_cfg_r ;  
   wire _res_cur_cfg_w_T_8 ;  
   wire res_cur_4_cfg_w ;  
   wire _res_cur_cfg_x_T_8 ;  
   wire res_cur_4_cfg_x ;  
   wire _res_T_224_cfg_x ;  
   wire _res_T_224_cfg_w ;  
   wire _res_T_224_cfg_r ;  
   wire [31:0] res_hit_lsbMask_5 ;  
   wire [28:0] _res_hit_msbMatch_T_59 ;  
   wire res_hit_msbMatch_5 ;  
   wire [2:0] _res_hit_lsbMatch_T_57 ;  
   wire [2:0] _res_hit_lsbMatch_T_59 ;  
   wire res_hit_lsbMatch_5 ;  
   wire _res_hit_T_71 ;  
   wire [31:0] _res_hit_msbsLess_T_61 ;  
   wire [31:0] _res_hit_msbsLess_T_63 ;  
   wire [28:0] _res_hit_msbsLess_T_65 ;  
   wire res_hit_msbsLess_10 ;  
   wire [28:0] _res_hit_msbsEqual_T_76 ;  
   wire res_hit_msbsEqual_10 ;  
   wire [2:0] _res_hit_lsbsLess_T_76 ;  
   wire res_hit_lsbsLess_10 ;  
   wire _res_hit_T_77 ;  
   wire _res_hit_T_78 ;  
   wire res_hit_lsbsLess_11 ;  
   wire _res_hit_T_80 ;  
   wire _res_hit_T_81 ;  
   wire _res_hit_T_82 ;  
   wire _res_hit_T_83 ;  
   wire res_hit_5 ;  
   wire res_ignore_5 ;  
   wire [2:0] _res_aligned_straddlesLowerBound_T_100 ;  
   wire _res_aligned_straddlesLowerBound_T_101 ;  
   wire res_aligned_straddlesLowerBound_5 ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_100 ;  
   wire _res_aligned_straddlesUpperBound_T_101 ;  
   wire res_aligned_straddlesUpperBound_5 ;  
   wire _res_aligned_rangeAligned_T_5 ;  
   wire res_aligned_rangeAligned_5 ;  
   wire [2:0] _res_aligned_pow2Aligned_T_17 ;  
   wire res_aligned_pow2Aligned_5 ;  
   wire res_aligned_5 ;  
   wire _res_cur_cfg_r_T_10 ;  
   wire res_cur_5_cfg_r ;  
   wire _res_cur_cfg_w_T_10 ;  
   wire res_cur_5_cfg_w ;  
   wire _res_cur_cfg_x_T_10 ;  
   wire res_cur_5_cfg_x ;  
   wire _res_T_269_cfg_x ;  
   wire _res_T_269_cfg_w ;  
   wire _res_T_269_cfg_r ;  
   wire [31:0] res_hit_lsbMask_6 ;  
   wire [28:0] _res_hit_msbMatch_T_69 ;  
   wire res_hit_msbMatch_6 ;  
   wire [2:0] _res_hit_lsbMatch_T_67 ;  
   wire [2:0] _res_hit_lsbMatch_T_69 ;  
   wire res_hit_lsbMatch_6 ;  
   wire _res_hit_T_85 ;  
   wire [31:0] _res_hit_msbsLess_T_73 ;  
   wire [31:0] _res_hit_msbsLess_T_75 ;  
   wire [28:0] _res_hit_msbsLess_T_77 ;  
   wire res_hit_msbsLess_12 ;  
   wire [28:0] _res_hit_msbsEqual_T_90 ;  
   wire res_hit_msbsEqual_12 ;  
   wire [2:0] _res_hit_lsbsLess_T_90 ;  
   wire res_hit_lsbsLess_12 ;  
   wire _res_hit_T_91 ;  
   wire _res_hit_T_92 ;  
   wire res_hit_lsbsLess_13 ;  
   wire _res_hit_T_94 ;  
   wire _res_hit_T_95 ;  
   wire _res_hit_T_96 ;  
   wire _res_hit_T_97 ;  
   wire res_hit_6 ;  
   wire res_ignore_6 ;  
   wire [2:0] _res_aligned_straddlesLowerBound_T_117 ;  
   wire _res_aligned_straddlesLowerBound_T_118 ;  
   wire res_aligned_straddlesLowerBound_6 ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_117 ;  
   wire _res_aligned_straddlesUpperBound_T_118 ;  
   wire res_aligned_straddlesUpperBound_6 ;  
   wire _res_aligned_rangeAligned_T_6 ;  
   wire res_aligned_rangeAligned_6 ;  
   wire [2:0] _res_aligned_pow2Aligned_T_20 ;  
   wire res_aligned_pow2Aligned_6 ;  
   wire res_aligned_6 ;  
   wire _res_cur_cfg_r_T_12 ;  
   wire res_cur_6_cfg_r ;  
   wire _res_cur_cfg_w_T_12 ;  
   wire res_cur_6_cfg_w ;  
   wire _res_cur_cfg_x_T_12 ;  
   wire res_cur_6_cfg_x ;  
   wire _res_T_314_cfg_x ;  
   wire _res_T_314_cfg_w ;  
   wire _res_T_314_cfg_r ;  
   wire [31:0] res_hit_lsbMask_7 ;  
   wire [28:0] _res_hit_msbMatch_T_79 ;  
   wire res_hit_msbMatch_7 ;  
   wire [2:0] _res_hit_lsbMatch_T_77 ;  
   wire [2:0] _res_hit_lsbMatch_T_79 ;  
   wire res_hit_lsbMatch_7 ;  
   wire _res_hit_T_99 ;  
   wire res_hit_lsbsLess_15 ;  
   wire _res_hit_T_108 ;  
   wire _res_hit_T_109 ;  
   wire _res_hit_T_111 ;  
   wire res_hit_7 ;  
   wire res_ignore_7 ;  
   wire [2:0] _res_aligned_straddlesUpperBound_T_134 ;  
   wire _res_aligned_straddlesUpperBound_T_135 ;  
   wire res_aligned_straddlesUpperBound_7 ;  
   wire res_aligned_rangeAligned_7 ;  
   wire [2:0] _res_aligned_pow2Aligned_T_23 ;  
   wire res_aligned_pow2Aligned_7 ;  
   wire res_aligned_7 ;  
   wire _res_cur_cfg_r_T_14 ;  
   wire res_cur_7_cfg_r ;  
   wire _res_cur_cfg_w_T_14 ;  
   wire res_cur_7_cfg_w ;  
   wire _res_cur_cfg_x_T_14 ;  
   wire res_cur_7_cfg_x ;  
   wire [29:0] PMPChecker_covSum ;  
  assign default_=io_prv>2'h1; 
  assign _res_hit_lsbMask_T_1=6'h7<<io_size; 
  assign _GEN_0={29'b0,~_res_hit_lsbMask_T_1[2:0]}; 
  assign res_hit_lsbMask=io_pmp_7_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_1={io_pmp_7_addr,2'h0}; 
  assign _res_hit_msbMatch_T_3=~_res_hit_msbMatch_T_1|32'h3; 
  assign _res_hit_msbMatch_T_5=~_res_hit_msbMatch_T_3[31:3]; 
  assign _res_hit_msbMatch_T_7=io_addr[31:3]^_res_hit_msbMatch_T_5; 
  assign _res_hit_msbMatch_T_9=_res_hit_msbMatch_T_7&~io_pmp_7_mask[31:3]; 
  assign res_hit_msbMatch=_res_hit_msbMatch_T_9==29'h0; 
  assign _res_hit_lsbMatch_T_5=~_res_hit_msbMatch_T_3[2:0]; 
  assign _res_hit_lsbMatch_T_7=io_addr[2:0]^_res_hit_lsbMatch_T_5; 
  assign _res_hit_lsbMatch_T_9=_res_hit_lsbMatch_T_7&~res_hit_lsbMask[2:0]; 
  assign res_hit_lsbMatch=_res_hit_lsbMatch_T_9==3'h0; 
  assign _res_hit_T_1=res_hit_msbMatch&res_hit_lsbMatch; 
  assign _res_hit_msbsLess_T_1={io_pmp_6_addr,2'h0}; 
  assign _res_hit_msbsLess_T_3=~_res_hit_msbsLess_T_1|32'h3; 
  assign _res_hit_msbsLess_T_5=~_res_hit_msbsLess_T_3[31:3]; 
  assign res_hit_msbsLess=io_addr[31:3]<_res_hit_msbsLess_T_5; 
  assign _res_hit_msbsEqual_T_6=io_addr[31:3]^_res_hit_msbsLess_T_5; 
  assign res_hit_msbsEqual=_res_hit_msbsEqual_T_6==29'h0; 
  assign _res_hit_lsbsLess_T_1=io_addr[2:0]|~_res_hit_lsbMask_T_1[2:0]; 
  assign _res_hit_lsbsLess_T_6=~_res_hit_msbsLess_T_3[2:0]; 
  assign res_hit_lsbsLess=_res_hit_lsbsLess_T_1<_res_hit_lsbsLess_T_6; 
  assign _res_hit_T_7=res_hit_msbsEqual&res_hit_lsbsLess; 
  assign _res_hit_T_8=res_hit_msbsLess|_res_hit_T_7; 
  assign res_hit_msbsLess_1=io_addr[31:3]<_res_hit_msbMatch_T_5; 
  assign res_hit_msbsEqual_1=_res_hit_msbMatch_T_7==29'h0; 
  assign res_hit_lsbsLess_1=io_addr[2:0]<_res_hit_lsbMatch_T_5; 
  assign _res_hit_T_10=res_hit_msbsEqual_1&res_hit_lsbsLess_1; 
  assign _res_hit_T_11=res_hit_msbsLess_1|_res_hit_T_10; 
  assign _res_hit_T_12=~_res_hit_T_8&_res_hit_T_11; 
  assign _res_hit_T_13=io_pmp_7_cfg_a[0]&_res_hit_T_12; 
  assign res_hit=io_pmp_7_cfg_a[1] ? _res_hit_T_1:_res_hit_T_13; 
  assign res_ignore=default_&~io_pmp_7_cfg_l; 
  assign _res_aligned_straddlesLowerBound_T_15=_res_hit_lsbsLess_T_6&~io_addr[2:0]; 
  assign _res_aligned_straddlesLowerBound_T_16=_res_aligned_straddlesLowerBound_T_15!=3'h0; 
  assign res_aligned_straddlesLowerBound=res_hit_msbsEqual&_res_aligned_straddlesLowerBound_T_16; 
  assign _res_aligned_straddlesUpperBound_T_15=_res_hit_lsbMatch_T_5&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_16=_res_aligned_straddlesUpperBound_T_15!=3'h0; 
  assign res_aligned_straddlesUpperBound=res_hit_msbsEqual_1&_res_aligned_straddlesUpperBound_T_16; 
  assign _res_aligned_rangeAligned_T=res_aligned_straddlesLowerBound|res_aligned_straddlesUpperBound; 
  assign res_aligned_rangeAligned=~_res_aligned_rangeAligned_T; 
  assign _res_aligned_pow2Aligned_T_2=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_7_mask[2:0]; 
  assign res_aligned_pow2Aligned=_res_aligned_pow2Aligned_T_2==3'h0; 
  assign res_aligned=io_pmp_7_cfg_a[1] ? res_aligned_pow2Aligned:res_aligned_rangeAligned; 
  assign _res_cur_cfg_r_T=io_pmp_7_cfg_r|res_ignore; 
  assign res_cur_cfg_r=res_aligned&_res_cur_cfg_r_T; 
  assign _res_cur_cfg_w_T=io_pmp_7_cfg_w|res_ignore; 
  assign res_cur_cfg_w=res_aligned&_res_cur_cfg_w_T; 
  assign _res_cur_cfg_x_T=io_pmp_7_cfg_x|res_ignore; 
  assign res_cur_cfg_x=res_aligned&_res_cur_cfg_x_T; 
  assign _res_T_44_cfg_x=res_hit ? res_cur_cfg_x:default_; 
  assign _res_T_44_cfg_w=res_hit ? res_cur_cfg_w:default_; 
  assign _res_T_44_cfg_r=res_hit ? res_cur_cfg_r:default_; 
  assign res_hit_lsbMask_1=io_pmp_6_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_19=_res_hit_msbsEqual_T_6&~io_pmp_6_mask[31:3]; 
  assign res_hit_msbMatch_1=_res_hit_msbMatch_T_19==29'h0; 
  assign _res_hit_lsbMatch_T_17=io_addr[2:0]^_res_hit_lsbsLess_T_6; 
  assign _res_hit_lsbMatch_T_19=_res_hit_lsbMatch_T_17&~res_hit_lsbMask_1[2:0]; 
  assign res_hit_lsbMatch_1=_res_hit_lsbMatch_T_19==3'h0; 
  assign _res_hit_T_15=res_hit_msbMatch_1&res_hit_lsbMatch_1; 
  assign _res_hit_msbsLess_T_13={io_pmp_5_addr,2'h0}; 
  assign _res_hit_msbsLess_T_15=~_res_hit_msbsLess_T_13|32'h3; 
  assign _res_hit_msbsLess_T_17=~_res_hit_msbsLess_T_15[31:3]; 
  assign res_hit_msbsLess_2=io_addr[31:3]<_res_hit_msbsLess_T_17; 
  assign _res_hit_msbsEqual_T_20=io_addr[31:3]^_res_hit_msbsLess_T_17; 
  assign res_hit_msbsEqual_2=_res_hit_msbsEqual_T_20==29'h0; 
  assign _res_hit_lsbsLess_T_20=~_res_hit_msbsLess_T_15[2:0]; 
  assign res_hit_lsbsLess_2=_res_hit_lsbsLess_T_1<_res_hit_lsbsLess_T_20; 
  assign _res_hit_T_21=res_hit_msbsEqual_2&res_hit_lsbsLess_2; 
  assign _res_hit_T_22=res_hit_msbsLess_2|_res_hit_T_21; 
  assign res_hit_lsbsLess_3=io_addr[2:0]<_res_hit_lsbsLess_T_6; 
  assign _res_hit_T_24=res_hit_msbsEqual&res_hit_lsbsLess_3; 
  assign _res_hit_T_25=res_hit_msbsLess|_res_hit_T_24; 
  assign _res_hit_T_26=~_res_hit_T_22&_res_hit_T_25; 
  assign _res_hit_T_27=io_pmp_6_cfg_a[0]&_res_hit_T_26; 
  assign res_hit_1=io_pmp_6_cfg_a[1] ? _res_hit_T_15:_res_hit_T_27; 
  assign res_ignore_1=default_&~io_pmp_6_cfg_l; 
  assign _res_aligned_straddlesLowerBound_T_32=_res_hit_lsbsLess_T_20&~io_addr[2:0]; 
  assign _res_aligned_straddlesLowerBound_T_33=_res_aligned_straddlesLowerBound_T_32!=3'h0; 
  assign res_aligned_straddlesLowerBound_1=res_hit_msbsEqual_2&_res_aligned_straddlesLowerBound_T_33; 
  assign _res_aligned_straddlesUpperBound_T_32=_res_hit_lsbsLess_T_6&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_33=_res_aligned_straddlesUpperBound_T_32!=3'h0; 
  assign res_aligned_straddlesUpperBound_1=res_hit_msbsEqual&_res_aligned_straddlesUpperBound_T_33; 
  assign _res_aligned_rangeAligned_T_1=res_aligned_straddlesLowerBound_1|res_aligned_straddlesUpperBound_1; 
  assign res_aligned_rangeAligned_1=~_res_aligned_rangeAligned_T_1; 
  assign _res_aligned_pow2Aligned_T_5=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_6_mask[2:0]; 
  assign res_aligned_pow2Aligned_1=_res_aligned_pow2Aligned_T_5==3'h0; 
  assign res_aligned_1=io_pmp_6_cfg_a[1] ? res_aligned_pow2Aligned_1:res_aligned_rangeAligned_1; 
  assign _res_cur_cfg_r_T_2=io_pmp_6_cfg_r|res_ignore_1; 
  assign res_cur_1_cfg_r=res_aligned_1&_res_cur_cfg_r_T_2; 
  assign _res_cur_cfg_w_T_2=io_pmp_6_cfg_w|res_ignore_1; 
  assign res_cur_1_cfg_w=res_aligned_1&_res_cur_cfg_w_T_2; 
  assign _res_cur_cfg_x_T_2=io_pmp_6_cfg_x|res_ignore_1; 
  assign res_cur_1_cfg_x=res_aligned_1&_res_cur_cfg_x_T_2; 
  assign _res_T_89_cfg_x=res_hit_1 ? res_cur_1_cfg_x:_res_T_44_cfg_x; 
  assign _res_T_89_cfg_w=res_hit_1 ? res_cur_1_cfg_w:_res_T_44_cfg_w; 
  assign _res_T_89_cfg_r=res_hit_1 ? res_cur_1_cfg_r:_res_T_44_cfg_r; 
  assign res_hit_lsbMask_2=io_pmp_5_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_29=_res_hit_msbsEqual_T_20&~io_pmp_5_mask[31:3]; 
  assign res_hit_msbMatch_2=_res_hit_msbMatch_T_29==29'h0; 
  assign _res_hit_lsbMatch_T_27=io_addr[2:0]^_res_hit_lsbsLess_T_20; 
  assign _res_hit_lsbMatch_T_29=_res_hit_lsbMatch_T_27&~res_hit_lsbMask_2[2:0]; 
  assign res_hit_lsbMatch_2=_res_hit_lsbMatch_T_29==3'h0; 
  assign _res_hit_T_29=res_hit_msbMatch_2&res_hit_lsbMatch_2; 
  assign _res_hit_msbsLess_T_25={io_pmp_4_addr,2'h0}; 
  assign _res_hit_msbsLess_T_27=~_res_hit_msbsLess_T_25|32'h3; 
  assign _res_hit_msbsLess_T_29=~_res_hit_msbsLess_T_27[31:3]; 
  assign res_hit_msbsLess_4=io_addr[31:3]<_res_hit_msbsLess_T_29; 
  assign _res_hit_msbsEqual_T_34=io_addr[31:3]^_res_hit_msbsLess_T_29; 
  assign res_hit_msbsEqual_4=_res_hit_msbsEqual_T_34==29'h0; 
  assign _res_hit_lsbsLess_T_34=~_res_hit_msbsLess_T_27[2:0]; 
  assign res_hit_lsbsLess_4=_res_hit_lsbsLess_T_1<_res_hit_lsbsLess_T_34; 
  assign _res_hit_T_35=res_hit_msbsEqual_4&res_hit_lsbsLess_4; 
  assign _res_hit_T_36=res_hit_msbsLess_4|_res_hit_T_35; 
  assign res_hit_lsbsLess_5=io_addr[2:0]<_res_hit_lsbsLess_T_20; 
  assign _res_hit_T_38=res_hit_msbsEqual_2&res_hit_lsbsLess_5; 
  assign _res_hit_T_39=res_hit_msbsLess_2|_res_hit_T_38; 
  assign _res_hit_T_40=~_res_hit_T_36&_res_hit_T_39; 
  assign _res_hit_T_41=io_pmp_5_cfg_a[0]&_res_hit_T_40; 
  assign res_hit_2=io_pmp_5_cfg_a[1] ? _res_hit_T_29:_res_hit_T_41; 
  assign res_ignore_2=default_&~io_pmp_5_cfg_l; 
  assign _res_aligned_straddlesLowerBound_T_49=_res_hit_lsbsLess_T_34&~io_addr[2:0]; 
  assign _res_aligned_straddlesLowerBound_T_50=_res_aligned_straddlesLowerBound_T_49!=3'h0; 
  assign res_aligned_straddlesLowerBound_2=res_hit_msbsEqual_4&_res_aligned_straddlesLowerBound_T_50; 
  assign _res_aligned_straddlesUpperBound_T_49=_res_hit_lsbsLess_T_20&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_50=_res_aligned_straddlesUpperBound_T_49!=3'h0; 
  assign res_aligned_straddlesUpperBound_2=res_hit_msbsEqual_2&_res_aligned_straddlesUpperBound_T_50; 
  assign _res_aligned_rangeAligned_T_2=res_aligned_straddlesLowerBound_2|res_aligned_straddlesUpperBound_2; 
  assign res_aligned_rangeAligned_2=~_res_aligned_rangeAligned_T_2; 
  assign _res_aligned_pow2Aligned_T_8=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_5_mask[2:0]; 
  assign res_aligned_pow2Aligned_2=_res_aligned_pow2Aligned_T_8==3'h0; 
  assign res_aligned_2=io_pmp_5_cfg_a[1] ? res_aligned_pow2Aligned_2:res_aligned_rangeAligned_2; 
  assign _res_cur_cfg_r_T_4=io_pmp_5_cfg_r|res_ignore_2; 
  assign res_cur_2_cfg_r=res_aligned_2&_res_cur_cfg_r_T_4; 
  assign _res_cur_cfg_w_T_4=io_pmp_5_cfg_w|res_ignore_2; 
  assign res_cur_2_cfg_w=res_aligned_2&_res_cur_cfg_w_T_4; 
  assign _res_cur_cfg_x_T_4=io_pmp_5_cfg_x|res_ignore_2; 
  assign res_cur_2_cfg_x=res_aligned_2&_res_cur_cfg_x_T_4; 
  assign _res_T_134_cfg_x=res_hit_2 ? res_cur_2_cfg_x:_res_T_89_cfg_x; 
  assign _res_T_134_cfg_w=res_hit_2 ? res_cur_2_cfg_w:_res_T_89_cfg_w; 
  assign _res_T_134_cfg_r=res_hit_2 ? res_cur_2_cfg_r:_res_T_89_cfg_r; 
  assign res_hit_lsbMask_3=io_pmp_4_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_39=_res_hit_msbsEqual_T_34&~io_pmp_4_mask[31:3]; 
  assign res_hit_msbMatch_3=_res_hit_msbMatch_T_39==29'h0; 
  assign _res_hit_lsbMatch_T_37=io_addr[2:0]^_res_hit_lsbsLess_T_34; 
  assign _res_hit_lsbMatch_T_39=_res_hit_lsbMatch_T_37&~res_hit_lsbMask_3[2:0]; 
  assign res_hit_lsbMatch_3=_res_hit_lsbMatch_T_39==3'h0; 
  assign _res_hit_T_43=res_hit_msbMatch_3&res_hit_lsbMatch_3; 
  assign _res_hit_msbsLess_T_37={io_pmp_3_addr,2'h0}; 
  assign _res_hit_msbsLess_T_39=~_res_hit_msbsLess_T_37|32'h3; 
  assign _res_hit_msbsLess_T_41=~_res_hit_msbsLess_T_39[31:3]; 
  assign res_hit_msbsLess_6=io_addr[31:3]<_res_hit_msbsLess_T_41; 
  assign _res_hit_msbsEqual_T_48=io_addr[31:3]^_res_hit_msbsLess_T_41; 
  assign res_hit_msbsEqual_6=_res_hit_msbsEqual_T_48==29'h0; 
  assign _res_hit_lsbsLess_T_48=~_res_hit_msbsLess_T_39[2:0]; 
  assign res_hit_lsbsLess_6=_res_hit_lsbsLess_T_1<_res_hit_lsbsLess_T_48; 
  assign _res_hit_T_49=res_hit_msbsEqual_6&res_hit_lsbsLess_6; 
  assign _res_hit_T_50=res_hit_msbsLess_6|_res_hit_T_49; 
  assign res_hit_lsbsLess_7=io_addr[2:0]<_res_hit_lsbsLess_T_34; 
  assign _res_hit_T_52=res_hit_msbsEqual_4&res_hit_lsbsLess_7; 
  assign _res_hit_T_53=res_hit_msbsLess_4|_res_hit_T_52; 
  assign _res_hit_T_54=~_res_hit_T_50&_res_hit_T_53; 
  assign _res_hit_T_55=io_pmp_4_cfg_a[0]&_res_hit_T_54; 
  assign res_hit_3=io_pmp_4_cfg_a[1] ? _res_hit_T_43:_res_hit_T_55; 
  assign res_ignore_3=default_&~io_pmp_4_cfg_l; 
  assign _res_aligned_straddlesLowerBound_T_66=_res_hit_lsbsLess_T_48&~io_addr[2:0]; 
  assign _res_aligned_straddlesLowerBound_T_67=_res_aligned_straddlesLowerBound_T_66!=3'h0; 
  assign res_aligned_straddlesLowerBound_3=res_hit_msbsEqual_6&_res_aligned_straddlesLowerBound_T_67; 
  assign _res_aligned_straddlesUpperBound_T_66=_res_hit_lsbsLess_T_34&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_67=_res_aligned_straddlesUpperBound_T_66!=3'h0; 
  assign res_aligned_straddlesUpperBound_3=res_hit_msbsEqual_4&_res_aligned_straddlesUpperBound_T_67; 
  assign _res_aligned_rangeAligned_T_3=res_aligned_straddlesLowerBound_3|res_aligned_straddlesUpperBound_3; 
  assign res_aligned_rangeAligned_3=~_res_aligned_rangeAligned_T_3; 
  assign _res_aligned_pow2Aligned_T_11=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_4_mask[2:0]; 
  assign res_aligned_pow2Aligned_3=_res_aligned_pow2Aligned_T_11==3'h0; 
  assign res_aligned_3=io_pmp_4_cfg_a[1] ? res_aligned_pow2Aligned_3:res_aligned_rangeAligned_3; 
  assign _res_cur_cfg_r_T_6=io_pmp_4_cfg_r|res_ignore_3; 
  assign res_cur_3_cfg_r=res_aligned_3&_res_cur_cfg_r_T_6; 
  assign _res_cur_cfg_w_T_6=io_pmp_4_cfg_w|res_ignore_3; 
  assign res_cur_3_cfg_w=res_aligned_3&_res_cur_cfg_w_T_6; 
  assign _res_cur_cfg_x_T_6=io_pmp_4_cfg_x|res_ignore_3; 
  assign res_cur_3_cfg_x=res_aligned_3&_res_cur_cfg_x_T_6; 
  assign _res_T_179_cfg_x=res_hit_3 ? res_cur_3_cfg_x:_res_T_134_cfg_x; 
  assign _res_T_179_cfg_w=res_hit_3 ? res_cur_3_cfg_w:_res_T_134_cfg_w; 
  assign _res_T_179_cfg_r=res_hit_3 ? res_cur_3_cfg_r:_res_T_134_cfg_r; 
  assign res_hit_lsbMask_4=io_pmp_3_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_49=_res_hit_msbsEqual_T_48&~io_pmp_3_mask[31:3]; 
  assign res_hit_msbMatch_4=_res_hit_msbMatch_T_49==29'h0; 
  assign _res_hit_lsbMatch_T_47=io_addr[2:0]^_res_hit_lsbsLess_T_48; 
  assign _res_hit_lsbMatch_T_49=_res_hit_lsbMatch_T_47&~res_hit_lsbMask_4[2:0]; 
  assign res_hit_lsbMatch_4=_res_hit_lsbMatch_T_49==3'h0; 
  assign _res_hit_T_57=res_hit_msbMatch_4&res_hit_lsbMatch_4; 
  assign _res_hit_msbsLess_T_49={io_pmp_2_addr,2'h0}; 
  assign _res_hit_msbsLess_T_51=~_res_hit_msbsLess_T_49|32'h3; 
  assign _res_hit_msbsLess_T_53=~_res_hit_msbsLess_T_51[31:3]; 
  assign res_hit_msbsLess_8=io_addr[31:3]<_res_hit_msbsLess_T_53; 
  assign _res_hit_msbsEqual_T_62=io_addr[31:3]^_res_hit_msbsLess_T_53; 
  assign res_hit_msbsEqual_8=_res_hit_msbsEqual_T_62==29'h0; 
  assign _res_hit_lsbsLess_T_62=~_res_hit_msbsLess_T_51[2:0]; 
  assign res_hit_lsbsLess_8=_res_hit_lsbsLess_T_1<_res_hit_lsbsLess_T_62; 
  assign _res_hit_T_63=res_hit_msbsEqual_8&res_hit_lsbsLess_8; 
  assign _res_hit_T_64=res_hit_msbsLess_8|_res_hit_T_63; 
  assign res_hit_lsbsLess_9=io_addr[2:0]<_res_hit_lsbsLess_T_48; 
  assign _res_hit_T_66=res_hit_msbsEqual_6&res_hit_lsbsLess_9; 
  assign _res_hit_T_67=res_hit_msbsLess_6|_res_hit_T_66; 
  assign _res_hit_T_68=~_res_hit_T_64&_res_hit_T_67; 
  assign _res_hit_T_69=io_pmp_3_cfg_a[0]&_res_hit_T_68; 
  assign res_hit_4=io_pmp_3_cfg_a[1] ? _res_hit_T_57:_res_hit_T_69; 
  assign res_ignore_4=default_&~io_pmp_3_cfg_l; 
  assign _res_aligned_straddlesLowerBound_T_83=_res_hit_lsbsLess_T_62&~io_addr[2:0]; 
  assign _res_aligned_straddlesLowerBound_T_84=_res_aligned_straddlesLowerBound_T_83!=3'h0; 
  assign res_aligned_straddlesLowerBound_4=res_hit_msbsEqual_8&_res_aligned_straddlesLowerBound_T_84; 
  assign _res_aligned_straddlesUpperBound_T_83=_res_hit_lsbsLess_T_48&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_84=_res_aligned_straddlesUpperBound_T_83!=3'h0; 
  assign res_aligned_straddlesUpperBound_4=res_hit_msbsEqual_6&_res_aligned_straddlesUpperBound_T_84; 
  assign _res_aligned_rangeAligned_T_4=res_aligned_straddlesLowerBound_4|res_aligned_straddlesUpperBound_4; 
  assign res_aligned_rangeAligned_4=~_res_aligned_rangeAligned_T_4; 
  assign _res_aligned_pow2Aligned_T_14=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_3_mask[2:0]; 
  assign res_aligned_pow2Aligned_4=_res_aligned_pow2Aligned_T_14==3'h0; 
  assign res_aligned_4=io_pmp_3_cfg_a[1] ? res_aligned_pow2Aligned_4:res_aligned_rangeAligned_4; 
  assign _res_cur_cfg_r_T_8=io_pmp_3_cfg_r|res_ignore_4; 
  assign res_cur_4_cfg_r=res_aligned_4&_res_cur_cfg_r_T_8; 
  assign _res_cur_cfg_w_T_8=io_pmp_3_cfg_w|res_ignore_4; 
  assign res_cur_4_cfg_w=res_aligned_4&_res_cur_cfg_w_T_8; 
  assign _res_cur_cfg_x_T_8=io_pmp_3_cfg_x|res_ignore_4; 
  assign res_cur_4_cfg_x=res_aligned_4&_res_cur_cfg_x_T_8; 
  assign _res_T_224_cfg_x=res_hit_4 ? res_cur_4_cfg_x:_res_T_179_cfg_x; 
  assign _res_T_224_cfg_w=res_hit_4 ? res_cur_4_cfg_w:_res_T_179_cfg_w; 
  assign _res_T_224_cfg_r=res_hit_4 ? res_cur_4_cfg_r:_res_T_179_cfg_r; 
  assign res_hit_lsbMask_5=io_pmp_2_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_59=_res_hit_msbsEqual_T_62&~io_pmp_2_mask[31:3]; 
  assign res_hit_msbMatch_5=_res_hit_msbMatch_T_59==29'h0; 
  assign _res_hit_lsbMatch_T_57=io_addr[2:0]^_res_hit_lsbsLess_T_62; 
  assign _res_hit_lsbMatch_T_59=_res_hit_lsbMatch_T_57&~res_hit_lsbMask_5[2:0]; 
  assign res_hit_lsbMatch_5=_res_hit_lsbMatch_T_59==3'h0; 
  assign _res_hit_T_71=res_hit_msbMatch_5&res_hit_lsbMatch_5; 
  assign _res_hit_msbsLess_T_61={io_pmp_1_addr,2'h0}; 
  assign _res_hit_msbsLess_T_63=~_res_hit_msbsLess_T_61|32'h3; 
  assign _res_hit_msbsLess_T_65=~_res_hit_msbsLess_T_63[31:3]; 
  assign res_hit_msbsLess_10=io_addr[31:3]<_res_hit_msbsLess_T_65; 
  assign _res_hit_msbsEqual_T_76=io_addr[31:3]^_res_hit_msbsLess_T_65; 
  assign res_hit_msbsEqual_10=_res_hit_msbsEqual_T_76==29'h0; 
  assign _res_hit_lsbsLess_T_76=~_res_hit_msbsLess_T_63[2:0]; 
  assign res_hit_lsbsLess_10=_res_hit_lsbsLess_T_1<_res_hit_lsbsLess_T_76; 
  assign _res_hit_T_77=res_hit_msbsEqual_10&res_hit_lsbsLess_10; 
  assign _res_hit_T_78=res_hit_msbsLess_10|_res_hit_T_77; 
  assign res_hit_lsbsLess_11=io_addr[2:0]<_res_hit_lsbsLess_T_62; 
  assign _res_hit_T_80=res_hit_msbsEqual_8&res_hit_lsbsLess_11; 
  assign _res_hit_T_81=res_hit_msbsLess_8|_res_hit_T_80; 
  assign _res_hit_T_82=~_res_hit_T_78&_res_hit_T_81; 
  assign _res_hit_T_83=io_pmp_2_cfg_a[0]&_res_hit_T_82; 
  assign res_hit_5=io_pmp_2_cfg_a[1] ? _res_hit_T_71:_res_hit_T_83; 
  assign res_ignore_5=default_&~io_pmp_2_cfg_l; 
  assign _res_aligned_straddlesLowerBound_T_100=_res_hit_lsbsLess_T_76&~io_addr[2:0]; 
  assign _res_aligned_straddlesLowerBound_T_101=_res_aligned_straddlesLowerBound_T_100!=3'h0; 
  assign res_aligned_straddlesLowerBound_5=res_hit_msbsEqual_10&_res_aligned_straddlesLowerBound_T_101; 
  assign _res_aligned_straddlesUpperBound_T_100=_res_hit_lsbsLess_T_62&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_101=_res_aligned_straddlesUpperBound_T_100!=3'h0; 
  assign res_aligned_straddlesUpperBound_5=res_hit_msbsEqual_8&_res_aligned_straddlesUpperBound_T_101; 
  assign _res_aligned_rangeAligned_T_5=res_aligned_straddlesLowerBound_5|res_aligned_straddlesUpperBound_5; 
  assign res_aligned_rangeAligned_5=~_res_aligned_rangeAligned_T_5; 
  assign _res_aligned_pow2Aligned_T_17=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_2_mask[2:0]; 
  assign res_aligned_pow2Aligned_5=_res_aligned_pow2Aligned_T_17==3'h0; 
  assign res_aligned_5=io_pmp_2_cfg_a[1] ? res_aligned_pow2Aligned_5:res_aligned_rangeAligned_5; 
  assign _res_cur_cfg_r_T_10=io_pmp_2_cfg_r|res_ignore_5; 
  assign res_cur_5_cfg_r=res_aligned_5&_res_cur_cfg_r_T_10; 
  assign _res_cur_cfg_w_T_10=io_pmp_2_cfg_w|res_ignore_5; 
  assign res_cur_5_cfg_w=res_aligned_5&_res_cur_cfg_w_T_10; 
  assign _res_cur_cfg_x_T_10=io_pmp_2_cfg_x|res_ignore_5; 
  assign res_cur_5_cfg_x=res_aligned_5&_res_cur_cfg_x_T_10; 
  assign _res_T_269_cfg_x=res_hit_5 ? res_cur_5_cfg_x:_res_T_224_cfg_x; 
  assign _res_T_269_cfg_w=res_hit_5 ? res_cur_5_cfg_w:_res_T_224_cfg_w; 
  assign _res_T_269_cfg_r=res_hit_5 ? res_cur_5_cfg_r:_res_T_224_cfg_r; 
  assign res_hit_lsbMask_6=io_pmp_1_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_69=_res_hit_msbsEqual_T_76&~io_pmp_1_mask[31:3]; 
  assign res_hit_msbMatch_6=_res_hit_msbMatch_T_69==29'h0; 
  assign _res_hit_lsbMatch_T_67=io_addr[2:0]^_res_hit_lsbsLess_T_76; 
  assign _res_hit_lsbMatch_T_69=_res_hit_lsbMatch_T_67&~res_hit_lsbMask_6[2:0]; 
  assign res_hit_lsbMatch_6=_res_hit_lsbMatch_T_69==3'h0; 
  assign _res_hit_T_85=res_hit_msbMatch_6&res_hit_lsbMatch_6; 
  assign _res_hit_msbsLess_T_73={io_pmp_0_addr,2'h0}; 
  assign _res_hit_msbsLess_T_75=~_res_hit_msbsLess_T_73|32'h3; 
  assign _res_hit_msbsLess_T_77=~_res_hit_msbsLess_T_75[31:3]; 
  assign res_hit_msbsLess_12=io_addr[31:3]<_res_hit_msbsLess_T_77; 
  assign _res_hit_msbsEqual_T_90=io_addr[31:3]^_res_hit_msbsLess_T_77; 
  assign res_hit_msbsEqual_12=_res_hit_msbsEqual_T_90==29'h0; 
  assign _res_hit_lsbsLess_T_90=~_res_hit_msbsLess_T_75[2:0]; 
  assign res_hit_lsbsLess_12=_res_hit_lsbsLess_T_1<_res_hit_lsbsLess_T_90; 
  assign _res_hit_T_91=res_hit_msbsEqual_12&res_hit_lsbsLess_12; 
  assign _res_hit_T_92=res_hit_msbsLess_12|_res_hit_T_91; 
  assign res_hit_lsbsLess_13=io_addr[2:0]<_res_hit_lsbsLess_T_76; 
  assign _res_hit_T_94=res_hit_msbsEqual_10&res_hit_lsbsLess_13; 
  assign _res_hit_T_95=res_hit_msbsLess_10|_res_hit_T_94; 
  assign _res_hit_T_96=~_res_hit_T_92&_res_hit_T_95; 
  assign _res_hit_T_97=io_pmp_1_cfg_a[0]&_res_hit_T_96; 
  assign res_hit_6=io_pmp_1_cfg_a[1] ? _res_hit_T_85:_res_hit_T_97; 
  assign res_ignore_6=default_&~io_pmp_1_cfg_l; 
  assign _res_aligned_straddlesLowerBound_T_117=_res_hit_lsbsLess_T_90&~io_addr[2:0]; 
  assign _res_aligned_straddlesLowerBound_T_118=_res_aligned_straddlesLowerBound_T_117!=3'h0; 
  assign res_aligned_straddlesLowerBound_6=res_hit_msbsEqual_12&_res_aligned_straddlesLowerBound_T_118; 
  assign _res_aligned_straddlesUpperBound_T_117=_res_hit_lsbsLess_T_76&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_118=_res_aligned_straddlesUpperBound_T_117!=3'h0; 
  assign res_aligned_straddlesUpperBound_6=res_hit_msbsEqual_10&_res_aligned_straddlesUpperBound_T_118; 
  assign _res_aligned_rangeAligned_T_6=res_aligned_straddlesLowerBound_6|res_aligned_straddlesUpperBound_6; 
  assign res_aligned_rangeAligned_6=~_res_aligned_rangeAligned_T_6; 
  assign _res_aligned_pow2Aligned_T_20=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_1_mask[2:0]; 
  assign res_aligned_pow2Aligned_6=_res_aligned_pow2Aligned_T_20==3'h0; 
  assign res_aligned_6=io_pmp_1_cfg_a[1] ? res_aligned_pow2Aligned_6:res_aligned_rangeAligned_6; 
  assign _res_cur_cfg_r_T_12=io_pmp_1_cfg_r|res_ignore_6; 
  assign res_cur_6_cfg_r=res_aligned_6&_res_cur_cfg_r_T_12; 
  assign _res_cur_cfg_w_T_12=io_pmp_1_cfg_w|res_ignore_6; 
  assign res_cur_6_cfg_w=res_aligned_6&_res_cur_cfg_w_T_12; 
  assign _res_cur_cfg_x_T_12=io_pmp_1_cfg_x|res_ignore_6; 
  assign res_cur_6_cfg_x=res_aligned_6&_res_cur_cfg_x_T_12; 
  assign _res_T_314_cfg_x=res_hit_6 ? res_cur_6_cfg_x:_res_T_269_cfg_x; 
  assign _res_T_314_cfg_w=res_hit_6 ? res_cur_6_cfg_w:_res_T_269_cfg_w; 
  assign _res_T_314_cfg_r=res_hit_6 ? res_cur_6_cfg_r:_res_T_269_cfg_r; 
  assign res_hit_lsbMask_7=io_pmp_0_mask|_GEN_0; 
  assign _res_hit_msbMatch_T_79=_res_hit_msbsEqual_T_90&~io_pmp_0_mask[31:3]; 
  assign res_hit_msbMatch_7=_res_hit_msbMatch_T_79==29'h0; 
  assign _res_hit_lsbMatch_T_77=io_addr[2:0]^_res_hit_lsbsLess_T_90; 
  assign _res_hit_lsbMatch_T_79=_res_hit_lsbMatch_T_77&~res_hit_lsbMask_7[2:0]; 
  assign res_hit_lsbMatch_7=_res_hit_lsbMatch_T_79==3'h0; 
  assign _res_hit_T_99=res_hit_msbMatch_7&res_hit_lsbMatch_7; 
  assign res_hit_lsbsLess_15=io_addr[2:0]<_res_hit_lsbsLess_T_90; 
  assign _res_hit_T_108=res_hit_msbsEqual_12&res_hit_lsbsLess_15; 
  assign _res_hit_T_109=res_hit_msbsLess_12|_res_hit_T_108; 
  assign _res_hit_T_111=io_pmp_0_cfg_a[0]&_res_hit_T_109; 
  assign res_hit_7=io_pmp_0_cfg_a[1] ? _res_hit_T_99:_res_hit_T_111; 
  assign res_ignore_7=default_&~io_pmp_0_cfg_l; 
  assign _res_aligned_straddlesUpperBound_T_134=_res_hit_lsbsLess_T_90&_res_hit_lsbsLess_T_1; 
  assign _res_aligned_straddlesUpperBound_T_135=_res_aligned_straddlesUpperBound_T_134!=3'h0; 
  assign res_aligned_straddlesUpperBound_7=res_hit_msbsEqual_12&_res_aligned_straddlesUpperBound_T_135; 
  assign res_aligned_rangeAligned_7=~res_aligned_straddlesUpperBound_7; 
  assign _res_aligned_pow2Aligned_T_23=~_res_hit_lsbMask_T_1[2:0]&~io_pmp_0_mask[2:0]; 
  assign res_aligned_pow2Aligned_7=_res_aligned_pow2Aligned_T_23==3'h0; 
  assign res_aligned_7=io_pmp_0_cfg_a[1] ? res_aligned_pow2Aligned_7:res_aligned_rangeAligned_7; 
  assign _res_cur_cfg_r_T_14=io_pmp_0_cfg_r|res_ignore_7; 
  assign res_cur_7_cfg_r=res_aligned_7&_res_cur_cfg_r_T_14; 
  assign _res_cur_cfg_w_T_14=io_pmp_0_cfg_w|res_ignore_7; 
  assign res_cur_7_cfg_w=res_aligned_7&_res_cur_cfg_w_T_14; 
  assign _res_cur_cfg_x_T_14=io_pmp_0_cfg_x|res_ignore_7; 
  assign res_cur_7_cfg_x=res_aligned_7&_res_cur_cfg_x_T_14; 
  assign io_r=res_hit_7 ? res_cur_7_cfg_r:_res_T_314_cfg_r; 
  assign io_w=res_hit_7 ? res_cur_7_cfg_w:_res_T_314_cfg_w; 
  assign io_x=res_hit_7 ? res_cur_7_cfg_x:_res_T_314_cfg_x; 
  assign PMPChecker_covSum=30'h0; 
  assign io_covSum=PMPChecker_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module PMPChecker_2 (
  input [1:0] io_prv,
  input io_pmp_0_cfg_l,
  input [1:0] io_pmp_0_cfg_a,
  input io_pmp_0_cfg_x,
  input io_pmp_0_cfg_w,
  input io_pmp_0_cfg_r,
  input [29:0] io_pmp_0_addr,
  input [31:0] io_pmp_0_mask,
  input io_pmp_1_cfg_l,
  input [1:0] io_pmp_1_cfg_a,
  input io_pmp_1_cfg_x,
  input io_pmp_1_cfg_w,
  input io_pmp_1_cfg_r,
  input [29:0] io_pmp_1_addr,
  input [31:0] io_pmp_1_mask,
  input io_pmp_2_cfg_l,
  input [1:0] io_pmp_2_cfg_a,
  input io_pmp_2_cfg_x,
  input io_pmp_2_cfg_w,
  input io_pmp_2_cfg_r,
  input [29:0] io_pmp_2_addr,
  input [31:0] io_pmp_2_mask,
  input io_pmp_3_cfg_l,
  input [1:0] io_pmp_3_cfg_a,
  input io_pmp_3_cfg_x,
  input io_pmp_3_cfg_w,
  input io_pmp_3_cfg_r,
  input [29:0] io_pmp_3_addr,
  input [31:0] io_pmp_3_mask,
  input io_pmp_4_cfg_l,
  input [1:0] io_pmp_4_cfg_a,
  input io_pmp_4_cfg_x,
  input io_pmp_4_cfg_w,
  input io_pmp_4_cfg_r,
  input [29:0] io_pmp_4_addr,
  input [31:0] io_pmp_4_mask,
  input io_pmp_5_cfg_l,
  input [1:0] io_pmp_5_cfg_a,
  input io_pmp_5_cfg_x,
  input io_pmp_5_cfg_w,
  input io_pmp_5_cfg_r,
  input [29:0] io_pmp_5_addr,
  input [31:0] io_pmp_5_mask,
  input io_pmp_6_cfg_l,
  input [1:0] io_pmp_6_cfg_a,
  input io_pmp_6_cfg_x,
  input io_pmp_6_cfg_w,
  input io_pmp_6_cfg_r,
  input [29:0] io_pmp_6_addr,
  input [31:0] io_pmp_6_mask,
  input io_pmp_7_cfg_l,
  input [1:0] io_pmp_7_cfg_a,
  input io_pmp_7_cfg_x,
  input io_pmp_7_cfg_w,
  input io_pmp_7_cfg_r,
  input [29:0] io_pmp_7_addr,
  input [31:0] io_pmp_7_mask,
  input [31:0] io_addr,
  output io_r,
  output io_w,
  output io_x,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire default_ ;  
   wire [31:0] _res_hit_T_1 ;  
   wire [31:0] _res_hit_T_3 ;  
   wire [31:0] _res_hit_T_5 ;  
   wire [31:0] _res_hit_T_7 ;  
   wire _res_hit_T_8 ;  
   wire [31:0] _res_hit_T_14 ;  
   wire [31:0] _res_hit_T_16 ;  
   wire _res_hit_T_18 ;  
   wire _res_hit_T_24 ;  
   wire _res_hit_T_25 ;  
   wire _res_hit_T_26 ;  
   wire res_hit ;  
   wire res_ignore ;  
   wire res_cur_cfg_r ;  
   wire res_cur_cfg_w ;  
   wire res_cur_cfg_x ;  
   wire _res_T_44_cfg_x ;  
   wire _res_T_44_cfg_w ;  
   wire _res_T_44_cfg_r ;  
   wire [31:0] _res_hit_T_32 ;  
   wire [31:0] _res_hit_T_34 ;  
   wire _res_hit_T_35 ;  
   wire [31:0] _res_hit_T_41 ;  
   wire [31:0] _res_hit_T_43 ;  
   wire _res_hit_T_45 ;  
   wire _res_hit_T_52 ;  
   wire _res_hit_T_53 ;  
   wire res_hit_1 ;  
   wire res_ignore_1 ;  
   wire res_cur_1_cfg_r ;  
   wire res_cur_1_cfg_w ;  
   wire res_cur_1_cfg_x ;  
   wire _res_T_89_cfg_x ;  
   wire _res_T_89_cfg_w ;  
   wire _res_T_89_cfg_r ;  
   wire [31:0] _res_hit_T_59 ;  
   wire [31:0] _res_hit_T_61 ;  
   wire _res_hit_T_62 ;  
   wire [31:0] _res_hit_T_68 ;  
   wire [31:0] _res_hit_T_70 ;  
   wire _res_hit_T_72 ;  
   wire _res_hit_T_79 ;  
   wire _res_hit_T_80 ;  
   wire res_hit_2 ;  
   wire res_ignore_2 ;  
   wire res_cur_2_cfg_r ;  
   wire res_cur_2_cfg_w ;  
   wire res_cur_2_cfg_x ;  
   wire _res_T_134_cfg_x ;  
   wire _res_T_134_cfg_w ;  
   wire _res_T_134_cfg_r ;  
   wire [31:0] _res_hit_T_86 ;  
   wire [31:0] _res_hit_T_88 ;  
   wire _res_hit_T_89 ;  
   wire [31:0] _res_hit_T_95 ;  
   wire [31:0] _res_hit_T_97 ;  
   wire _res_hit_T_99 ;  
   wire _res_hit_T_106 ;  
   wire _res_hit_T_107 ;  
   wire res_hit_3 ;  
   wire res_ignore_3 ;  
   wire res_cur_3_cfg_r ;  
   wire res_cur_3_cfg_w ;  
   wire res_cur_3_cfg_x ;  
   wire _res_T_179_cfg_x ;  
   wire _res_T_179_cfg_w ;  
   wire _res_T_179_cfg_r ;  
   wire [31:0] _res_hit_T_113 ;  
   wire [31:0] _res_hit_T_115 ;  
   wire _res_hit_T_116 ;  
   wire [31:0] _res_hit_T_122 ;  
   wire [31:0] _res_hit_T_124 ;  
   wire _res_hit_T_126 ;  
   wire _res_hit_T_133 ;  
   wire _res_hit_T_134 ;  
   wire res_hit_4 ;  
   wire res_ignore_4 ;  
   wire res_cur_4_cfg_r ;  
   wire res_cur_4_cfg_w ;  
   wire res_cur_4_cfg_x ;  
   wire _res_T_224_cfg_x ;  
   wire _res_T_224_cfg_w ;  
   wire _res_T_224_cfg_r ;  
   wire [31:0] _res_hit_T_140 ;  
   wire [31:0] _res_hit_T_142 ;  
   wire _res_hit_T_143 ;  
   wire [31:0] _res_hit_T_149 ;  
   wire [31:0] _res_hit_T_151 ;  
   wire _res_hit_T_153 ;  
   wire _res_hit_T_160 ;  
   wire _res_hit_T_161 ;  
   wire res_hit_5 ;  
   wire res_ignore_5 ;  
   wire res_cur_5_cfg_r ;  
   wire res_cur_5_cfg_w ;  
   wire res_cur_5_cfg_x ;  
   wire _res_T_269_cfg_x ;  
   wire _res_T_269_cfg_w ;  
   wire _res_T_269_cfg_r ;  
   wire [31:0] _res_hit_T_167 ;  
   wire [31:0] _res_hit_T_169 ;  
   wire _res_hit_T_170 ;  
   wire [31:0] _res_hit_T_176 ;  
   wire [31:0] _res_hit_T_178 ;  
   wire _res_hit_T_180 ;  
   wire _res_hit_T_187 ;  
   wire _res_hit_T_188 ;  
   wire res_hit_6 ;  
   wire res_ignore_6 ;  
   wire res_cur_6_cfg_r ;  
   wire res_cur_6_cfg_w ;  
   wire res_cur_6_cfg_x ;  
   wire _res_T_314_cfg_x ;  
   wire _res_T_314_cfg_w ;  
   wire _res_T_314_cfg_r ;  
   wire [31:0] _res_hit_T_194 ;  
   wire [31:0] _res_hit_T_196 ;  
   wire _res_hit_T_197 ;  
   wire _res_hit_T_215 ;  
   wire res_hit_7 ;  
   wire res_ignore_7 ;  
   wire res_cur_7_cfg_r ;  
   wire res_cur_7_cfg_w ;  
   wire res_cur_7_cfg_x ;  
   wire [29:0] PMPChecker_2_covSum ;  
  assign default_=io_prv>2'h1; 
  assign _res_hit_T_1={io_pmp_7_addr,2'h0}; 
  assign _res_hit_T_3=~_res_hit_T_1|32'h3; 
  assign _res_hit_T_5=io_addr^~_res_hit_T_3; 
  assign _res_hit_T_7=_res_hit_T_5&~io_pmp_7_mask; 
  assign _res_hit_T_8=_res_hit_T_7==32'h0; 
  assign _res_hit_T_14={io_pmp_6_addr,2'h0}; 
  assign _res_hit_T_16=~_res_hit_T_14|32'h3; 
  assign _res_hit_T_18=io_addr<~_res_hit_T_16; 
  assign _res_hit_T_24=io_addr<~_res_hit_T_3; 
  assign _res_hit_T_25=~_res_hit_T_18&_res_hit_T_24; 
  assign _res_hit_T_26=io_pmp_7_cfg_a[0]&_res_hit_T_25; 
  assign res_hit=io_pmp_7_cfg_a[1] ? _res_hit_T_8:_res_hit_T_26; 
  assign res_ignore=default_&~io_pmp_7_cfg_l; 
  assign res_cur_cfg_r=io_pmp_7_cfg_r|res_ignore; 
  assign res_cur_cfg_w=io_pmp_7_cfg_w|res_ignore; 
  assign res_cur_cfg_x=io_pmp_7_cfg_x|res_ignore; 
  assign _res_T_44_cfg_x=res_hit ? res_cur_cfg_x:default_; 
  assign _res_T_44_cfg_w=res_hit ? res_cur_cfg_w:default_; 
  assign _res_T_44_cfg_r=res_hit ? res_cur_cfg_r:default_; 
  assign _res_hit_T_32=io_addr^~_res_hit_T_16; 
  assign _res_hit_T_34=_res_hit_T_32&~io_pmp_6_mask; 
  assign _res_hit_T_35=_res_hit_T_34==32'h0; 
  assign _res_hit_T_41={io_pmp_5_addr,2'h0}; 
  assign _res_hit_T_43=~_res_hit_T_41|32'h3; 
  assign _res_hit_T_45=io_addr<~_res_hit_T_43; 
  assign _res_hit_T_52=~_res_hit_T_45&_res_hit_T_18; 
  assign _res_hit_T_53=io_pmp_6_cfg_a[0]&_res_hit_T_52; 
  assign res_hit_1=io_pmp_6_cfg_a[1] ? _res_hit_T_35:_res_hit_T_53; 
  assign res_ignore_1=default_&~io_pmp_6_cfg_l; 
  assign res_cur_1_cfg_r=io_pmp_6_cfg_r|res_ignore_1; 
  assign res_cur_1_cfg_w=io_pmp_6_cfg_w|res_ignore_1; 
  assign res_cur_1_cfg_x=io_pmp_6_cfg_x|res_ignore_1; 
  assign _res_T_89_cfg_x=res_hit_1 ? res_cur_1_cfg_x:_res_T_44_cfg_x; 
  assign _res_T_89_cfg_w=res_hit_1 ? res_cur_1_cfg_w:_res_T_44_cfg_w; 
  assign _res_T_89_cfg_r=res_hit_1 ? res_cur_1_cfg_r:_res_T_44_cfg_r; 
  assign _res_hit_T_59=io_addr^~_res_hit_T_43; 
  assign _res_hit_T_61=_res_hit_T_59&~io_pmp_5_mask; 
  assign _res_hit_T_62=_res_hit_T_61==32'h0; 
  assign _res_hit_T_68={io_pmp_4_addr,2'h0}; 
  assign _res_hit_T_70=~_res_hit_T_68|32'h3; 
  assign _res_hit_T_72=io_addr<~_res_hit_T_70; 
  assign _res_hit_T_79=~_res_hit_T_72&_res_hit_T_45; 
  assign _res_hit_T_80=io_pmp_5_cfg_a[0]&_res_hit_T_79; 
  assign res_hit_2=io_pmp_5_cfg_a[1] ? _res_hit_T_62:_res_hit_T_80; 
  assign res_ignore_2=default_&~io_pmp_5_cfg_l; 
  assign res_cur_2_cfg_r=io_pmp_5_cfg_r|res_ignore_2; 
  assign res_cur_2_cfg_w=io_pmp_5_cfg_w|res_ignore_2; 
  assign res_cur_2_cfg_x=io_pmp_5_cfg_x|res_ignore_2; 
  assign _res_T_134_cfg_x=res_hit_2 ? res_cur_2_cfg_x:_res_T_89_cfg_x; 
  assign _res_T_134_cfg_w=res_hit_2 ? res_cur_2_cfg_w:_res_T_89_cfg_w; 
  assign _res_T_134_cfg_r=res_hit_2 ? res_cur_2_cfg_r:_res_T_89_cfg_r; 
  assign _res_hit_T_86=io_addr^~_res_hit_T_70; 
  assign _res_hit_T_88=_res_hit_T_86&~io_pmp_4_mask; 
  assign _res_hit_T_89=_res_hit_T_88==32'h0; 
  assign _res_hit_T_95={io_pmp_3_addr,2'h0}; 
  assign _res_hit_T_97=~_res_hit_T_95|32'h3; 
  assign _res_hit_T_99=io_addr<~_res_hit_T_97; 
  assign _res_hit_T_106=~_res_hit_T_99&_res_hit_T_72; 
  assign _res_hit_T_107=io_pmp_4_cfg_a[0]&_res_hit_T_106; 
  assign res_hit_3=io_pmp_4_cfg_a[1] ? _res_hit_T_89:_res_hit_T_107; 
  assign res_ignore_3=default_&~io_pmp_4_cfg_l; 
  assign res_cur_3_cfg_r=io_pmp_4_cfg_r|res_ignore_3; 
  assign res_cur_3_cfg_w=io_pmp_4_cfg_w|res_ignore_3; 
  assign res_cur_3_cfg_x=io_pmp_4_cfg_x|res_ignore_3; 
  assign _res_T_179_cfg_x=res_hit_3 ? res_cur_3_cfg_x:_res_T_134_cfg_x; 
  assign _res_T_179_cfg_w=res_hit_3 ? res_cur_3_cfg_w:_res_T_134_cfg_w; 
  assign _res_T_179_cfg_r=res_hit_3 ? res_cur_3_cfg_r:_res_T_134_cfg_r; 
  assign _res_hit_T_113=io_addr^~_res_hit_T_97; 
  assign _res_hit_T_115=_res_hit_T_113&~io_pmp_3_mask; 
  assign _res_hit_T_116=_res_hit_T_115==32'h0; 
  assign _res_hit_T_122={io_pmp_2_addr,2'h0}; 
  assign _res_hit_T_124=~_res_hit_T_122|32'h3; 
  assign _res_hit_T_126=io_addr<~_res_hit_T_124; 
  assign _res_hit_T_133=~_res_hit_T_126&_res_hit_T_99; 
  assign _res_hit_T_134=io_pmp_3_cfg_a[0]&_res_hit_T_133; 
  assign res_hit_4=io_pmp_3_cfg_a[1] ? _res_hit_T_116:_res_hit_T_134; 
  assign res_ignore_4=default_&~io_pmp_3_cfg_l; 
  assign res_cur_4_cfg_r=io_pmp_3_cfg_r|res_ignore_4; 
  assign res_cur_4_cfg_w=io_pmp_3_cfg_w|res_ignore_4; 
  assign res_cur_4_cfg_x=io_pmp_3_cfg_x|res_ignore_4; 
  assign _res_T_224_cfg_x=res_hit_4 ? res_cur_4_cfg_x:_res_T_179_cfg_x; 
  assign _res_T_224_cfg_w=res_hit_4 ? res_cur_4_cfg_w:_res_T_179_cfg_w; 
  assign _res_T_224_cfg_r=res_hit_4 ? res_cur_4_cfg_r:_res_T_179_cfg_r; 
  assign _res_hit_T_140=io_addr^~_res_hit_T_124; 
  assign _res_hit_T_142=_res_hit_T_140&~io_pmp_2_mask; 
  assign _res_hit_T_143=_res_hit_T_142==32'h0; 
  assign _res_hit_T_149={io_pmp_1_addr,2'h0}; 
  assign _res_hit_T_151=~_res_hit_T_149|32'h3; 
  assign _res_hit_T_153=io_addr<~_res_hit_T_151; 
  assign _res_hit_T_160=~_res_hit_T_153&_res_hit_T_126; 
  assign _res_hit_T_161=io_pmp_2_cfg_a[0]&_res_hit_T_160; 
  assign res_hit_5=io_pmp_2_cfg_a[1] ? _res_hit_T_143:_res_hit_T_161; 
  assign res_ignore_5=default_&~io_pmp_2_cfg_l; 
  assign res_cur_5_cfg_r=io_pmp_2_cfg_r|res_ignore_5; 
  assign res_cur_5_cfg_w=io_pmp_2_cfg_w|res_ignore_5; 
  assign res_cur_5_cfg_x=io_pmp_2_cfg_x|res_ignore_5; 
  assign _res_T_269_cfg_x=res_hit_5 ? res_cur_5_cfg_x:_res_T_224_cfg_x; 
  assign _res_T_269_cfg_w=res_hit_5 ? res_cur_5_cfg_w:_res_T_224_cfg_w; 
  assign _res_T_269_cfg_r=res_hit_5 ? res_cur_5_cfg_r:_res_T_224_cfg_r; 
  assign _res_hit_T_167=io_addr^~_res_hit_T_151; 
  assign _res_hit_T_169=_res_hit_T_167&~io_pmp_1_mask; 
  assign _res_hit_T_170=_res_hit_T_169==32'h0; 
  assign _res_hit_T_176={io_pmp_0_addr,2'h0}; 
  assign _res_hit_T_178=~_res_hit_T_176|32'h3; 
  assign _res_hit_T_180=io_addr<~_res_hit_T_178; 
  assign _res_hit_T_187=~_res_hit_T_180&_res_hit_T_153; 
  assign _res_hit_T_188=io_pmp_1_cfg_a[0]&_res_hit_T_187; 
  assign res_hit_6=io_pmp_1_cfg_a[1] ? _res_hit_T_170:_res_hit_T_188; 
  assign res_ignore_6=default_&~io_pmp_1_cfg_l; 
  assign res_cur_6_cfg_r=io_pmp_1_cfg_r|res_ignore_6; 
  assign res_cur_6_cfg_w=io_pmp_1_cfg_w|res_ignore_6; 
  assign res_cur_6_cfg_x=io_pmp_1_cfg_x|res_ignore_6; 
  assign _res_T_314_cfg_x=res_hit_6 ? res_cur_6_cfg_x:_res_T_269_cfg_x; 
  assign _res_T_314_cfg_w=res_hit_6 ? res_cur_6_cfg_w:_res_T_269_cfg_w; 
  assign _res_T_314_cfg_r=res_hit_6 ? res_cur_6_cfg_r:_res_T_269_cfg_r; 
  assign _res_hit_T_194=io_addr^~_res_hit_T_178; 
  assign _res_hit_T_196=_res_hit_T_194&~io_pmp_0_mask; 
  assign _res_hit_T_197=_res_hit_T_196==32'h0; 
  assign _res_hit_T_215=io_pmp_0_cfg_a[0]&_res_hit_T_180; 
  assign res_hit_7=io_pmp_0_cfg_a[1] ? _res_hit_T_197:_res_hit_T_215; 
  assign res_ignore_7=default_&~io_pmp_0_cfg_l; 
  assign res_cur_7_cfg_r=io_pmp_0_cfg_r|res_ignore_7; 
  assign res_cur_7_cfg_w=io_pmp_0_cfg_w|res_ignore_7; 
  assign res_cur_7_cfg_x=io_pmp_0_cfg_x|res_ignore_7; 
  assign io_r=res_hit_7 ? res_cur_7_cfg_r:_res_T_314_cfg_r; 
  assign io_w=res_hit_7 ? res_cur_7_cfg_w:_res_T_314_cfg_w; 
  assign io_x=res_hit_7 ? res_cur_7_cfg_x:_res_T_314_cfg_x; 
  assign PMPChecker_2_covSum=30'h0; 
  assign io_covSum=PMPChecker_2_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module MulAddRecFNPipe (
  input clock,
  input reset,
  input io_validin,
  input [1:0] io_op,
  input [32:0] io_a,
  input [32:0] io_b,
  input [32:0] io_c,
  input [2:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [1:0] mulAddRecFNToRaw_preMul_io_op ;  
   wire [32:0] mulAddRecFNToRaw_preMul_io_a ;  
   wire [32:0] mulAddRecFNToRaw_preMul_io_b ;  
   wire [32:0] mulAddRecFNToRaw_preMul_io_c ;  
   wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA ;  
   wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB ;  
   wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfA ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfB ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_signProd ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC ;  
   wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant ;  
   wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist ;  
   wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC ;  
   wire [29:0] mulAddRecFNToRaw_preMul_io_covSum ;  
   wire mulAddRecFNToRaw_preMul_metaAssert ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_signProd ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC ;  
   wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant ;  
   wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist ;  
   wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC ;  
   wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult ;  
   wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode ;  
   wire mulAddRecFNToRaw_postMul_io_invalidExc ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_isNaN ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_isInf ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_isZero ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_sign ;  
   wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp ;  
   wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig ;  
   wire [29:0] mulAddRecFNToRaw_postMul_io_covSum ;  
   wire mulAddRecFNToRaw_postMul_metaAssert ;  
   wire roundRawFNToRecFN_io_invalidExc ;  
   wire roundRawFNToRecFN_io_infiniteExc ;  
   wire roundRawFNToRecFN_io_in_isNaN ;  
   wire roundRawFNToRecFN_io_in_isInf ;  
   wire roundRawFNToRecFN_io_in_isZero ;  
   wire roundRawFNToRecFN_io_in_sign ;  
   wire [9:0] roundRawFNToRecFN_io_in_sExp ;  
   wire [26:0] roundRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundRawFNToRecFN_io_roundingMode ;  
   wire roundRawFNToRecFN_io_detectTininess ;  
   wire [32:0] roundRawFNToRecFN_io_out ;  
   wire [4:0] roundRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundRawFNToRecFN_io_covSum ;  
   wire roundRawFNToRecFN_metaAssert ;  
   wire [47:0] _mulAddResult_T ;  
   wire [48:0] mulAddResult ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny ;  
   reg [31:0] _RAND_0 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB ;  
   reg [31:0] _RAND_1 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA ;  
   reg [31:0] _RAND_2 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA ;  
   reg [31:0] _RAND_3 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB ;  
   reg [31:0] _RAND_4 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB ;  
   reg [31:0] _RAND_5 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd ;  
   reg [31:0] _RAND_6 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC ;  
   reg [31:0] _RAND_7 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC ;  
   reg [31:0] _RAND_8 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC ;  
   reg [31:0] _RAND_9 ;  
   reg [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum ;  
   reg [31:0] _RAND_10 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags ;  
   reg [31:0] _RAND_11 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant ;  
   reg [31:0] _RAND_12 ;  
   reg [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist ;  
   reg [31:0] _RAND_13 ;  
   reg [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC ;  
   reg [31:0] _RAND_14 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC ;  
   reg [31:0] _RAND_15 ;  
   reg [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult_b ;  
   reg [63:0] _RAND_16 ;  
   reg [2:0] mulAddRecFNToRaw_postMul_io_roundingMode_b ;  
   reg [31:0] _RAND_17 ;  
   reg [2:0] roundingMode_stage0_b ;  
   reg [31:0] _RAND_18 ;  
   reg detectTininess_stage0_b ;  
   reg [31:0] _RAND_19 ;  
   reg valid_stage0_v ;  
   reg [31:0] _RAND_20 ;  
   reg roundRawFNToRecFN_io_invalidExc_b ;  
   reg [31:0] _RAND_21 ;  
   reg roundRawFNToRecFN_io_in_b_isNaN ;  
   reg [31:0] _RAND_22 ;  
   reg roundRawFNToRecFN_io_in_b_isInf ;  
   reg [31:0] _RAND_23 ;  
   reg roundRawFNToRecFN_io_in_b_isZero ;  
   reg [31:0] _RAND_24 ;  
   reg roundRawFNToRecFN_io_in_b_sign ;  
   reg [31:0] _RAND_25 ;  
   reg [9:0] roundRawFNToRecFN_io_in_b_sExp ;  
   reg [31:0] _RAND_26 ;  
   reg [26:0] roundRawFNToRecFN_io_in_b_sig ;  
   reg [31:0] _RAND_27 ;  
   reg [2:0] roundRawFNToRecFN_io_roundingMode_b ;  
   reg [31:0] _RAND_28 ;  
   reg roundRawFNToRecFN_io_detectTininess_b ;  
   reg [31:0] _RAND_29 ;  
   reg MulAddRecFNPipe_state ;  
   reg [31:0] _RAND_30 ;  
   reg MulAddRecFNPipe_cov[0:1] ;  
   reg [31:0] _RAND_31 ;  
   wire MulAddRecFNPipe_cov_read_data ;  
   wire MulAddRecFNPipe_cov_read_addr ;  
   wire MulAddRecFNPipe_cov_write_data ;  
   wire MulAddRecFNPipe_cov_write_addr ;  
   wire MulAddRecFNPipe_cov_write_mask ;  
   wire MulAddRecFNPipe_cov_write_en ;  
   reg [29:0] MulAddRecFNPipe_covSum ;  
   reg [31:0] _RAND_32 ;  
   wire valid_stage0_v_shl ;  
   wire valid_stage0_v_pad ;  
   wire [29:0] mulAddRecFNToRaw_preMul_sum ;  
   wire [29:0] mulAddRecFNToRaw_postMul_sum ;  
   wire [29:0] roundRawFNToRecFN_sum ;  
   wire mulAddRecFNToRaw_preMul_metaAssert_wire ;  
   wire mulAddRecFNToRaw_postMul_metaAssert_wire ;  
   wire roundRawFNToRecFN_metaAssert_wire ;  
   wire MulAddRecFNPipe_or2 ;  
   wire MulAddRecFNPipe_or0 ;  
   reg MulAddRecFNPipe_metaAssert ;  
   reg [31:0] _RAND_33 ;  
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul(.io_op(mulAddRecFNToRaw_preMul_io_op),.io_a(mulAddRecFNToRaw_preMul_io_a),.io_b(mulAddRecFNToRaw_preMul_io_b),.io_c(mulAddRecFNToRaw_preMul_io_c),.io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),.io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),.io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),.io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),.io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),.io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),.io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),.io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),.io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),.io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),.io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),.io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),.io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),.io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),.io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),.io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),.io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),.io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),.io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),.io_covSum(mulAddRecFNToRaw_preMul_io_covSum),.metaAssert(mulAddRecFNToRaw_preMul_metaAssert)); 
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul(.io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),.io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),.io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),.io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),.io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),.io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),.io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),.io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),.io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),.io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),.io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),.io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),.io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),.io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),.io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),.io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),.io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),.io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),.io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),.io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),.io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),.io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),.io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),.io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),.io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),.io_covSum(mulAddRecFNToRaw_postMul_io_covSum),.metaAssert(mulAddRecFNToRaw_postMul_metaAssert)); 
  RoundRawFNToRecFN_2 roundRawFNToRecFN(.io_invalidExc(roundRawFNToRecFN_io_invalidExc),.io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),.io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),.io_in_isInf(roundRawFNToRecFN_io_in_isInf),.io_in_isZero(roundRawFNToRecFN_io_in_isZero),.io_in_sign(roundRawFNToRecFN_io_in_sign),.io_in_sExp(roundRawFNToRecFN_io_in_sExp),.io_in_sig(roundRawFNToRecFN_io_in_sig),.io_roundingMode(roundRawFNToRecFN_io_roundingMode),.io_detectTininess(roundRawFNToRecFN_io_detectTininess),.io_out(roundRawFNToRecFN_io_out),.io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),.io_covSum(roundRawFNToRecFN_io_covSum),.metaAssert(roundRawFNToRecFN_metaAssert)); 
  assign _mulAddResult_T=mulAddRecFNToRaw_preMul_io_mulAddA*mulAddRecFNToRaw_preMul_io_mulAddB; 
  assign mulAddResult=_mulAddResult_T+mulAddRecFNToRaw_preMul_io_mulAddC; 
  assign io_out=roundRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundRawFNToRecFN_io_exceptionFlags; 
  assign mulAddRecFNToRaw_preMul_io_op=io_op; 
  assign mulAddRecFNToRaw_preMul_io_a=io_a; 
  assign mulAddRecFNToRaw_preMul_io_b=io_b; 
  assign mulAddRecFNToRaw_preMul_io_c=io_c; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd=mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum=mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags=mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant=mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist=mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC; 
  assign mulAddRecFNToRaw_postMul_io_mulAddResult=mulAddRecFNToRaw_postMul_io_mulAddResult_b; 
  assign mulAddRecFNToRaw_postMul_io_roundingMode=mulAddRecFNToRaw_postMul_io_roundingMode_b; 
  assign roundRawFNToRecFN_io_invalidExc=roundRawFNToRecFN_io_invalidExc_b; 
  assign roundRawFNToRecFN_io_infiniteExc=1'h0; 
  assign roundRawFNToRecFN_io_in_isNaN=roundRawFNToRecFN_io_in_b_isNaN; 
  assign roundRawFNToRecFN_io_in_isInf=roundRawFNToRecFN_io_in_b_isInf; 
  assign roundRawFNToRecFN_io_in_isZero=roundRawFNToRecFN_io_in_b_isZero; 
  assign roundRawFNToRecFN_io_in_sign=roundRawFNToRecFN_io_in_b_sign; 
  assign roundRawFNToRecFN_io_in_sExp=roundRawFNToRecFN_io_in_b_sExp; 
  assign roundRawFNToRecFN_io_in_sig=roundRawFNToRecFN_io_in_b_sig; 
  assign roundRawFNToRecFN_io_roundingMode=roundRawFNToRecFN_io_roundingMode_b; 
  assign roundRawFNToRecFN_io_detectTininess=roundRawFNToRecFN_io_detectTininess_b; 
  assign MulAddRecFNPipe_cov_read_addr=MulAddRecFNPipe_state; 
  assign MulAddRecFNPipe_cov_read_data=MulAddRecFNPipe_cov[MulAddRecFNPipe_cov_read_addr]; 
  assign MulAddRecFNPipe_cov_write_data=1'h1; 
  assign MulAddRecFNPipe_cov_write_addr=MulAddRecFNPipe_state; 
  assign MulAddRecFNPipe_cov_write_mask=1'h1; 
  assign MulAddRecFNPipe_cov_write_en=1'h1; 
  assign valid_stage0_v_shl=valid_stage0_v; 
  assign valid_stage0_v_pad=valid_stage0_v_shl; 
  assign mulAddRecFNToRaw_preMul_sum=MulAddRecFNPipe_covSum+mulAddRecFNToRaw_preMul_io_covSum; 
  assign mulAddRecFNToRaw_postMul_sum=mulAddRecFNToRaw_preMul_sum+mulAddRecFNToRaw_postMul_io_covSum; 
  assign roundRawFNToRecFN_sum=mulAddRecFNToRaw_postMul_sum+roundRawFNToRecFN_io_covSum; 
  assign io_covSum=roundRawFNToRecFN_sum; 
  assign mulAddRecFNToRaw_preMul_metaAssert_wire=mulAddRecFNToRaw_preMul_metaAssert; 
  assign mulAddRecFNToRaw_postMul_metaAssert_wire=mulAddRecFNToRaw_postMul_metaAssert; 
  assign roundRawFNToRecFN_metaAssert_wire=roundRawFNToRecFN_metaAssert; 
  assign MulAddRecFNPipe_or2=mulAddRecFNToRaw_postMul_metaAssert_wire|roundRawFNToRecFN_metaAssert_wire; 
  assign MulAddRecFNPipe_or0=mulAddRecFNToRaw_preMul_metaAssert_wire|MulAddRecFNPipe_or2; 
  assign metaAssert=MulAddRecFNPipe_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <=mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <=mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <=mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <=mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <=mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <=mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <=mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <=mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <=mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <=mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <=10'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <=mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <=mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <=mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <=5'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <=mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <=26'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <=mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <=mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_mulAddResult_b <=49'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_mulAddResult_b <=mulAddResult;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_roundingMode_b <=3'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_roundingMode_b <=io_roundingMode;
               end 
         if (metaReset)
            begin 
              roundingMode_stage0_b <=3'h0;
            end 
          else 
            if (io_validin)
               begin 
                 roundingMode_stage0_b <=io_roundingMode;
               end 
         if (metaReset)
            begin 
              detectTininess_stage0_b <=1'h0;
            end 
          else 
            begin 
              detectTininess_stage0_b <=io_validin|detectTininess_stage0_b;
            end 
         if (metaReset)
            begin 
              valid_stage0_v <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 valid_stage0_v <=1'h0;
               end 
             else 
               begin 
                 valid_stage0_v <=io_validin;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_invalidExc_b <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_invalidExc_b <=mulAddRecFNToRaw_postMul_io_invalidExc;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_isNaN <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_isNaN <=mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_isInf <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_isInf <=mulAddRecFNToRaw_postMul_io_rawOut_isInf;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_isZero <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_isZero <=mulAddRecFNToRaw_postMul_io_rawOut_isZero;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_sign <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_sign <=mulAddRecFNToRaw_postMul_io_rawOut_sign;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_sExp <=10'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_sExp <=mulAddRecFNToRaw_postMul_io_rawOut_sExp;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_sig <=27'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_sig <=mulAddRecFNToRaw_postMul_io_rawOut_sig;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_roundingMode_b <=3'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_roundingMode_b <=roundingMode_stage0_b;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_detectTininess_b <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_detectTininess_b <=detectTininess_stage0_b;
               end 
         MulAddRecFNPipe_state <=valid_stage0_v_pad;
         if (!(MulAddRecFNPipe_cov_read_data))
            begin 
              MulAddRecFNPipe_covSum <=MulAddRecFNPipe_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              MulAddRecFNPipe_metaAssert <=1'h0;
            end 
          else 
            begin 
              MulAddRecFNPipe_metaAssert <=MulAddRecFNPipe_metaAssert|MulAddRecFNPipe_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (MulAddRecFNPipe_cov_write_en&MulAddRecFNPipe_cov_write_mask)
            begin 
              MulAddRecFNPipe_cov [MulAddRecFNPipe_cov_write_addr]<=MulAddRecFNPipe_cov_write_data;
            end 
       end
  
endmodule
 
module CompareRecFN (
  input [64:0] io_a,
  input [64:0] io_b,
  input io_signaling,
  output io_lt,
  output io_eq,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [11:0] rawA_exp ;  
   wire rawA_isZero ;  
   wire rawA_isSpecial ;  
   wire rawA__isNaN ;  
   wire rawA__isInf ;  
   wire rawA__sign ;  
   wire [12:0] rawA__sExp ;  
   wire rawA_out_sig_hi_lo ;  
   wire [51:0] rawA_out_sig_lo ;  
   wire [53:0] rawA__sig ;  
   wire [11:0] rawB_exp ;  
   wire rawB_isZero ;  
   wire rawB_isSpecial ;  
   wire rawB__isNaN ;  
   wire rawB__isInf ;  
   wire rawB__sign ;  
   wire [12:0] rawB__sExp ;  
   wire rawB_out_sig_hi_lo ;  
   wire [51:0] rawB_out_sig_lo ;  
   wire [53:0] rawB__sig ;  
   wire ordered ;  
   wire bothInfs ;  
   wire bothZeros ;  
   wire eqExps ;  
   wire _common_ltMags_T ;  
   wire _common_ltMags_T_1 ;  
   wire _common_ltMags_T_2 ;  
   wire common_ltMags ;  
   wire _common_eqMags_T ;  
   wire common_eqMags ;  
   wire _ordered_lt_T_2 ;  
   wire _ordered_lt_T_5 ;  
   wire _ordered_lt_T_7 ;  
   wire _ordered_lt_T_9 ;  
   wire _ordered_lt_T_10 ;  
   wire _ordered_lt_T_11 ;  
   wire _ordered_lt_T_12 ;  
   wire ordered_lt ;  
   wire _ordered_eq_T ;  
   wire _ordered_eq_T_1 ;  
   wire _ordered_eq_T_2 ;  
   wire ordered_eq ;  
   wire _invalid_T_2 ;  
   wire _invalid_T_5 ;  
   wire _invalid_T_6 ;  
   wire _invalid_T_8 ;  
   wire invalid ;  
   wire [29:0] CompareRecFN_covSum ;  
  assign rawA_exp=io_a[63:52]; 
  assign rawA_isZero=rawA_exp[11:9]==3'h0; 
  assign rawA_isSpecial=rawA_exp[11:10]==2'h3; 
  assign rawA__isNaN=rawA_isSpecial&rawA_exp[9]; 
  assign rawA__isInf=rawA_isSpecial&~rawA_exp[9]; 
  assign rawA__sign=io_a[64]; 
  assign rawA__sExp={1'b0,$signed(rawA_exp)}; 
  assign rawA_out_sig_hi_lo=~rawA_isZero; 
  assign rawA_out_sig_lo=io_a[51:0]; 
  assign rawA__sig={1'h0,rawA_out_sig_hi_lo,rawA_out_sig_lo}; 
  assign rawB_exp=io_b[63:52]; 
  assign rawB_isZero=rawB_exp[11:9]==3'h0; 
  assign rawB_isSpecial=rawB_exp[11:10]==2'h3; 
  assign rawB__isNaN=rawB_isSpecial&rawB_exp[9]; 
  assign rawB__isInf=rawB_isSpecial&~rawB_exp[9]; 
  assign rawB__sign=io_b[64]; 
  assign rawB__sExp={1'b0,$signed(rawB_exp)}; 
  assign rawB_out_sig_hi_lo=~rawB_isZero; 
  assign rawB_out_sig_lo=io_b[51:0]; 
  assign rawB__sig={1'h0,rawB_out_sig_hi_lo,rawB_out_sig_lo}; 
  assign ordered=~rawA__isNaN&~rawB__isNaN; 
  assign bothInfs=rawA__isInf&rawB__isInf; 
  assign bothZeros=rawA_isZero&rawB_isZero; 
  assign eqExps=$signed(rawA__sExp)==$signed(rawB__sExp); 
  assign _common_ltMags_T=$signed(rawA__sExp)<$signed(rawB__sExp); 
  assign _common_ltMags_T_1=rawA__sig<rawB__sig; 
  assign _common_ltMags_T_2=eqExps&_common_ltMags_T_1; 
  assign common_ltMags=_common_ltMags_T|_common_ltMags_T_2; 
  assign _common_eqMags_T=rawA__sig==rawB__sig; 
  assign common_eqMags=eqExps&_common_eqMags_T; 
  assign _ordered_lt_T_2=rawA__sign&~rawB__sign; 
  assign _ordered_lt_T_5=rawA__sign&~common_ltMags; 
  assign _ordered_lt_T_7=_ordered_lt_T_5&~common_eqMags; 
  assign _ordered_lt_T_9=~rawB__sign&common_ltMags; 
  assign _ordered_lt_T_10=_ordered_lt_T_7|_ordered_lt_T_9; 
  assign _ordered_lt_T_11=~bothInfs&_ordered_lt_T_10; 
  assign _ordered_lt_T_12=_ordered_lt_T_2|_ordered_lt_T_11; 
  assign ordered_lt=~bothZeros&_ordered_lt_T_12; 
  assign _ordered_eq_T=rawA__sign==rawB__sign; 
  assign _ordered_eq_T_1=bothInfs|common_eqMags; 
  assign _ordered_eq_T_2=_ordered_eq_T&_ordered_eq_T_1; 
  assign ordered_eq=bothZeros|_ordered_eq_T_2; 
  assign _invalid_T_2=rawA__isNaN&~rawA__sig[51]; 
  assign _invalid_T_5=rawB__isNaN&~rawB__sig[51]; 
  assign _invalid_T_6=_invalid_T_2|_invalid_T_5; 
  assign _invalid_T_8=io_signaling&~ordered; 
  assign invalid=_invalid_T_6|_invalid_T_8; 
  assign io_lt=ordered&ordered_lt; 
  assign io_eq=ordered&ordered_eq; 
  assign io_exceptionFlags={invalid,4'h0}; 
  assign CompareRecFN_covSum=30'h0; 
  assign io_covSum=CompareRecFN_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module RecFNToIN (
  input [64:0] io_in,
  input [2:0] io_roundingMode,
  input io_signedOut,
  output [63:0] io_out,
  output [2:0] io_intExceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [11:0] rawIn_exp ;  
   wire rawIn_isZero ;  
   wire rawIn_isSpecial ;  
   wire rawIn__isNaN ;  
   wire rawIn__isInf ;  
   wire rawIn__sign ;  
   wire [12:0] rawIn__sExp ;  
   wire rawIn_out_sig_hi_lo ;  
   wire [51:0] rawIn_out_sig_lo ;  
   wire [53:0] rawIn__sig ;  
   wire magGeOne ;  
   wire [10:0] posExp ;  
   wire _magJustBelowOne_T_1 ;  
   wire magJustBelowOne ;  
   wire roundingMode_near_even ;  
   wire roundingMode_min ;  
   wire roundingMode_max ;  
   wire roundingMode_near_maxMag ;  
   wire roundingMode_odd ;  
   wire [51:0] shiftedSig_lo ;  
   wire [52:0] _shiftedSig_T ;  
   wire [5:0] _shiftedSig_T_2 ;  
   wire [115:0] _GEN_0 ;  
   wire [115:0] shiftedSig ;  
   wire [64:0] alignedSig_hi ;  
   wire alignedSig_lo ;  
   wire [65:0] alignedSig ;  
   wire [63:0] unroundedInt ;  
   wire _common_inexact_T_1 ;  
   wire common_inexact ;  
   wire _roundIncr_near_even_T_1 ;  
   wire _roundIncr_near_even_T_3 ;  
   wire _roundIncr_near_even_T_4 ;  
   wire _roundIncr_near_even_T_5 ;  
   wire _roundIncr_near_even_T_8 ;  
   wire roundIncr_near_even ;  
   wire _roundIncr_near_maxMag_T_1 ;  
   wire roundIncr_near_maxMag ;  
   wire _roundIncr_T ;  
   wire _roundIncr_T_1 ;  
   wire _roundIncr_T_2 ;  
   wire _roundIncr_T_3 ;  
   wire _roundIncr_T_4 ;  
   wire _roundIncr_T_5 ;  
   wire _roundIncr_T_6 ;  
   wire _roundIncr_T_8 ;  
   wire _roundIncr_T_9 ;  
   wire roundIncr ;  
   wire [63:0] complUnroundedInt ;  
   wire _roundedInt_T ;  
   wire [63:0] _roundedInt_T_2 ;  
   wire [63:0] _roundedInt_T_3 ;  
   wire _roundedInt_T_4 ;  
   wire [63:0] _GEN_1 ;  
   wire [63:0] roundedInt ;  
   wire magGeOne_atOverflowEdge ;  
   wire _roundCarryBut2_T_1 ;  
   wire roundCarryBut2 ;  
   wire _common_overflow_T ;  
   wire _common_overflow_T_2 ;  
   wire _common_overflow_T_3 ;  
   wire _common_overflow_T_4 ;  
   wire _common_overflow_T_5 ;  
   wire _common_overflow_T_6 ;  
   wire _common_overflow_T_7 ;  
   wire _common_overflow_T_8 ;  
   wire _common_overflow_T_10 ;  
   wire _common_overflow_T_11 ;  
   wire _common_overflow_T_12 ;  
   wire _common_overflow_T_13 ;  
   wire _common_overflow_T_14 ;  
   wire _common_overflow_T_16 ;  
   wire _common_overflow_T_17 ;  
   wire common_overflow ;  
   wire invalidExc ;  
   wire overflow ;  
   wire _inexact_T_2 ;  
   wire inexact ;  
   wire excSign ;  
   wire _excOut_T ;  
   wire [63:0] _excOut_T_1 ;  
   wire [62:0] _excOut_T_3 ;  
   wire [63:0] _GEN_2 ;  
   wire [63:0] excOut ;  
   wire _io_out_T ;  
   wire [1:0] io_intExceptionFlags_hi ;  
   wire [29:0] RecFNToIN_covSum ;  
  assign rawIn_exp=io_in[63:52]; 
  assign rawIn_isZero=rawIn_exp[11:9]==3'h0; 
  assign rawIn_isSpecial=rawIn_exp[11:10]==2'h3; 
  assign rawIn__isNaN=rawIn_isSpecial&rawIn_exp[9]; 
  assign rawIn__isInf=rawIn_isSpecial&~rawIn_exp[9]; 
  assign rawIn__sign=io_in[64]; 
  assign rawIn__sExp={1'b0,$signed(rawIn_exp)}; 
  assign rawIn_out_sig_hi_lo=~rawIn_isZero; 
  assign rawIn_out_sig_lo=io_in[51:0]; 
  assign rawIn__sig={1'h0,rawIn_out_sig_hi_lo,rawIn_out_sig_lo}; 
  assign magGeOne=rawIn__sExp[11]; 
  assign posExp=rawIn__sExp[10:0]; 
  assign _magJustBelowOne_T_1=&posExp; 
  assign magJustBelowOne=~magGeOne&_magJustBelowOne_T_1; 
  assign roundingMode_near_even=io_roundingMode==3'h0; 
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign roundingMode_max=io_roundingMode==3'h3; 
  assign roundingMode_near_maxMag=io_roundingMode==3'h4; 
  assign roundingMode_odd=io_roundingMode==3'h6; 
  assign shiftedSig_lo=rawIn__sig[51:0]; 
  assign _shiftedSig_T={magGeOne,shiftedSig_lo}; 
  assign _shiftedSig_T_2=magGeOne ? rawIn__sExp[5:0]:6'h0; 
  assign _GEN_0={63'b0,_shiftedSig_T}; 
  assign shiftedSig=_GEN_0<<_shiftedSig_T_2; 
  assign alignedSig_hi=shiftedSig[115:51]; 
  assign alignedSig_lo=|shiftedSig[50:0]; 
  assign alignedSig={alignedSig_hi,alignedSig_lo}; 
  assign unroundedInt=alignedSig[65:2]; 
  assign _common_inexact_T_1=|alignedSig[1:0]; 
  assign common_inexact=magGeOne ? _common_inexact_T_1:rawIn_out_sig_hi_lo; 
  assign _roundIncr_near_even_T_1=&alignedSig[2:1]; 
  assign _roundIncr_near_even_T_3=&alignedSig[1:0]; 
  assign _roundIncr_near_even_T_4=_roundIncr_near_even_T_1|_roundIncr_near_even_T_3; 
  assign _roundIncr_near_even_T_5=magGeOne&_roundIncr_near_even_T_4; 
  assign _roundIncr_near_even_T_8=magJustBelowOne&_common_inexact_T_1; 
  assign roundIncr_near_even=_roundIncr_near_even_T_5|_roundIncr_near_even_T_8; 
  assign _roundIncr_near_maxMag_T_1=magGeOne&alignedSig[1]; 
  assign roundIncr_near_maxMag=_roundIncr_near_maxMag_T_1|magJustBelowOne; 
  assign _roundIncr_T=roundingMode_near_even&roundIncr_near_even; 
  assign _roundIncr_T_1=roundingMode_near_maxMag&roundIncr_near_maxMag; 
  assign _roundIncr_T_2=_roundIncr_T|_roundIncr_T_1; 
  assign _roundIncr_T_3=roundingMode_min|roundingMode_odd; 
  assign _roundIncr_T_4=rawIn__sign&common_inexact; 
  assign _roundIncr_T_5=_roundIncr_T_3&_roundIncr_T_4; 
  assign _roundIncr_T_6=_roundIncr_T_2|_roundIncr_T_5; 
  assign _roundIncr_T_8=~rawIn__sign&common_inexact; 
  assign _roundIncr_T_9=roundingMode_max&_roundIncr_T_8; 
  assign roundIncr=_roundIncr_T_6|_roundIncr_T_9; 
  assign complUnroundedInt=rawIn__sign ? ~unroundedInt:unroundedInt; 
  assign _roundedInt_T=roundIncr^rawIn__sign; 
  assign _roundedInt_T_2=complUnroundedInt+64'h1; 
  assign _roundedInt_T_3=_roundedInt_T ? _roundedInt_T_2:complUnroundedInt; 
  assign _roundedInt_T_4=roundingMode_odd&common_inexact; 
  assign _GEN_1={63'b0,_roundedInt_T_4}; 
  assign roundedInt=_roundedInt_T_3|_GEN_1; 
  assign magGeOne_atOverflowEdge=posExp==11'h3f; 
  assign _roundCarryBut2_T_1=&unroundedInt[61:0]; 
  assign roundCarryBut2=_roundCarryBut2_T_1&roundIncr; 
  assign _common_overflow_T=posExp>=11'h40; 
  assign _common_overflow_T_2=|unroundedInt[62:0]; 
  assign _common_overflow_T_3=_common_overflow_T_2|roundIncr; 
  assign _common_overflow_T_4=magGeOne_atOverflowEdge&_common_overflow_T_3; 
  assign _common_overflow_T_5=posExp==11'h3e; 
  assign _common_overflow_T_6=_common_overflow_T_5&roundCarryBut2; 
  assign _common_overflow_T_7=magGeOne_atOverflowEdge|_common_overflow_T_6; 
  assign _common_overflow_T_8=rawIn__sign ? _common_overflow_T_4:_common_overflow_T_7; 
  assign _common_overflow_T_10=magGeOne_atOverflowEdge&unroundedInt[62]; 
  assign _common_overflow_T_11=_common_overflow_T_10&roundCarryBut2; 
  assign _common_overflow_T_12=rawIn__sign|_common_overflow_T_11; 
  assign _common_overflow_T_13=io_signedOut ? _common_overflow_T_8:_common_overflow_T_12; 
  assign _common_overflow_T_14=_common_overflow_T|_common_overflow_T_13; 
  assign _common_overflow_T_16=~io_signedOut&rawIn__sign; 
  assign _common_overflow_T_17=_common_overflow_T_16&roundIncr; 
  assign common_overflow=magGeOne ? _common_overflow_T_14:_common_overflow_T_17; 
  assign invalidExc=rawIn__isNaN|rawIn__isInf; 
  assign overflow=~invalidExc&common_overflow; 
  assign _inexact_T_2=~invalidExc&~common_overflow; 
  assign inexact=_inexact_T_2&common_inexact; 
  assign excSign=~rawIn__isNaN&rawIn__sign; 
  assign _excOut_T=io_signedOut==excSign; 
  assign _excOut_T_1=_excOut_T ? 64'h8000000000000000:64'h0; 
  assign _excOut_T_3=excSign ? 63'h0:63'h7fffffffffffffff; 
  assign _GEN_2={1'b0,_excOut_T_3}; 
  assign excOut=_excOut_T_1|_GEN_2; 
  assign _io_out_T=invalidExc|common_overflow; 
  assign io_intExceptionFlags_hi={invalidExc,overflow}; 
  assign io_out=_io_out_T ? excOut:roundedInt; 
  assign io_intExceptionFlags={io_intExceptionFlags_hi,inexact}; 
  assign RecFNToIN_covSum=30'h0; 
  assign io_covSum=RecFNToIN_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module RecFNToIN_1 (
  input [64:0] io_in,
  input [2:0] io_roundingMode,
  input io_signedOut,
  output [2:0] io_intExceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [11:0] rawIn_exp ;  
   wire rawIn_isZero ;  
   wire rawIn_isSpecial ;  
   wire rawIn__isNaN ;  
   wire rawIn__isInf ;  
   wire rawIn__sign ;  
   wire [12:0] rawIn__sExp ;  
   wire rawIn_out_sig_hi_lo ;  
   wire [51:0] rawIn_out_sig_lo ;  
   wire [53:0] rawIn__sig ;  
   wire magGeOne ;  
   wire [10:0] posExp ;  
   wire _magJustBelowOne_T_1 ;  
   wire magJustBelowOne ;  
   wire roundingMode_near_even ;  
   wire roundingMode_min ;  
   wire roundingMode_max ;  
   wire roundingMode_near_maxMag ;  
   wire roundingMode_odd ;  
   wire [51:0] shiftedSig_lo ;  
   wire [52:0] _shiftedSig_T ;  
   wire [4:0] _shiftedSig_T_2 ;  
   wire [83:0] _GEN_0 ;  
   wire [83:0] shiftedSig ;  
   wire [32:0] alignedSig_hi ;  
   wire alignedSig_lo ;  
   wire [33:0] alignedSig ;  
   wire [31:0] unroundedInt ;  
   wire _common_inexact_T_1 ;  
   wire common_inexact ;  
   wire _roundIncr_near_even_T_1 ;  
   wire _roundIncr_near_even_T_3 ;  
   wire _roundIncr_near_even_T_4 ;  
   wire _roundIncr_near_even_T_5 ;  
   wire _roundIncr_near_even_T_8 ;  
   wire roundIncr_near_even ;  
   wire _roundIncr_near_maxMag_T_1 ;  
   wire roundIncr_near_maxMag ;  
   wire _roundIncr_T ;  
   wire _roundIncr_T_1 ;  
   wire _roundIncr_T_2 ;  
   wire _roundIncr_T_3 ;  
   wire _roundIncr_T_4 ;  
   wire _roundIncr_T_5 ;  
   wire _roundIncr_T_6 ;  
   wire _roundIncr_T_8 ;  
   wire _roundIncr_T_9 ;  
   wire roundIncr ;  
   wire magGeOne_atOverflowEdge ;  
   wire _roundCarryBut2_T_1 ;  
   wire roundCarryBut2 ;  
   wire _common_overflow_T ;  
   wire _common_overflow_T_2 ;  
   wire _common_overflow_T_3 ;  
   wire _common_overflow_T_4 ;  
   wire _common_overflow_T_5 ;  
   wire _common_overflow_T_6 ;  
   wire _common_overflow_T_7 ;  
   wire _common_overflow_T_8 ;  
   wire _common_overflow_T_10 ;  
   wire _common_overflow_T_11 ;  
   wire _common_overflow_T_12 ;  
   wire _common_overflow_T_13 ;  
   wire _common_overflow_T_14 ;  
   wire _common_overflow_T_16 ;  
   wire _common_overflow_T_17 ;  
   wire common_overflow ;  
   wire invalidExc ;  
   wire overflow ;  
   wire _inexact_T_2 ;  
   wire inexact ;  
   wire [1:0] io_intExceptionFlags_hi ;  
   wire [29:0] RecFNToIN_1_covSum ;  
  assign rawIn_exp=io_in[63:52]; 
  assign rawIn_isZero=rawIn_exp[11:9]==3'h0; 
  assign rawIn_isSpecial=rawIn_exp[11:10]==2'h3; 
  assign rawIn__isNaN=rawIn_isSpecial&rawIn_exp[9]; 
  assign rawIn__isInf=rawIn_isSpecial&~rawIn_exp[9]; 
  assign rawIn__sign=io_in[64]; 
  assign rawIn__sExp={1'b0,$signed(rawIn_exp)}; 
  assign rawIn_out_sig_hi_lo=~rawIn_isZero; 
  assign rawIn_out_sig_lo=io_in[51:0]; 
  assign rawIn__sig={1'h0,rawIn_out_sig_hi_lo,rawIn_out_sig_lo}; 
  assign magGeOne=rawIn__sExp[11]; 
  assign posExp=rawIn__sExp[10:0]; 
  assign _magJustBelowOne_T_1=&posExp; 
  assign magJustBelowOne=~magGeOne&_magJustBelowOne_T_1; 
  assign roundingMode_near_even=io_roundingMode==3'h0; 
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign roundingMode_max=io_roundingMode==3'h3; 
  assign roundingMode_near_maxMag=io_roundingMode==3'h4; 
  assign roundingMode_odd=io_roundingMode==3'h6; 
  assign shiftedSig_lo=rawIn__sig[51:0]; 
  assign _shiftedSig_T={magGeOne,shiftedSig_lo}; 
  assign _shiftedSig_T_2=magGeOne ? rawIn__sExp[4:0]:5'h0; 
  assign _GEN_0={31'b0,_shiftedSig_T}; 
  assign shiftedSig=_GEN_0<<_shiftedSig_T_2; 
  assign alignedSig_hi=shiftedSig[83:51]; 
  assign alignedSig_lo=|shiftedSig[50:0]; 
  assign alignedSig={alignedSig_hi,alignedSig_lo}; 
  assign unroundedInt=alignedSig[33:2]; 
  assign _common_inexact_T_1=|alignedSig[1:0]; 
  assign common_inexact=magGeOne ? _common_inexact_T_1:rawIn_out_sig_hi_lo; 
  assign _roundIncr_near_even_T_1=&alignedSig[2:1]; 
  assign _roundIncr_near_even_T_3=&alignedSig[1:0]; 
  assign _roundIncr_near_even_T_4=_roundIncr_near_even_T_1|_roundIncr_near_even_T_3; 
  assign _roundIncr_near_even_T_5=magGeOne&_roundIncr_near_even_T_4; 
  assign _roundIncr_near_even_T_8=magJustBelowOne&_common_inexact_T_1; 
  assign roundIncr_near_even=_roundIncr_near_even_T_5|_roundIncr_near_even_T_8; 
  assign _roundIncr_near_maxMag_T_1=magGeOne&alignedSig[1]; 
  assign roundIncr_near_maxMag=_roundIncr_near_maxMag_T_1|magJustBelowOne; 
  assign _roundIncr_T=roundingMode_near_even&roundIncr_near_even; 
  assign _roundIncr_T_1=roundingMode_near_maxMag&roundIncr_near_maxMag; 
  assign _roundIncr_T_2=_roundIncr_T|_roundIncr_T_1; 
  assign _roundIncr_T_3=roundingMode_min|roundingMode_odd; 
  assign _roundIncr_T_4=rawIn__sign&common_inexact; 
  assign _roundIncr_T_5=_roundIncr_T_3&_roundIncr_T_4; 
  assign _roundIncr_T_6=_roundIncr_T_2|_roundIncr_T_5; 
  assign _roundIncr_T_8=~rawIn__sign&common_inexact; 
  assign _roundIncr_T_9=roundingMode_max&_roundIncr_T_8; 
  assign roundIncr=_roundIncr_T_6|_roundIncr_T_9; 
  assign magGeOne_atOverflowEdge=posExp==11'h1f; 
  assign _roundCarryBut2_T_1=&unroundedInt[29:0]; 
  assign roundCarryBut2=_roundCarryBut2_T_1&roundIncr; 
  assign _common_overflow_T=posExp>=11'h20; 
  assign _common_overflow_T_2=|unroundedInt[30:0]; 
  assign _common_overflow_T_3=_common_overflow_T_2|roundIncr; 
  assign _common_overflow_T_4=magGeOne_atOverflowEdge&_common_overflow_T_3; 
  assign _common_overflow_T_5=posExp==11'h1e; 
  assign _common_overflow_T_6=_common_overflow_T_5&roundCarryBut2; 
  assign _common_overflow_T_7=magGeOne_atOverflowEdge|_common_overflow_T_6; 
  assign _common_overflow_T_8=rawIn__sign ? _common_overflow_T_4:_common_overflow_T_7; 
  assign _common_overflow_T_10=magGeOne_atOverflowEdge&unroundedInt[30]; 
  assign _common_overflow_T_11=_common_overflow_T_10&roundCarryBut2; 
  assign _common_overflow_T_12=rawIn__sign|_common_overflow_T_11; 
  assign _common_overflow_T_13=io_signedOut ? _common_overflow_T_8:_common_overflow_T_12; 
  assign _common_overflow_T_14=_common_overflow_T|_common_overflow_T_13; 
  assign _common_overflow_T_16=~io_signedOut&rawIn__sign; 
  assign _common_overflow_T_17=_common_overflow_T_16&roundIncr; 
  assign common_overflow=magGeOne ? _common_overflow_T_14:_common_overflow_T_17; 
  assign invalidExc=rawIn__isNaN|rawIn__isInf; 
  assign overflow=~invalidExc&common_overflow; 
  assign _inexact_T_2=~invalidExc&~common_overflow; 
  assign inexact=_inexact_T_2&common_inexact; 
  assign io_intExceptionFlags_hi={invalidExc,overflow}; 
  assign io_intExceptionFlags={io_intExceptionFlags_hi,inexact}; 
  assign RecFNToIN_1_covSum=30'h0; 
  assign io_covSum=RecFNToIN_1_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module INToRecFN (
  input io_signedIn,
  input [63:0] io_in,
  input [2:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundAnyRawFNToRecFN_io_in_isZero ;  
   wire roundAnyRawFNToRecFN_io_in_sign ;  
   wire [8:0] roundAnyRawFNToRecFN_io_in_sExp ;  
   wire [64:0] roundAnyRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundAnyRawFNToRecFN_io_roundingMode ;  
   wire [32:0] roundAnyRawFNToRecFN_io_out ;  
   wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundAnyRawFNToRecFN_io_covSum ;  
   wire roundAnyRawFNToRecFN_metaAssert ;  
   wire intAsRawFloat_sign ;  
   wire [63:0] _intAsRawFloat_absIn_T_1 ;  
   wire [63:0] intAsRawFloat_extAbsIn_lo ;  
   wire [127:0] _intAsRawFloat_extAbsIn_T ;  
   wire [63:0] intAsRawFloat_extAbsIn ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_64 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_65 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_66 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_67 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_68 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_69 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_70 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_71 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_72 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_73 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_74 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_75 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_76 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_77 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_78 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_79 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_80 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_81 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_82 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_83 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_84 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_85 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_86 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_87 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_88 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_89 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_90 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_91 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_92 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_93 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_94 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_95 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_96 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_97 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_98 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_99 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_100 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_101 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_102 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_103 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_104 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_105 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_106 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_107 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_108 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_109 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_110 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_111 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_112 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_113 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_114 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_115 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_116 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_117 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_118 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_119 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_120 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_121 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_122 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_123 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_124 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_125 ;  
   wire [5:0] intAsRawFloat_adjustedNormDist ;  
   wire [126:0] _GEN_0 ;  
   wire [126:0] _intAsRawFloat_sig_T ;  
   wire [63:0] intAsRawFloat_sig ;  
   wire [5:0] intAsRawFloat_out_sExp_lo ;  
   wire [7:0] _intAsRawFloat_out_sExp_T_1 ;  
   wire [29:0] INToRecFN_covSum ;  
   wire [29:0] roundAnyRawFNToRecFN_sum ;  
   wire roundAnyRawFNToRecFN_metaAssert_wire ;  
  RoundAnyRawFNToRecFN_1 roundAnyRawFNToRecFN(.io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),.io_in_sign(roundAnyRawFNToRecFN_io_in_sign),.io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),.io_in_sig(roundAnyRawFNToRecFN_io_in_sig),.io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),.io_out(roundAnyRawFNToRecFN_io_out),.io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),.io_covSum(roundAnyRawFNToRecFN_io_covSum),.metaAssert(roundAnyRawFNToRecFN_metaAssert)); 
  assign intAsRawFloat_sign=io_signedIn&io_in[63]; 
  assign _intAsRawFloat_absIn_T_1=64'h0-io_in; 
  assign intAsRawFloat_extAbsIn_lo=intAsRawFloat_sign ? _intAsRawFloat_absIn_T_1:io_in; 
  assign _intAsRawFloat_extAbsIn_T={64'h0,intAsRawFloat_extAbsIn_lo}; 
  assign intAsRawFloat_extAbsIn=_intAsRawFloat_extAbsIn_T[63:0]; 
  assign _intAsRawFloat_adjustedNormDist_T_64=intAsRawFloat_extAbsIn[1] ? 6'h3e:6'h3f; 
  assign _intAsRawFloat_adjustedNormDist_T_65=intAsRawFloat_extAbsIn[2] ? 6'h3d:_intAsRawFloat_adjustedNormDist_T_64; 
  assign _intAsRawFloat_adjustedNormDist_T_66=intAsRawFloat_extAbsIn[3] ? 6'h3c:_intAsRawFloat_adjustedNormDist_T_65; 
  assign _intAsRawFloat_adjustedNormDist_T_67=intAsRawFloat_extAbsIn[4] ? 6'h3b:_intAsRawFloat_adjustedNormDist_T_66; 
  assign _intAsRawFloat_adjustedNormDist_T_68=intAsRawFloat_extAbsIn[5] ? 6'h3a:_intAsRawFloat_adjustedNormDist_T_67; 
  assign _intAsRawFloat_adjustedNormDist_T_69=intAsRawFloat_extAbsIn[6] ? 6'h39:_intAsRawFloat_adjustedNormDist_T_68; 
  assign _intAsRawFloat_adjustedNormDist_T_70=intAsRawFloat_extAbsIn[7] ? 6'h38:_intAsRawFloat_adjustedNormDist_T_69; 
  assign _intAsRawFloat_adjustedNormDist_T_71=intAsRawFloat_extAbsIn[8] ? 6'h37:_intAsRawFloat_adjustedNormDist_T_70; 
  assign _intAsRawFloat_adjustedNormDist_T_72=intAsRawFloat_extAbsIn[9] ? 6'h36:_intAsRawFloat_adjustedNormDist_T_71; 
  assign _intAsRawFloat_adjustedNormDist_T_73=intAsRawFloat_extAbsIn[10] ? 6'h35:_intAsRawFloat_adjustedNormDist_T_72; 
  assign _intAsRawFloat_adjustedNormDist_T_74=intAsRawFloat_extAbsIn[11] ? 6'h34:_intAsRawFloat_adjustedNormDist_T_73; 
  assign _intAsRawFloat_adjustedNormDist_T_75=intAsRawFloat_extAbsIn[12] ? 6'h33:_intAsRawFloat_adjustedNormDist_T_74; 
  assign _intAsRawFloat_adjustedNormDist_T_76=intAsRawFloat_extAbsIn[13] ? 6'h32:_intAsRawFloat_adjustedNormDist_T_75; 
  assign _intAsRawFloat_adjustedNormDist_T_77=intAsRawFloat_extAbsIn[14] ? 6'h31:_intAsRawFloat_adjustedNormDist_T_76; 
  assign _intAsRawFloat_adjustedNormDist_T_78=intAsRawFloat_extAbsIn[15] ? 6'h30:_intAsRawFloat_adjustedNormDist_T_77; 
  assign _intAsRawFloat_adjustedNormDist_T_79=intAsRawFloat_extAbsIn[16] ? 6'h2f:_intAsRawFloat_adjustedNormDist_T_78; 
  assign _intAsRawFloat_adjustedNormDist_T_80=intAsRawFloat_extAbsIn[17] ? 6'h2e:_intAsRawFloat_adjustedNormDist_T_79; 
  assign _intAsRawFloat_adjustedNormDist_T_81=intAsRawFloat_extAbsIn[18] ? 6'h2d:_intAsRawFloat_adjustedNormDist_T_80; 
  assign _intAsRawFloat_adjustedNormDist_T_82=intAsRawFloat_extAbsIn[19] ? 6'h2c:_intAsRawFloat_adjustedNormDist_T_81; 
  assign _intAsRawFloat_adjustedNormDist_T_83=intAsRawFloat_extAbsIn[20] ? 6'h2b:_intAsRawFloat_adjustedNormDist_T_82; 
  assign _intAsRawFloat_adjustedNormDist_T_84=intAsRawFloat_extAbsIn[21] ? 6'h2a:_intAsRawFloat_adjustedNormDist_T_83; 
  assign _intAsRawFloat_adjustedNormDist_T_85=intAsRawFloat_extAbsIn[22] ? 6'h29:_intAsRawFloat_adjustedNormDist_T_84; 
  assign _intAsRawFloat_adjustedNormDist_T_86=intAsRawFloat_extAbsIn[23] ? 6'h28:_intAsRawFloat_adjustedNormDist_T_85; 
  assign _intAsRawFloat_adjustedNormDist_T_87=intAsRawFloat_extAbsIn[24] ? 6'h27:_intAsRawFloat_adjustedNormDist_T_86; 
  assign _intAsRawFloat_adjustedNormDist_T_88=intAsRawFloat_extAbsIn[25] ? 6'h26:_intAsRawFloat_adjustedNormDist_T_87; 
  assign _intAsRawFloat_adjustedNormDist_T_89=intAsRawFloat_extAbsIn[26] ? 6'h25:_intAsRawFloat_adjustedNormDist_T_88; 
  assign _intAsRawFloat_adjustedNormDist_T_90=intAsRawFloat_extAbsIn[27] ? 6'h24:_intAsRawFloat_adjustedNormDist_T_89; 
  assign _intAsRawFloat_adjustedNormDist_T_91=intAsRawFloat_extAbsIn[28] ? 6'h23:_intAsRawFloat_adjustedNormDist_T_90; 
  assign _intAsRawFloat_adjustedNormDist_T_92=intAsRawFloat_extAbsIn[29] ? 6'h22:_intAsRawFloat_adjustedNormDist_T_91; 
  assign _intAsRawFloat_adjustedNormDist_T_93=intAsRawFloat_extAbsIn[30] ? 6'h21:_intAsRawFloat_adjustedNormDist_T_92; 
  assign _intAsRawFloat_adjustedNormDist_T_94=intAsRawFloat_extAbsIn[31] ? 6'h20:_intAsRawFloat_adjustedNormDist_T_93; 
  assign _intAsRawFloat_adjustedNormDist_T_95=intAsRawFloat_extAbsIn[32] ? 6'h1f:_intAsRawFloat_adjustedNormDist_T_94; 
  assign _intAsRawFloat_adjustedNormDist_T_96=intAsRawFloat_extAbsIn[33] ? 6'h1e:_intAsRawFloat_adjustedNormDist_T_95; 
  assign _intAsRawFloat_adjustedNormDist_T_97=intAsRawFloat_extAbsIn[34] ? 6'h1d:_intAsRawFloat_adjustedNormDist_T_96; 
  assign _intAsRawFloat_adjustedNormDist_T_98=intAsRawFloat_extAbsIn[35] ? 6'h1c:_intAsRawFloat_adjustedNormDist_T_97; 
  assign _intAsRawFloat_adjustedNormDist_T_99=intAsRawFloat_extAbsIn[36] ? 6'h1b:_intAsRawFloat_adjustedNormDist_T_98; 
  assign _intAsRawFloat_adjustedNormDist_T_100=intAsRawFloat_extAbsIn[37] ? 6'h1a:_intAsRawFloat_adjustedNormDist_T_99; 
  assign _intAsRawFloat_adjustedNormDist_T_101=intAsRawFloat_extAbsIn[38] ? 6'h19:_intAsRawFloat_adjustedNormDist_T_100; 
  assign _intAsRawFloat_adjustedNormDist_T_102=intAsRawFloat_extAbsIn[39] ? 6'h18:_intAsRawFloat_adjustedNormDist_T_101; 
  assign _intAsRawFloat_adjustedNormDist_T_103=intAsRawFloat_extAbsIn[40] ? 6'h17:_intAsRawFloat_adjustedNormDist_T_102; 
  assign _intAsRawFloat_adjustedNormDist_T_104=intAsRawFloat_extAbsIn[41] ? 6'h16:_intAsRawFloat_adjustedNormDist_T_103; 
  assign _intAsRawFloat_adjustedNormDist_T_105=intAsRawFloat_extAbsIn[42] ? 6'h15:_intAsRawFloat_adjustedNormDist_T_104; 
  assign _intAsRawFloat_adjustedNormDist_T_106=intAsRawFloat_extAbsIn[43] ? 6'h14:_intAsRawFloat_adjustedNormDist_T_105; 
  assign _intAsRawFloat_adjustedNormDist_T_107=intAsRawFloat_extAbsIn[44] ? 6'h13:_intAsRawFloat_adjustedNormDist_T_106; 
  assign _intAsRawFloat_adjustedNormDist_T_108=intAsRawFloat_extAbsIn[45] ? 6'h12:_intAsRawFloat_adjustedNormDist_T_107; 
  assign _intAsRawFloat_adjustedNormDist_T_109=intAsRawFloat_extAbsIn[46] ? 6'h11:_intAsRawFloat_adjustedNormDist_T_108; 
  assign _intAsRawFloat_adjustedNormDist_T_110=intAsRawFloat_extAbsIn[47] ? 6'h10:_intAsRawFloat_adjustedNormDist_T_109; 
  assign _intAsRawFloat_adjustedNormDist_T_111=intAsRawFloat_extAbsIn[48] ? 6'hf:_intAsRawFloat_adjustedNormDist_T_110; 
  assign _intAsRawFloat_adjustedNormDist_T_112=intAsRawFloat_extAbsIn[49] ? 6'he:_intAsRawFloat_adjustedNormDist_T_111; 
  assign _intAsRawFloat_adjustedNormDist_T_113=intAsRawFloat_extAbsIn[50] ? 6'hd:_intAsRawFloat_adjustedNormDist_T_112; 
  assign _intAsRawFloat_adjustedNormDist_T_114=intAsRawFloat_extAbsIn[51] ? 6'hc:_intAsRawFloat_adjustedNormDist_T_113; 
  assign _intAsRawFloat_adjustedNormDist_T_115=intAsRawFloat_extAbsIn[52] ? 6'hb:_intAsRawFloat_adjustedNormDist_T_114; 
  assign _intAsRawFloat_adjustedNormDist_T_116=intAsRawFloat_extAbsIn[53] ? 6'ha:_intAsRawFloat_adjustedNormDist_T_115; 
  assign _intAsRawFloat_adjustedNormDist_T_117=intAsRawFloat_extAbsIn[54] ? 6'h9:_intAsRawFloat_adjustedNormDist_T_116; 
  assign _intAsRawFloat_adjustedNormDist_T_118=intAsRawFloat_extAbsIn[55] ? 6'h8:_intAsRawFloat_adjustedNormDist_T_117; 
  assign _intAsRawFloat_adjustedNormDist_T_119=intAsRawFloat_extAbsIn[56] ? 6'h7:_intAsRawFloat_adjustedNormDist_T_118; 
  assign _intAsRawFloat_adjustedNormDist_T_120=intAsRawFloat_extAbsIn[57] ? 6'h6:_intAsRawFloat_adjustedNormDist_T_119; 
  assign _intAsRawFloat_adjustedNormDist_T_121=intAsRawFloat_extAbsIn[58] ? 6'h5:_intAsRawFloat_adjustedNormDist_T_120; 
  assign _intAsRawFloat_adjustedNormDist_T_122=intAsRawFloat_extAbsIn[59] ? 6'h4:_intAsRawFloat_adjustedNormDist_T_121; 
  assign _intAsRawFloat_adjustedNormDist_T_123=intAsRawFloat_extAbsIn[60] ? 6'h3:_intAsRawFloat_adjustedNormDist_T_122; 
  assign _intAsRawFloat_adjustedNormDist_T_124=intAsRawFloat_extAbsIn[61] ? 6'h2:_intAsRawFloat_adjustedNormDist_T_123; 
  assign _intAsRawFloat_adjustedNormDist_T_125=intAsRawFloat_extAbsIn[62] ? 6'h1:_intAsRawFloat_adjustedNormDist_T_124; 
  assign intAsRawFloat_adjustedNormDist=intAsRawFloat_extAbsIn[63] ? 6'h0:_intAsRawFloat_adjustedNormDist_T_125; 
  assign _GEN_0={63'b0,intAsRawFloat_extAbsIn}; 
  assign _intAsRawFloat_sig_T=_GEN_0<<intAsRawFloat_adjustedNormDist; 
  assign intAsRawFloat_sig=_intAsRawFloat_sig_T[63:0]; 
  assign intAsRawFloat_out_sExp_lo=~intAsRawFloat_adjustedNormDist; 
  assign _intAsRawFloat_out_sExp_T_1={2'h2,intAsRawFloat_out_sExp_lo}; 
  assign io_out=roundAnyRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundAnyRawFNToRecFN_io_exceptionFlags; 
  assign roundAnyRawFNToRecFN_io_in_isZero=~intAsRawFloat_sig[63]; 
  assign roundAnyRawFNToRecFN_io_in_sign=io_signedIn&io_in[63]; 
  assign roundAnyRawFNToRecFN_io_in_sExp={1'b0,$signed(_intAsRawFloat_out_sExp_T_1)}; 
  assign roundAnyRawFNToRecFN_io_in_sig={1'b0,intAsRawFloat_sig}; 
  assign roundAnyRawFNToRecFN_io_roundingMode=io_roundingMode; 
  assign INToRecFN_covSum=30'h0; 
  assign roundAnyRawFNToRecFN_sum=INToRecFN_covSum+roundAnyRawFNToRecFN_io_covSum; 
  assign io_covSum=roundAnyRawFNToRecFN_sum; 
  assign roundAnyRawFNToRecFN_metaAssert_wire=roundAnyRawFNToRecFN_metaAssert; 
  assign metaAssert=roundAnyRawFNToRecFN_metaAssert_wire; 
endmodule
 
module INToRecFN_1 (
  input io_signedIn,
  input [63:0] io_in,
  input [2:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundAnyRawFNToRecFN_io_in_isZero ;  
   wire roundAnyRawFNToRecFN_io_in_sign ;  
   wire [8:0] roundAnyRawFNToRecFN_io_in_sExp ;  
   wire [64:0] roundAnyRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundAnyRawFNToRecFN_io_roundingMode ;  
   wire [64:0] roundAnyRawFNToRecFN_io_out ;  
   wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundAnyRawFNToRecFN_io_covSum ;  
   wire roundAnyRawFNToRecFN_metaAssert ;  
   wire intAsRawFloat_sign ;  
   wire [63:0] _intAsRawFloat_absIn_T_1 ;  
   wire [63:0] intAsRawFloat_extAbsIn_lo ;  
   wire [127:0] _intAsRawFloat_extAbsIn_T ;  
   wire [63:0] intAsRawFloat_extAbsIn ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_64 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_65 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_66 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_67 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_68 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_69 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_70 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_71 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_72 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_73 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_74 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_75 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_76 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_77 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_78 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_79 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_80 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_81 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_82 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_83 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_84 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_85 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_86 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_87 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_88 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_89 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_90 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_91 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_92 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_93 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_94 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_95 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_96 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_97 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_98 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_99 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_100 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_101 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_102 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_103 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_104 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_105 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_106 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_107 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_108 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_109 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_110 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_111 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_112 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_113 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_114 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_115 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_116 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_117 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_118 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_119 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_120 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_121 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_122 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_123 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_124 ;  
   wire [5:0] _intAsRawFloat_adjustedNormDist_T_125 ;  
   wire [5:0] intAsRawFloat_adjustedNormDist ;  
   wire [126:0] _GEN_0 ;  
   wire [126:0] _intAsRawFloat_sig_T ;  
   wire [63:0] intAsRawFloat_sig ;  
   wire [5:0] intAsRawFloat_out_sExp_lo ;  
   wire [7:0] _intAsRawFloat_out_sExp_T_1 ;  
   wire [29:0] INToRecFN_1_covSum ;  
   wire [29:0] roundAnyRawFNToRecFN_sum ;  
   wire roundAnyRawFNToRecFN_metaAssert_wire ;  
  RoundAnyRawFNToRecFN_2 roundAnyRawFNToRecFN(.io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),.io_in_sign(roundAnyRawFNToRecFN_io_in_sign),.io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),.io_in_sig(roundAnyRawFNToRecFN_io_in_sig),.io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),.io_out(roundAnyRawFNToRecFN_io_out),.io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),.io_covSum(roundAnyRawFNToRecFN_io_covSum),.metaAssert(roundAnyRawFNToRecFN_metaAssert)); 
  assign intAsRawFloat_sign=io_signedIn&io_in[63]; 
  assign _intAsRawFloat_absIn_T_1=64'h0-io_in; 
  assign intAsRawFloat_extAbsIn_lo=intAsRawFloat_sign ? _intAsRawFloat_absIn_T_1:io_in; 
  assign _intAsRawFloat_extAbsIn_T={64'h0,intAsRawFloat_extAbsIn_lo}; 
  assign intAsRawFloat_extAbsIn=_intAsRawFloat_extAbsIn_T[63:0]; 
  assign _intAsRawFloat_adjustedNormDist_T_64=intAsRawFloat_extAbsIn[1] ? 6'h3e:6'h3f; 
  assign _intAsRawFloat_adjustedNormDist_T_65=intAsRawFloat_extAbsIn[2] ? 6'h3d:_intAsRawFloat_adjustedNormDist_T_64; 
  assign _intAsRawFloat_adjustedNormDist_T_66=intAsRawFloat_extAbsIn[3] ? 6'h3c:_intAsRawFloat_adjustedNormDist_T_65; 
  assign _intAsRawFloat_adjustedNormDist_T_67=intAsRawFloat_extAbsIn[4] ? 6'h3b:_intAsRawFloat_adjustedNormDist_T_66; 
  assign _intAsRawFloat_adjustedNormDist_T_68=intAsRawFloat_extAbsIn[5] ? 6'h3a:_intAsRawFloat_adjustedNormDist_T_67; 
  assign _intAsRawFloat_adjustedNormDist_T_69=intAsRawFloat_extAbsIn[6] ? 6'h39:_intAsRawFloat_adjustedNormDist_T_68; 
  assign _intAsRawFloat_adjustedNormDist_T_70=intAsRawFloat_extAbsIn[7] ? 6'h38:_intAsRawFloat_adjustedNormDist_T_69; 
  assign _intAsRawFloat_adjustedNormDist_T_71=intAsRawFloat_extAbsIn[8] ? 6'h37:_intAsRawFloat_adjustedNormDist_T_70; 
  assign _intAsRawFloat_adjustedNormDist_T_72=intAsRawFloat_extAbsIn[9] ? 6'h36:_intAsRawFloat_adjustedNormDist_T_71; 
  assign _intAsRawFloat_adjustedNormDist_T_73=intAsRawFloat_extAbsIn[10] ? 6'h35:_intAsRawFloat_adjustedNormDist_T_72; 
  assign _intAsRawFloat_adjustedNormDist_T_74=intAsRawFloat_extAbsIn[11] ? 6'h34:_intAsRawFloat_adjustedNormDist_T_73; 
  assign _intAsRawFloat_adjustedNormDist_T_75=intAsRawFloat_extAbsIn[12] ? 6'h33:_intAsRawFloat_adjustedNormDist_T_74; 
  assign _intAsRawFloat_adjustedNormDist_T_76=intAsRawFloat_extAbsIn[13] ? 6'h32:_intAsRawFloat_adjustedNormDist_T_75; 
  assign _intAsRawFloat_adjustedNormDist_T_77=intAsRawFloat_extAbsIn[14] ? 6'h31:_intAsRawFloat_adjustedNormDist_T_76; 
  assign _intAsRawFloat_adjustedNormDist_T_78=intAsRawFloat_extAbsIn[15] ? 6'h30:_intAsRawFloat_adjustedNormDist_T_77; 
  assign _intAsRawFloat_adjustedNormDist_T_79=intAsRawFloat_extAbsIn[16] ? 6'h2f:_intAsRawFloat_adjustedNormDist_T_78; 
  assign _intAsRawFloat_adjustedNormDist_T_80=intAsRawFloat_extAbsIn[17] ? 6'h2e:_intAsRawFloat_adjustedNormDist_T_79; 
  assign _intAsRawFloat_adjustedNormDist_T_81=intAsRawFloat_extAbsIn[18] ? 6'h2d:_intAsRawFloat_adjustedNormDist_T_80; 
  assign _intAsRawFloat_adjustedNormDist_T_82=intAsRawFloat_extAbsIn[19] ? 6'h2c:_intAsRawFloat_adjustedNormDist_T_81; 
  assign _intAsRawFloat_adjustedNormDist_T_83=intAsRawFloat_extAbsIn[20] ? 6'h2b:_intAsRawFloat_adjustedNormDist_T_82; 
  assign _intAsRawFloat_adjustedNormDist_T_84=intAsRawFloat_extAbsIn[21] ? 6'h2a:_intAsRawFloat_adjustedNormDist_T_83; 
  assign _intAsRawFloat_adjustedNormDist_T_85=intAsRawFloat_extAbsIn[22] ? 6'h29:_intAsRawFloat_adjustedNormDist_T_84; 
  assign _intAsRawFloat_adjustedNormDist_T_86=intAsRawFloat_extAbsIn[23] ? 6'h28:_intAsRawFloat_adjustedNormDist_T_85; 
  assign _intAsRawFloat_adjustedNormDist_T_87=intAsRawFloat_extAbsIn[24] ? 6'h27:_intAsRawFloat_adjustedNormDist_T_86; 
  assign _intAsRawFloat_adjustedNormDist_T_88=intAsRawFloat_extAbsIn[25] ? 6'h26:_intAsRawFloat_adjustedNormDist_T_87; 
  assign _intAsRawFloat_adjustedNormDist_T_89=intAsRawFloat_extAbsIn[26] ? 6'h25:_intAsRawFloat_adjustedNormDist_T_88; 
  assign _intAsRawFloat_adjustedNormDist_T_90=intAsRawFloat_extAbsIn[27] ? 6'h24:_intAsRawFloat_adjustedNormDist_T_89; 
  assign _intAsRawFloat_adjustedNormDist_T_91=intAsRawFloat_extAbsIn[28] ? 6'h23:_intAsRawFloat_adjustedNormDist_T_90; 
  assign _intAsRawFloat_adjustedNormDist_T_92=intAsRawFloat_extAbsIn[29] ? 6'h22:_intAsRawFloat_adjustedNormDist_T_91; 
  assign _intAsRawFloat_adjustedNormDist_T_93=intAsRawFloat_extAbsIn[30] ? 6'h21:_intAsRawFloat_adjustedNormDist_T_92; 
  assign _intAsRawFloat_adjustedNormDist_T_94=intAsRawFloat_extAbsIn[31] ? 6'h20:_intAsRawFloat_adjustedNormDist_T_93; 
  assign _intAsRawFloat_adjustedNormDist_T_95=intAsRawFloat_extAbsIn[32] ? 6'h1f:_intAsRawFloat_adjustedNormDist_T_94; 
  assign _intAsRawFloat_adjustedNormDist_T_96=intAsRawFloat_extAbsIn[33] ? 6'h1e:_intAsRawFloat_adjustedNormDist_T_95; 
  assign _intAsRawFloat_adjustedNormDist_T_97=intAsRawFloat_extAbsIn[34] ? 6'h1d:_intAsRawFloat_adjustedNormDist_T_96; 
  assign _intAsRawFloat_adjustedNormDist_T_98=intAsRawFloat_extAbsIn[35] ? 6'h1c:_intAsRawFloat_adjustedNormDist_T_97; 
  assign _intAsRawFloat_adjustedNormDist_T_99=intAsRawFloat_extAbsIn[36] ? 6'h1b:_intAsRawFloat_adjustedNormDist_T_98; 
  assign _intAsRawFloat_adjustedNormDist_T_100=intAsRawFloat_extAbsIn[37] ? 6'h1a:_intAsRawFloat_adjustedNormDist_T_99; 
  assign _intAsRawFloat_adjustedNormDist_T_101=intAsRawFloat_extAbsIn[38] ? 6'h19:_intAsRawFloat_adjustedNormDist_T_100; 
  assign _intAsRawFloat_adjustedNormDist_T_102=intAsRawFloat_extAbsIn[39] ? 6'h18:_intAsRawFloat_adjustedNormDist_T_101; 
  assign _intAsRawFloat_adjustedNormDist_T_103=intAsRawFloat_extAbsIn[40] ? 6'h17:_intAsRawFloat_adjustedNormDist_T_102; 
  assign _intAsRawFloat_adjustedNormDist_T_104=intAsRawFloat_extAbsIn[41] ? 6'h16:_intAsRawFloat_adjustedNormDist_T_103; 
  assign _intAsRawFloat_adjustedNormDist_T_105=intAsRawFloat_extAbsIn[42] ? 6'h15:_intAsRawFloat_adjustedNormDist_T_104; 
  assign _intAsRawFloat_adjustedNormDist_T_106=intAsRawFloat_extAbsIn[43] ? 6'h14:_intAsRawFloat_adjustedNormDist_T_105; 
  assign _intAsRawFloat_adjustedNormDist_T_107=intAsRawFloat_extAbsIn[44] ? 6'h13:_intAsRawFloat_adjustedNormDist_T_106; 
  assign _intAsRawFloat_adjustedNormDist_T_108=intAsRawFloat_extAbsIn[45] ? 6'h12:_intAsRawFloat_adjustedNormDist_T_107; 
  assign _intAsRawFloat_adjustedNormDist_T_109=intAsRawFloat_extAbsIn[46] ? 6'h11:_intAsRawFloat_adjustedNormDist_T_108; 
  assign _intAsRawFloat_adjustedNormDist_T_110=intAsRawFloat_extAbsIn[47] ? 6'h10:_intAsRawFloat_adjustedNormDist_T_109; 
  assign _intAsRawFloat_adjustedNormDist_T_111=intAsRawFloat_extAbsIn[48] ? 6'hf:_intAsRawFloat_adjustedNormDist_T_110; 
  assign _intAsRawFloat_adjustedNormDist_T_112=intAsRawFloat_extAbsIn[49] ? 6'he:_intAsRawFloat_adjustedNormDist_T_111; 
  assign _intAsRawFloat_adjustedNormDist_T_113=intAsRawFloat_extAbsIn[50] ? 6'hd:_intAsRawFloat_adjustedNormDist_T_112; 
  assign _intAsRawFloat_adjustedNormDist_T_114=intAsRawFloat_extAbsIn[51] ? 6'hc:_intAsRawFloat_adjustedNormDist_T_113; 
  assign _intAsRawFloat_adjustedNormDist_T_115=intAsRawFloat_extAbsIn[52] ? 6'hb:_intAsRawFloat_adjustedNormDist_T_114; 
  assign _intAsRawFloat_adjustedNormDist_T_116=intAsRawFloat_extAbsIn[53] ? 6'ha:_intAsRawFloat_adjustedNormDist_T_115; 
  assign _intAsRawFloat_adjustedNormDist_T_117=intAsRawFloat_extAbsIn[54] ? 6'h9:_intAsRawFloat_adjustedNormDist_T_116; 
  assign _intAsRawFloat_adjustedNormDist_T_118=intAsRawFloat_extAbsIn[55] ? 6'h8:_intAsRawFloat_adjustedNormDist_T_117; 
  assign _intAsRawFloat_adjustedNormDist_T_119=intAsRawFloat_extAbsIn[56] ? 6'h7:_intAsRawFloat_adjustedNormDist_T_118; 
  assign _intAsRawFloat_adjustedNormDist_T_120=intAsRawFloat_extAbsIn[57] ? 6'h6:_intAsRawFloat_adjustedNormDist_T_119; 
  assign _intAsRawFloat_adjustedNormDist_T_121=intAsRawFloat_extAbsIn[58] ? 6'h5:_intAsRawFloat_adjustedNormDist_T_120; 
  assign _intAsRawFloat_adjustedNormDist_T_122=intAsRawFloat_extAbsIn[59] ? 6'h4:_intAsRawFloat_adjustedNormDist_T_121; 
  assign _intAsRawFloat_adjustedNormDist_T_123=intAsRawFloat_extAbsIn[60] ? 6'h3:_intAsRawFloat_adjustedNormDist_T_122; 
  assign _intAsRawFloat_adjustedNormDist_T_124=intAsRawFloat_extAbsIn[61] ? 6'h2:_intAsRawFloat_adjustedNormDist_T_123; 
  assign _intAsRawFloat_adjustedNormDist_T_125=intAsRawFloat_extAbsIn[62] ? 6'h1:_intAsRawFloat_adjustedNormDist_T_124; 
  assign intAsRawFloat_adjustedNormDist=intAsRawFloat_extAbsIn[63] ? 6'h0:_intAsRawFloat_adjustedNormDist_T_125; 
  assign _GEN_0={63'b0,intAsRawFloat_extAbsIn}; 
  assign _intAsRawFloat_sig_T=_GEN_0<<intAsRawFloat_adjustedNormDist; 
  assign intAsRawFloat_sig=_intAsRawFloat_sig_T[63:0]; 
  assign intAsRawFloat_out_sExp_lo=~intAsRawFloat_adjustedNormDist; 
  assign _intAsRawFloat_out_sExp_T_1={2'h2,intAsRawFloat_out_sExp_lo}; 
  assign io_out=roundAnyRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundAnyRawFNToRecFN_io_exceptionFlags; 
  assign roundAnyRawFNToRecFN_io_in_isZero=~intAsRawFloat_sig[63]; 
  assign roundAnyRawFNToRecFN_io_in_sign=io_signedIn&io_in[63]; 
  assign roundAnyRawFNToRecFN_io_in_sExp={1'b0,$signed(_intAsRawFloat_out_sExp_T_1)}; 
  assign roundAnyRawFNToRecFN_io_in_sig={1'b0,intAsRawFloat_sig}; 
  assign roundAnyRawFNToRecFN_io_roundingMode=io_roundingMode; 
  assign INToRecFN_1_covSum=30'h0; 
  assign roundAnyRawFNToRecFN_sum=INToRecFN_1_covSum+roundAnyRawFNToRecFN_io_covSum; 
  assign io_covSum=roundAnyRawFNToRecFN_sum; 
  assign roundAnyRawFNToRecFN_metaAssert_wire=roundAnyRawFNToRecFN_metaAssert; 
  assign metaAssert=roundAnyRawFNToRecFN_metaAssert_wire; 
endmodule
 
module RecFNToRecFN (
  input [64:0] io_in,
  input [2:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundAnyRawFNToRecFN_io_invalidExc ;  
   wire roundAnyRawFNToRecFN_io_in_isNaN ;  
   wire roundAnyRawFNToRecFN_io_in_isInf ;  
   wire roundAnyRawFNToRecFN_io_in_isZero ;  
   wire roundAnyRawFNToRecFN_io_in_sign ;  
   wire [12:0] roundAnyRawFNToRecFN_io_in_sExp ;  
   wire [53:0] roundAnyRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundAnyRawFNToRecFN_io_roundingMode ;  
   wire [32:0] roundAnyRawFNToRecFN_io_out ;  
   wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundAnyRawFNToRecFN_io_covSum ;  
   wire roundAnyRawFNToRecFN_metaAssert ;  
   wire [11:0] rawIn_exp ;  
   wire rawIn_isZero ;  
   wire rawIn_isSpecial ;  
   wire rawIn__isNaN ;  
   wire rawIn_out_sig_hi_lo ;  
   wire [51:0] rawIn_out_sig_lo ;  
   wire [1:0] rawIn_out_sig_hi ;  
   wire [53:0] rawIn__sig ;  
   wire [29:0] RecFNToRecFN_covSum ;  
   wire [29:0] roundAnyRawFNToRecFN_sum ;  
   wire roundAnyRawFNToRecFN_metaAssert_wire ;  
  RoundAnyRawFNToRecFN_3 roundAnyRawFNToRecFN(.io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),.io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),.io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),.io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),.io_in_sign(roundAnyRawFNToRecFN_io_in_sign),.io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),.io_in_sig(roundAnyRawFNToRecFN_io_in_sig),.io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),.io_out(roundAnyRawFNToRecFN_io_out),.io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),.io_covSum(roundAnyRawFNToRecFN_io_covSum),.metaAssert(roundAnyRawFNToRecFN_metaAssert)); 
  assign rawIn_exp=io_in[63:52]; 
  assign rawIn_isZero=rawIn_exp[11:9]==3'h0; 
  assign rawIn_isSpecial=rawIn_exp[11:10]==2'h3; 
  assign rawIn__isNaN=rawIn_isSpecial&rawIn_exp[9]; 
  assign rawIn_out_sig_hi_lo=~rawIn_isZero; 
  assign rawIn_out_sig_lo=io_in[51:0]; 
  assign rawIn_out_sig_hi={1'h0,rawIn_out_sig_hi_lo}; 
  assign rawIn__sig={1'h0,rawIn_out_sig_hi_lo,rawIn_out_sig_lo}; 
  assign io_out=roundAnyRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundAnyRawFNToRecFN_io_exceptionFlags; 
  assign roundAnyRawFNToRecFN_io_invalidExc=rawIn__isNaN&~rawIn__sig[51]; 
  assign roundAnyRawFNToRecFN_io_in_isNaN=rawIn_isSpecial&rawIn_exp[9]; 
  assign roundAnyRawFNToRecFN_io_in_isInf=rawIn_isSpecial&~rawIn_exp[9]; 
  assign roundAnyRawFNToRecFN_io_in_isZero=rawIn_exp[11:9]==3'h0; 
  assign roundAnyRawFNToRecFN_io_in_sign=io_in[64]; 
  assign roundAnyRawFNToRecFN_io_in_sExp={1'b0,$signed(rawIn_exp)}; 
  assign roundAnyRawFNToRecFN_io_in_sig={rawIn_out_sig_hi,rawIn_out_sig_lo}; 
  assign roundAnyRawFNToRecFN_io_roundingMode=io_roundingMode; 
  assign RecFNToRecFN_covSum=30'h0; 
  assign roundAnyRawFNToRecFN_sum=RecFNToRecFN_covSum+roundAnyRawFNToRecFN_io_covSum; 
  assign io_covSum=roundAnyRawFNToRecFN_sum; 
  assign roundAnyRawFNToRecFN_metaAssert_wire=roundAnyRawFNToRecFN_metaAssert; 
  assign metaAssert=roundAnyRawFNToRecFN_metaAssert_wire; 
endmodule
 
module MulAddRecFNPipe_1 (
  input clock,
  input reset,
  input io_validin,
  input [1:0] io_op,
  input [64:0] io_a,
  input [64:0] io_b,
  input [64:0] io_c,
  input [2:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output io_validout,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   wire [1:0] mulAddRecFNToRaw_preMul_io_op ;  
   wire [64:0] mulAddRecFNToRaw_preMul_io_a ;  
   wire [64:0] mulAddRecFNToRaw_preMul_io_b ;  
   wire [64:0] mulAddRecFNToRaw_preMul_io_c ;  
   wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddA ;  
   wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddB ;  
   wire [105:0] mulAddRecFNToRaw_preMul_io_mulAddC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfA ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfB ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_signProd ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC ;  
   wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant ;  
   wire [5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist ;  
   wire [54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC ;  
   wire mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC ;  
   wire [29:0] mulAddRecFNToRaw_preMul_io_covSum ;  
   wire mulAddRecFNToRaw_preMul_metaAssert ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_signProd ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC ;  
   wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant ;  
   wire [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist ;  
   wire [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC ;  
   wire mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC ;  
   wire [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult ;  
   wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode ;  
   wire mulAddRecFNToRaw_postMul_io_invalidExc ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_isNaN ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_isInf ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_isZero ;  
   wire mulAddRecFNToRaw_postMul_io_rawOut_sign ;  
   wire [12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp ;  
   wire [55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig ;  
   wire [29:0] mulAddRecFNToRaw_postMul_io_covSum ;  
   wire mulAddRecFNToRaw_postMul_metaAssert ;  
   wire roundRawFNToRecFN_io_invalidExc ;  
   wire roundRawFNToRecFN_io_infiniteExc ;  
   wire roundRawFNToRecFN_io_in_isNaN ;  
   wire roundRawFNToRecFN_io_in_isInf ;  
   wire roundRawFNToRecFN_io_in_isZero ;  
   wire roundRawFNToRecFN_io_in_sign ;  
   wire [12:0] roundRawFNToRecFN_io_in_sExp ;  
   wire [55:0] roundRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundRawFNToRecFN_io_roundingMode ;  
   wire roundRawFNToRecFN_io_detectTininess ;  
   wire [64:0] roundRawFNToRecFN_io_out ;  
   wire [4:0] roundRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundRawFNToRecFN_io_covSum ;  
   wire roundRawFNToRecFN_metaAssert ;  
   wire [105:0] _mulAddResult_T ;  
   wire [106:0] mulAddResult ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny ;  
   reg [31:0] _RAND_0 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB ;  
   reg [31:0] _RAND_1 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA ;  
   reg [31:0] _RAND_2 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA ;  
   reg [31:0] _RAND_3 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB ;  
   reg [31:0] _RAND_4 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB ;  
   reg [31:0] _RAND_5 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd ;  
   reg [31:0] _RAND_6 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC ;  
   reg [31:0] _RAND_7 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC ;  
   reg [31:0] _RAND_8 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC ;  
   reg [31:0] _RAND_9 ;  
   reg [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum ;  
   reg [31:0] _RAND_10 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags ;  
   reg [31:0] _RAND_11 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant ;  
   reg [31:0] _RAND_12 ;  
   reg [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist ;  
   reg [31:0] _RAND_13 ;  
   reg [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC ;  
   reg [63:0] _RAND_14 ;  
   reg mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC ;  
   reg [31:0] _RAND_15 ;  
   reg [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult_b ;  
   reg [127:0] _RAND_16 ;  
   reg [2:0] mulAddRecFNToRaw_postMul_io_roundingMode_b ;  
   reg [31:0] _RAND_17 ;  
   reg [2:0] roundingMode_stage0_b ;  
   reg [31:0] _RAND_18 ;  
   reg detectTininess_stage0_b ;  
   reg [31:0] _RAND_19 ;  
   reg valid_stage0_v ;  
   reg [31:0] _RAND_20 ;  
   reg roundRawFNToRecFN_io_invalidExc_b ;  
   reg [31:0] _RAND_21 ;  
   reg roundRawFNToRecFN_io_in_b_isNaN ;  
   reg [31:0] _RAND_22 ;  
   reg roundRawFNToRecFN_io_in_b_isInf ;  
   reg [31:0] _RAND_23 ;  
   reg roundRawFNToRecFN_io_in_b_isZero ;  
   reg [31:0] _RAND_24 ;  
   reg roundRawFNToRecFN_io_in_b_sign ;  
   reg [31:0] _RAND_25 ;  
   reg [12:0] roundRawFNToRecFN_io_in_b_sExp ;  
   reg [31:0] _RAND_26 ;  
   reg [55:0] roundRawFNToRecFN_io_in_b_sig ;  
   reg [63:0] _RAND_27 ;  
   reg [2:0] roundRawFNToRecFN_io_roundingMode_b ;  
   reg [31:0] _RAND_28 ;  
   reg roundRawFNToRecFN_io_detectTininess_b ;  
   reg [31:0] _RAND_29 ;  
   reg io_validout_v ;  
   reg [31:0] _RAND_30 ;  
   reg MulAddRecFNPipe_1_state ;  
   reg [31:0] _RAND_31 ;  
   reg MulAddRecFNPipe_1_cov[0:1] ;  
   reg [31:0] _RAND_32 ;  
   wire MulAddRecFNPipe_1_cov_read_data ;  
   wire MulAddRecFNPipe_1_cov_read_addr ;  
   wire MulAddRecFNPipe_1_cov_write_data ;  
   wire MulAddRecFNPipe_1_cov_write_addr ;  
   wire MulAddRecFNPipe_1_cov_write_mask ;  
   wire MulAddRecFNPipe_1_cov_write_en ;  
   reg [29:0] MulAddRecFNPipe_1_covSum ;  
   reg [31:0] _RAND_33 ;  
   wire valid_stage0_v_shl ;  
   wire valid_stage0_v_pad ;  
   wire [29:0] mulAddRecFNToRaw_preMul_sum ;  
   wire [29:0] mulAddRecFNToRaw_postMul_sum ;  
   wire [29:0] roundRawFNToRecFN_sum ;  
   wire mulAddRecFNToRaw_preMul_metaAssert_wire ;  
   wire mulAddRecFNToRaw_postMul_metaAssert_wire ;  
   wire roundRawFNToRecFN_metaAssert_wire ;  
   wire MulAddRecFNPipe_1_or2 ;  
   wire MulAddRecFNPipe_1_or0 ;  
   reg MulAddRecFNPipe_1_metaAssert ;  
   reg [31:0] _RAND_34 ;  
  MulAddRecFNToRaw_preMul_1 mulAddRecFNToRaw_preMul(.io_op(mulAddRecFNToRaw_preMul_io_op),.io_a(mulAddRecFNToRaw_preMul_io_a),.io_b(mulAddRecFNToRaw_preMul_io_b),.io_c(mulAddRecFNToRaw_preMul_io_c),.io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),.io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),.io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),.io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),.io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),.io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),.io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),.io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),.io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),.io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),.io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),.io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),.io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),.io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),.io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),.io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),.io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),.io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),.io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC),.io_covSum(mulAddRecFNToRaw_preMul_io_covSum),.metaAssert(mulAddRecFNToRaw_preMul_metaAssert)); 
  MulAddRecFNToRaw_postMul_1 mulAddRecFNToRaw_postMul(.io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),.io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),.io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),.io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),.io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),.io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),.io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),.io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),.io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),.io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),.io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),.io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),.io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),.io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),.io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),.io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),.io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),.io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),.io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),.io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),.io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),.io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),.io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),.io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),.io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig),.io_covSum(mulAddRecFNToRaw_postMul_io_covSum),.metaAssert(mulAddRecFNToRaw_postMul_metaAssert)); 
  RoundRawFNToRecFN_3 roundRawFNToRecFN(.io_invalidExc(roundRawFNToRecFN_io_invalidExc),.io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),.io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),.io_in_isInf(roundRawFNToRecFN_io_in_isInf),.io_in_isZero(roundRawFNToRecFN_io_in_isZero),.io_in_sign(roundRawFNToRecFN_io_in_sign),.io_in_sExp(roundRawFNToRecFN_io_in_sExp),.io_in_sig(roundRawFNToRecFN_io_in_sig),.io_roundingMode(roundRawFNToRecFN_io_roundingMode),.io_detectTininess(roundRawFNToRecFN_io_detectTininess),.io_out(roundRawFNToRecFN_io_out),.io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags),.io_covSum(roundRawFNToRecFN_io_covSum),.metaAssert(roundRawFNToRecFN_metaAssert)); 
  assign _mulAddResult_T=mulAddRecFNToRaw_preMul_io_mulAddA*mulAddRecFNToRaw_preMul_io_mulAddB; 
  assign mulAddResult=_mulAddResult_T+mulAddRecFNToRaw_preMul_io_mulAddC; 
  assign io_out=roundRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundRawFNToRecFN_io_exceptionFlags; 
  assign io_validout=io_validout_v; 
  assign mulAddRecFNToRaw_preMul_io_op=io_op; 
  assign mulAddRecFNToRaw_preMul_io_a=io_a; 
  assign mulAddRecFNToRaw_preMul_io_b=io_b; 
  assign mulAddRecFNToRaw_preMul_io_c=io_c; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd=mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum=mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags=mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant=mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist=mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC; 
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC=mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC; 
  assign mulAddRecFNToRaw_postMul_io_mulAddResult=mulAddRecFNToRaw_postMul_io_mulAddResult_b; 
  assign mulAddRecFNToRaw_postMul_io_roundingMode=mulAddRecFNToRaw_postMul_io_roundingMode_b; 
  assign roundRawFNToRecFN_io_invalidExc=roundRawFNToRecFN_io_invalidExc_b; 
  assign roundRawFNToRecFN_io_infiniteExc=1'h0; 
  assign roundRawFNToRecFN_io_in_isNaN=roundRawFNToRecFN_io_in_b_isNaN; 
  assign roundRawFNToRecFN_io_in_isInf=roundRawFNToRecFN_io_in_b_isInf; 
  assign roundRawFNToRecFN_io_in_isZero=roundRawFNToRecFN_io_in_b_isZero; 
  assign roundRawFNToRecFN_io_in_sign=roundRawFNToRecFN_io_in_b_sign; 
  assign roundRawFNToRecFN_io_in_sExp=roundRawFNToRecFN_io_in_b_sExp; 
  assign roundRawFNToRecFN_io_in_sig=roundRawFNToRecFN_io_in_b_sig; 
  assign roundRawFNToRecFN_io_roundingMode=roundRawFNToRecFN_io_roundingMode_b; 
  assign roundRawFNToRecFN_io_detectTininess=roundRawFNToRecFN_io_detectTininess_b; 
  assign MulAddRecFNPipe_1_cov_read_addr=MulAddRecFNPipe_1_state; 
  assign MulAddRecFNPipe_1_cov_read_data=MulAddRecFNPipe_1_cov[MulAddRecFNPipe_1_cov_read_addr]; 
  assign MulAddRecFNPipe_1_cov_write_data=1'h1; 
  assign MulAddRecFNPipe_1_cov_write_addr=MulAddRecFNPipe_1_state; 
  assign MulAddRecFNPipe_1_cov_write_mask=1'h1; 
  assign MulAddRecFNPipe_1_cov_write_en=1'h1; 
  assign valid_stage0_v_shl=valid_stage0_v; 
  assign valid_stage0_v_pad=valid_stage0_v_shl; 
  assign mulAddRecFNToRaw_preMul_sum=MulAddRecFNPipe_1_covSum+mulAddRecFNToRaw_preMul_io_covSum; 
  assign mulAddRecFNToRaw_postMul_sum=mulAddRecFNToRaw_preMul_sum+mulAddRecFNToRaw_postMul_io_covSum; 
  assign roundRawFNToRecFN_sum=mulAddRecFNToRaw_postMul_sum+roundRawFNToRecFN_io_covSum; 
  assign io_covSum=roundRawFNToRecFN_sum; 
  assign mulAddRecFNToRaw_preMul_metaAssert_wire=mulAddRecFNToRaw_preMul_metaAssert; 
  assign mulAddRecFNToRaw_postMul_metaAssert_wire=mulAddRecFNToRaw_postMul_metaAssert; 
  assign roundRawFNToRecFN_metaAssert_wire=roundRawFNToRecFN_metaAssert; 
  assign MulAddRecFNPipe_1_or2=mulAddRecFNToRaw_postMul_metaAssert_wire|roundRawFNToRecFN_metaAssert_wire; 
  assign MulAddRecFNPipe_1_or0=mulAddRecFNToRaw_preMul_metaAssert_wire|MulAddRecFNPipe_1_or2; 
  assign metaAssert=MulAddRecFNPipe_1_metaAssert; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isSigNaNAny <=mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNAOrB <=mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfA <=mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroA <=mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfB <=mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroB <=mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_signProd <=mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isNaNC <=mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isInfC <=mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_isZeroC <=mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <=13'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_sExpSum <=mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_doSubMags <=mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_CIsDominant <=mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <=6'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_CDom_CAlignDist <=mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <=55'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_highAlignedSigC <=mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <=1'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_fromPreMul_b_bit0AlignedSigC <=mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_mulAddResult_b <=107'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_mulAddResult_b <=mulAddResult;
               end 
         if (metaReset)
            begin 
              mulAddRecFNToRaw_postMul_io_roundingMode_b <=3'h0;
            end 
          else 
            if (io_validin)
               begin 
                 mulAddRecFNToRaw_postMul_io_roundingMode_b <=io_roundingMode;
               end 
         if (metaReset)
            begin 
              roundingMode_stage0_b <=3'h0;
            end 
          else 
            if (io_validin)
               begin 
                 roundingMode_stage0_b <=io_roundingMode;
               end 
         if (metaReset)
            begin 
              detectTininess_stage0_b <=1'h0;
            end 
          else 
            begin 
              detectTininess_stage0_b <=io_validin|detectTininess_stage0_b;
            end 
         if (metaReset)
            begin 
              valid_stage0_v <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 valid_stage0_v <=1'h0;
               end 
             else 
               begin 
                 valid_stage0_v <=io_validin;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_invalidExc_b <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_invalidExc_b <=mulAddRecFNToRaw_postMul_io_invalidExc;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_isNaN <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_isNaN <=mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_isInf <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_isInf <=mulAddRecFNToRaw_postMul_io_rawOut_isInf;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_isZero <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_isZero <=mulAddRecFNToRaw_postMul_io_rawOut_isZero;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_sign <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_sign <=mulAddRecFNToRaw_postMul_io_rawOut_sign;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_sExp <=13'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_sExp <=mulAddRecFNToRaw_postMul_io_rawOut_sExp;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_in_b_sig <=56'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_in_b_sig <=mulAddRecFNToRaw_postMul_io_rawOut_sig;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_roundingMode_b <=3'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_roundingMode_b <=roundingMode_stage0_b;
               end 
         if (metaReset)
            begin 
              roundRawFNToRecFN_io_detectTininess_b <=1'h0;
            end 
          else 
            if (valid_stage0_v)
               begin 
                 roundRawFNToRecFN_io_detectTininess_b <=detectTininess_stage0_b;
               end 
         if (metaReset)
            begin 
              io_validout_v <=1'h0;
            end 
          else 
            if (reset)
               begin 
                 io_validout_v <=1'h0;
               end 
             else 
               begin 
                 io_validout_v <=valid_stage0_v;
               end 
         MulAddRecFNPipe_1_state <=valid_stage0_v_pad;
         if (!(MulAddRecFNPipe_1_cov_read_data))
            begin 
              MulAddRecFNPipe_1_covSum <=MulAddRecFNPipe_1_covSum+1'h1;
            end 
         if (metaReset)
            begin 
              MulAddRecFNPipe_1_metaAssert <=1'h0;
            end 
          else 
            begin 
              MulAddRecFNPipe_1_metaAssert <=MulAddRecFNPipe_1_metaAssert|MulAddRecFNPipe_1_or0;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (MulAddRecFNPipe_1_cov_write_en&MulAddRecFNPipe_1_cov_write_mask)
            begin 
              MulAddRecFNPipe_1_cov [MulAddRecFNPipe_1_cov_write_addr]<=MulAddRecFNPipe_1_cov_write_data;
            end 
       end
  
endmodule
 
module DivSqrtRecFNToRaw_small (
  input clock,
  input reset,
  output io_inReady,
  input io_inValid,
  input io_sqrtOp,
  input [32:0] io_a,
  input [32:0] io_b,
  input [2:0] io_roundingMode,
  output io_rawOutValid_div,
  output io_rawOutValid_sqrt,
  output [2:0] io_roundingModeOut,
  output io_invalidExc,
  output io_infiniteExc,
  output io_rawOut_isNaN,
  output io_rawOut_isInf,
  output io_rawOut_isZero,
  output io_rawOut_sign,
  output [9:0] io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input divSqrtRawFN__halt) ; 
   wire divSqrtRawFN__clock ;  
   wire divSqrtRawFN__reset ;  
   wire divSqrtRawFN__io_inReady ;  
   wire divSqrtRawFN__io_inValid ;  
   wire divSqrtRawFN__io_sqrtOp ;  
   wire divSqrtRawFN__io_a_isNaN ;  
   wire divSqrtRawFN__io_a_isInf ;  
   wire divSqrtRawFN__io_a_isZero ;  
   wire divSqrtRawFN__io_a_sign ;  
   wire [9:0] divSqrtRawFN__io_a_sExp ;  
   wire [24:0] divSqrtRawFN__io_a_sig ;  
   wire divSqrtRawFN__io_b_isNaN ;  
   wire divSqrtRawFN__io_b_isInf ;  
   wire divSqrtRawFN__io_b_isZero ;  
   wire divSqrtRawFN__io_b_sign ;  
   wire [9:0] divSqrtRawFN__io_b_sExp ;  
   wire [24:0] divSqrtRawFN__io_b_sig ;  
   wire [2:0] divSqrtRawFN__io_roundingMode ;  
   wire divSqrtRawFN__io_rawOutValid_div ;  
   wire divSqrtRawFN__io_rawOutValid_sqrt ;  
   wire [2:0] divSqrtRawFN__io_roundingModeOut ;  
   wire divSqrtRawFN__io_invalidExc ;  
   wire divSqrtRawFN__io_infiniteExc ;  
   wire divSqrtRawFN__io_rawOut_isNaN ;  
   wire divSqrtRawFN__io_rawOut_isInf ;  
   wire divSqrtRawFN__io_rawOut_isZero ;  
   wire divSqrtRawFN__io_rawOut_sign ;  
   wire [9:0] divSqrtRawFN__io_rawOut_sExp ;  
   wire [26:0] divSqrtRawFN__io_rawOut_sig ;  
   wire [29:0] divSqrtRawFN__io_covSum ;  
   wire divSqrtRawFN__metaAssert ;  
   wire divSqrtRawFN__metaReset ;  
   wire [8:0] divSqrtRawFN_io_a_exp ;  
   wire divSqrtRawFN_io_a_isZero ;  
   wire divSqrtRawFN_io_a_isSpecial ;  
   wire divSqrtRawFN_io_a_out_sig_hi_lo ;  
   wire [22:0] divSqrtRawFN_io_a_out_sig_lo ;  
   wire [1:0] divSqrtRawFN_io_a_out_sig_hi ;  
   wire [8:0] divSqrtRawFN_io_b_exp ;  
   wire divSqrtRawFN_io_b_isZero ;  
   wire divSqrtRawFN_io_b_isSpecial ;  
   wire divSqrtRawFN_io_b_out_sig_hi_lo ;  
   wire [22:0] divSqrtRawFN_io_b_out_sig_lo ;  
   wire [1:0] divSqrtRawFN_io_b_out_sig_hi ;  
   wire [29:0] DivSqrtRecFNToRaw_small_covSum ;  
   wire [29:0] divSqrtRawFN__sum ;  
   wire divSqrtRawFN__metaAssert_wire ;  
   reg DivSqrtRecFNToRaw_small_metaAssert ;  
   reg [31:0] _RAND_0 ;  
  DivSqrtRawFN_small divSqrtRawFN_(.clock(divSqrtRawFN__clock),.reset(divSqrtRawFN__reset),.io_inReady(divSqrtRawFN__io_inReady),.io_inValid(divSqrtRawFN__io_inValid),.io_sqrtOp(divSqrtRawFN__io_sqrtOp),.io_a_isNaN(divSqrtRawFN__io_a_isNaN),.io_a_isInf(divSqrtRawFN__io_a_isInf),.io_a_isZero(divSqrtRawFN__io_a_isZero),.io_a_sign(divSqrtRawFN__io_a_sign),.io_a_sExp(divSqrtRawFN__io_a_sExp),.io_a_sig(divSqrtRawFN__io_a_sig),.io_b_isNaN(divSqrtRawFN__io_b_isNaN),.io_b_isInf(divSqrtRawFN__io_b_isInf),.io_b_isZero(divSqrtRawFN__io_b_isZero),.io_b_sign(divSqrtRawFN__io_b_sign),.io_b_sExp(divSqrtRawFN__io_b_sExp),.io_b_sig(divSqrtRawFN__io_b_sig),.io_roundingMode(divSqrtRawFN__io_roundingMode),.io_rawOutValid_div(divSqrtRawFN__io_rawOutValid_div),.io_rawOutValid_sqrt(divSqrtRawFN__io_rawOutValid_sqrt),.io_roundingModeOut(divSqrtRawFN__io_roundingModeOut),.io_invalidExc(divSqrtRawFN__io_invalidExc),.io_infiniteExc(divSqrtRawFN__io_infiniteExc),.io_rawOut_isNaN(divSqrtRawFN__io_rawOut_isNaN),.io_rawOut_isInf(divSqrtRawFN__io_rawOut_isInf),.io_rawOut_isZero(divSqrtRawFN__io_rawOut_isZero),.io_rawOut_sign(divSqrtRawFN__io_rawOut_sign),.io_rawOut_sExp(divSqrtRawFN__io_rawOut_sExp),.io_rawOut_sig(divSqrtRawFN__io_rawOut_sig),.io_covSum(divSqrtRawFN__io_covSum),.metaAssert(divSqrtRawFN__metaAssert),.metaReset(divSqrtRawFN__metaReset)); 
  assign divSqrtRawFN_io_a_exp=io_a[31:23]; 
  assign divSqrtRawFN_io_a_isZero=divSqrtRawFN_io_a_exp[8:6]==3'h0; 
  assign divSqrtRawFN_io_a_isSpecial=divSqrtRawFN_io_a_exp[8:7]==2'h3; 
  assign divSqrtRawFN_io_a_out_sig_hi_lo=~divSqrtRawFN_io_a_isZero; 
  assign divSqrtRawFN_io_a_out_sig_lo=io_a[22:0]; 
  assign divSqrtRawFN_io_a_out_sig_hi={1'h0,divSqrtRawFN_io_a_out_sig_hi_lo}; 
  assign divSqrtRawFN_io_b_exp=io_b[31:23]; 
  assign divSqrtRawFN_io_b_isZero=divSqrtRawFN_io_b_exp[8:6]==3'h0; 
  assign divSqrtRawFN_io_b_isSpecial=divSqrtRawFN_io_b_exp[8:7]==2'h3; 
  assign divSqrtRawFN_io_b_out_sig_hi_lo=~divSqrtRawFN_io_b_isZero; 
  assign divSqrtRawFN_io_b_out_sig_lo=io_b[22:0]; 
  assign divSqrtRawFN_io_b_out_sig_hi={1'h0,divSqrtRawFN_io_b_out_sig_hi_lo}; 
  assign io_inReady=divSqrtRawFN__io_inReady; 
  assign io_rawOutValid_div=divSqrtRawFN__io_rawOutValid_div; 
  assign io_rawOutValid_sqrt=divSqrtRawFN__io_rawOutValid_sqrt; 
  assign io_roundingModeOut=divSqrtRawFN__io_roundingModeOut; 
  assign io_invalidExc=divSqrtRawFN__io_invalidExc; 
  assign io_infiniteExc=divSqrtRawFN__io_infiniteExc; 
  assign io_rawOut_isNaN=divSqrtRawFN__io_rawOut_isNaN; 
  assign io_rawOut_isInf=divSqrtRawFN__io_rawOut_isInf; 
  assign io_rawOut_isZero=divSqrtRawFN__io_rawOut_isZero; 
  assign io_rawOut_sign=divSqrtRawFN__io_rawOut_sign; 
  assign io_rawOut_sExp=divSqrtRawFN__io_rawOut_sExp; 
  assign io_rawOut_sig=divSqrtRawFN__io_rawOut_sig; 
  assign divSqrtRawFN__clock=clock; 
  assign divSqrtRawFN__reset=reset; 
  assign divSqrtRawFN__io_inValid=io_inValid; 
  assign divSqrtRawFN__io_sqrtOp=io_sqrtOp; 
  assign divSqrtRawFN__io_a_isNaN=divSqrtRawFN_io_a_isSpecial&divSqrtRawFN_io_a_exp[6]; 
  assign divSqrtRawFN__io_a_isInf=divSqrtRawFN_io_a_isSpecial&~divSqrtRawFN_io_a_exp[6]; 
  assign divSqrtRawFN__io_a_isZero=divSqrtRawFN_io_a_exp[8:6]==3'h0; 
  assign divSqrtRawFN__io_a_sign=io_a[32]; 
  assign divSqrtRawFN__io_a_sExp={1'b0,$signed(divSqrtRawFN_io_a_exp)}; 
  assign divSqrtRawFN__io_a_sig={divSqrtRawFN_io_a_out_sig_hi,divSqrtRawFN_io_a_out_sig_lo}; 
  assign divSqrtRawFN__io_b_isNaN=divSqrtRawFN_io_b_isSpecial&divSqrtRawFN_io_b_exp[6]; 
  assign divSqrtRawFN__io_b_isInf=divSqrtRawFN_io_b_isSpecial&~divSqrtRawFN_io_b_exp[6]; 
  assign divSqrtRawFN__io_b_isZero=divSqrtRawFN_io_b_exp[8:6]==3'h0; 
  assign divSqrtRawFN__io_b_sign=io_b[32]; 
  assign divSqrtRawFN__io_b_sExp={1'b0,$signed(divSqrtRawFN_io_b_exp)}; 
  assign divSqrtRawFN__io_b_sig={divSqrtRawFN_io_b_out_sig_hi,divSqrtRawFN_io_b_out_sig_lo}; 
  assign divSqrtRawFN__io_roundingMode=io_roundingMode; 
  assign DivSqrtRecFNToRaw_small_covSum=30'h0; 
  assign divSqrtRawFN__sum=DivSqrtRecFNToRaw_small_covSum+divSqrtRawFN__io_covSum; 
  assign io_covSum=divSqrtRawFN__sum; 
  assign divSqrtRawFN__metaAssert_wire=divSqrtRawFN__metaAssert; 
  assign metaAssert=DivSqrtRecFNToRaw_small_metaAssert; 
  assign divSqrtRawFN__metaReset=metaReset|divSqrtRawFN__halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              DivSqrtRecFNToRaw_small_metaAssert <=1'h0;
            end 
          else 
            begin 
              DivSqrtRecFNToRaw_small_metaAssert <=DivSqrtRecFNToRaw_small_metaAssert|divSqrtRawFN__metaAssert_wire;
            end 
       end
  
endmodule
 
module RoundRawFNToRecFN_2 (
  input io_invalidExc,
  input io_infiniteExc,
  input io_in_isNaN,
  input io_in_isInf,
  input io_in_isZero,
  input io_in_sign,
  input [9:0] io_in_sExp,
  input [26:0] io_in_sig,
  input [2:0] io_roundingMode,
  input io_detectTininess,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundAnyRawFNToRecFN_io_invalidExc ;  
   wire roundAnyRawFNToRecFN_io_infiniteExc ;  
   wire roundAnyRawFNToRecFN_io_in_isNaN ;  
   wire roundAnyRawFNToRecFN_io_in_isInf ;  
   wire roundAnyRawFNToRecFN_io_in_isZero ;  
   wire roundAnyRawFNToRecFN_io_in_sign ;  
   wire [9:0] roundAnyRawFNToRecFN_io_in_sExp ;  
   wire [26:0] roundAnyRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundAnyRawFNToRecFN_io_roundingMode ;  
   wire roundAnyRawFNToRecFN_io_detectTininess ;  
   wire [32:0] roundAnyRawFNToRecFN_io_out ;  
   wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundAnyRawFNToRecFN_io_covSum ;  
   wire roundAnyRawFNToRecFN_metaAssert ;  
   wire [29:0] RoundRawFNToRecFN_2_covSum ;  
   wire [29:0] roundAnyRawFNToRecFN_sum ;  
   wire roundAnyRawFNToRecFN_metaAssert_wire ;  
  RoundAnyRawFNToRecFN_5 roundAnyRawFNToRecFN(.io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),.io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),.io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),.io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),.io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),.io_in_sign(roundAnyRawFNToRecFN_io_in_sign),.io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),.io_in_sig(roundAnyRawFNToRecFN_io_in_sig),.io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),.io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),.io_out(roundAnyRawFNToRecFN_io_out),.io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),.io_covSum(roundAnyRawFNToRecFN_io_covSum),.metaAssert(roundAnyRawFNToRecFN_metaAssert)); 
  assign io_out=roundAnyRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundAnyRawFNToRecFN_io_exceptionFlags; 
  assign roundAnyRawFNToRecFN_io_invalidExc=io_invalidExc; 
  assign roundAnyRawFNToRecFN_io_infiniteExc=io_infiniteExc; 
  assign roundAnyRawFNToRecFN_io_in_isNaN=io_in_isNaN; 
  assign roundAnyRawFNToRecFN_io_in_isInf=io_in_isInf; 
  assign roundAnyRawFNToRecFN_io_in_isZero=io_in_isZero; 
  assign roundAnyRawFNToRecFN_io_in_sign=io_in_sign; 
  assign roundAnyRawFNToRecFN_io_in_sExp=io_in_sExp; 
  assign roundAnyRawFNToRecFN_io_in_sig=io_in_sig; 
  assign roundAnyRawFNToRecFN_io_roundingMode=io_roundingMode; 
  assign roundAnyRawFNToRecFN_io_detectTininess=io_detectTininess; 
  assign RoundRawFNToRecFN_2_covSum=30'h0; 
  assign roundAnyRawFNToRecFN_sum=RoundRawFNToRecFN_2_covSum+roundAnyRawFNToRecFN_io_covSum; 
  assign io_covSum=roundAnyRawFNToRecFN_sum; 
  assign roundAnyRawFNToRecFN_metaAssert_wire=roundAnyRawFNToRecFN_metaAssert; 
  assign metaAssert=roundAnyRawFNToRecFN_metaAssert_wire; 
endmodule
 
module DivSqrtRecFNToRaw_small_1 (
  input clock,
  input reset,
  output io_inReady,
  input io_inValid,
  input io_sqrtOp,
  input [64:0] io_a,
  input [64:0] io_b,
  input [2:0] io_roundingMode,
  output io_rawOutValid_div,
  output io_rawOutValid_sqrt,
  output [2:0] io_roundingModeOut,
  output io_invalidExc,
  output io_infiniteExc,
  output io_rawOut_isNaN,
  output io_rawOut_isInf,
  output io_rawOut_isZero,
  output io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset,
  input divSqrtRawFN__halt) ; 
   wire divSqrtRawFN__clock ;  
   wire divSqrtRawFN__reset ;  
   wire divSqrtRawFN__io_inReady ;  
   wire divSqrtRawFN__io_inValid ;  
   wire divSqrtRawFN__io_sqrtOp ;  
   wire divSqrtRawFN__io_a_isNaN ;  
   wire divSqrtRawFN__io_a_isInf ;  
   wire divSqrtRawFN__io_a_isZero ;  
   wire divSqrtRawFN__io_a_sign ;  
   wire [12:0] divSqrtRawFN__io_a_sExp ;  
   wire [53:0] divSqrtRawFN__io_a_sig ;  
   wire divSqrtRawFN__io_b_isNaN ;  
   wire divSqrtRawFN__io_b_isInf ;  
   wire divSqrtRawFN__io_b_isZero ;  
   wire divSqrtRawFN__io_b_sign ;  
   wire [12:0] divSqrtRawFN__io_b_sExp ;  
   wire [53:0] divSqrtRawFN__io_b_sig ;  
   wire [2:0] divSqrtRawFN__io_roundingMode ;  
   wire divSqrtRawFN__io_rawOutValid_div ;  
   wire divSqrtRawFN__io_rawOutValid_sqrt ;  
   wire [2:0] divSqrtRawFN__io_roundingModeOut ;  
   wire divSqrtRawFN__io_invalidExc ;  
   wire divSqrtRawFN__io_infiniteExc ;  
   wire divSqrtRawFN__io_rawOut_isNaN ;  
   wire divSqrtRawFN__io_rawOut_isInf ;  
   wire divSqrtRawFN__io_rawOut_isZero ;  
   wire divSqrtRawFN__io_rawOut_sign ;  
   wire [12:0] divSqrtRawFN__io_rawOut_sExp ;  
   wire [55:0] divSqrtRawFN__io_rawOut_sig ;  
   wire [29:0] divSqrtRawFN__io_covSum ;  
   wire divSqrtRawFN__metaAssert ;  
   wire divSqrtRawFN__metaReset ;  
   wire [11:0] divSqrtRawFN_io_a_exp ;  
   wire divSqrtRawFN_io_a_isZero ;  
   wire divSqrtRawFN_io_a_isSpecial ;  
   wire divSqrtRawFN_io_a_out_sig_hi_lo ;  
   wire [51:0] divSqrtRawFN_io_a_out_sig_lo ;  
   wire [1:0] divSqrtRawFN_io_a_out_sig_hi ;  
   wire [11:0] divSqrtRawFN_io_b_exp ;  
   wire divSqrtRawFN_io_b_isZero ;  
   wire divSqrtRawFN_io_b_isSpecial ;  
   wire divSqrtRawFN_io_b_out_sig_hi_lo ;  
   wire [51:0] divSqrtRawFN_io_b_out_sig_lo ;  
   wire [1:0] divSqrtRawFN_io_b_out_sig_hi ;  
   wire [29:0] DivSqrtRecFNToRaw_small_1_covSum ;  
   wire [29:0] divSqrtRawFN__sum ;  
   wire divSqrtRawFN__metaAssert_wire ;  
   reg DivSqrtRecFNToRaw_small_1_metaAssert ;  
   reg [31:0] _RAND_0 ;  
  DivSqrtRawFN_small_1 divSqrtRawFN_(.clock(divSqrtRawFN__clock),.reset(divSqrtRawFN__reset),.io_inReady(divSqrtRawFN__io_inReady),.io_inValid(divSqrtRawFN__io_inValid),.io_sqrtOp(divSqrtRawFN__io_sqrtOp),.io_a_isNaN(divSqrtRawFN__io_a_isNaN),.io_a_isInf(divSqrtRawFN__io_a_isInf),.io_a_isZero(divSqrtRawFN__io_a_isZero),.io_a_sign(divSqrtRawFN__io_a_sign),.io_a_sExp(divSqrtRawFN__io_a_sExp),.io_a_sig(divSqrtRawFN__io_a_sig),.io_b_isNaN(divSqrtRawFN__io_b_isNaN),.io_b_isInf(divSqrtRawFN__io_b_isInf),.io_b_isZero(divSqrtRawFN__io_b_isZero),.io_b_sign(divSqrtRawFN__io_b_sign),.io_b_sExp(divSqrtRawFN__io_b_sExp),.io_b_sig(divSqrtRawFN__io_b_sig),.io_roundingMode(divSqrtRawFN__io_roundingMode),.io_rawOutValid_div(divSqrtRawFN__io_rawOutValid_div),.io_rawOutValid_sqrt(divSqrtRawFN__io_rawOutValid_sqrt),.io_roundingModeOut(divSqrtRawFN__io_roundingModeOut),.io_invalidExc(divSqrtRawFN__io_invalidExc),.io_infiniteExc(divSqrtRawFN__io_infiniteExc),.io_rawOut_isNaN(divSqrtRawFN__io_rawOut_isNaN),.io_rawOut_isInf(divSqrtRawFN__io_rawOut_isInf),.io_rawOut_isZero(divSqrtRawFN__io_rawOut_isZero),.io_rawOut_sign(divSqrtRawFN__io_rawOut_sign),.io_rawOut_sExp(divSqrtRawFN__io_rawOut_sExp),.io_rawOut_sig(divSqrtRawFN__io_rawOut_sig),.io_covSum(divSqrtRawFN__io_covSum),.metaAssert(divSqrtRawFN__metaAssert),.metaReset(divSqrtRawFN__metaReset)); 
  assign divSqrtRawFN_io_a_exp=io_a[63:52]; 
  assign divSqrtRawFN_io_a_isZero=divSqrtRawFN_io_a_exp[11:9]==3'h0; 
  assign divSqrtRawFN_io_a_isSpecial=divSqrtRawFN_io_a_exp[11:10]==2'h3; 
  assign divSqrtRawFN_io_a_out_sig_hi_lo=~divSqrtRawFN_io_a_isZero; 
  assign divSqrtRawFN_io_a_out_sig_lo=io_a[51:0]; 
  assign divSqrtRawFN_io_a_out_sig_hi={1'h0,divSqrtRawFN_io_a_out_sig_hi_lo}; 
  assign divSqrtRawFN_io_b_exp=io_b[63:52]; 
  assign divSqrtRawFN_io_b_isZero=divSqrtRawFN_io_b_exp[11:9]==3'h0; 
  assign divSqrtRawFN_io_b_isSpecial=divSqrtRawFN_io_b_exp[11:10]==2'h3; 
  assign divSqrtRawFN_io_b_out_sig_hi_lo=~divSqrtRawFN_io_b_isZero; 
  assign divSqrtRawFN_io_b_out_sig_lo=io_b[51:0]; 
  assign divSqrtRawFN_io_b_out_sig_hi={1'h0,divSqrtRawFN_io_b_out_sig_hi_lo}; 
  assign io_inReady=divSqrtRawFN__io_inReady; 
  assign io_rawOutValid_div=divSqrtRawFN__io_rawOutValid_div; 
  assign io_rawOutValid_sqrt=divSqrtRawFN__io_rawOutValid_sqrt; 
  assign io_roundingModeOut=divSqrtRawFN__io_roundingModeOut; 
  assign io_invalidExc=divSqrtRawFN__io_invalidExc; 
  assign io_infiniteExc=divSqrtRawFN__io_infiniteExc; 
  assign io_rawOut_isNaN=divSqrtRawFN__io_rawOut_isNaN; 
  assign io_rawOut_isInf=divSqrtRawFN__io_rawOut_isInf; 
  assign io_rawOut_isZero=divSqrtRawFN__io_rawOut_isZero; 
  assign io_rawOut_sign=divSqrtRawFN__io_rawOut_sign; 
  assign io_rawOut_sExp=divSqrtRawFN__io_rawOut_sExp; 
  assign io_rawOut_sig=divSqrtRawFN__io_rawOut_sig; 
  assign divSqrtRawFN__clock=clock; 
  assign divSqrtRawFN__reset=reset; 
  assign divSqrtRawFN__io_inValid=io_inValid; 
  assign divSqrtRawFN__io_sqrtOp=io_sqrtOp; 
  assign divSqrtRawFN__io_a_isNaN=divSqrtRawFN_io_a_isSpecial&divSqrtRawFN_io_a_exp[9]; 
  assign divSqrtRawFN__io_a_isInf=divSqrtRawFN_io_a_isSpecial&~divSqrtRawFN_io_a_exp[9]; 
  assign divSqrtRawFN__io_a_isZero=divSqrtRawFN_io_a_exp[11:9]==3'h0; 
  assign divSqrtRawFN__io_a_sign=io_a[64]; 
  assign divSqrtRawFN__io_a_sExp={1'b0,$signed(divSqrtRawFN_io_a_exp)}; 
  assign divSqrtRawFN__io_a_sig={divSqrtRawFN_io_a_out_sig_hi,divSqrtRawFN_io_a_out_sig_lo}; 
  assign divSqrtRawFN__io_b_isNaN=divSqrtRawFN_io_b_isSpecial&divSqrtRawFN_io_b_exp[9]; 
  assign divSqrtRawFN__io_b_isInf=divSqrtRawFN_io_b_isSpecial&~divSqrtRawFN_io_b_exp[9]; 
  assign divSqrtRawFN__io_b_isZero=divSqrtRawFN_io_b_exp[11:9]==3'h0; 
  assign divSqrtRawFN__io_b_sign=io_b[64]; 
  assign divSqrtRawFN__io_b_sExp={1'b0,$signed(divSqrtRawFN_io_b_exp)}; 
  assign divSqrtRawFN__io_b_sig={divSqrtRawFN_io_b_out_sig_hi,divSqrtRawFN_io_b_out_sig_lo}; 
  assign divSqrtRawFN__io_roundingMode=io_roundingMode; 
  assign DivSqrtRecFNToRaw_small_1_covSum=30'h0; 
  assign divSqrtRawFN__sum=DivSqrtRecFNToRaw_small_1_covSum+divSqrtRawFN__io_covSum; 
  assign io_covSum=divSqrtRawFN__sum; 
  assign divSqrtRawFN__metaAssert_wire=divSqrtRawFN__metaAssert; 
  assign metaAssert=DivSqrtRecFNToRaw_small_1_metaAssert; 
  assign divSqrtRawFN__metaReset=metaReset|divSqrtRawFN__halt; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              DivSqrtRecFNToRaw_small_1_metaAssert <=1'h0;
            end 
          else 
            begin 
              DivSqrtRecFNToRaw_small_1_metaAssert <=DivSqrtRecFNToRaw_small_1_metaAssert|divSqrtRawFN__metaAssert_wire;
            end 
       end
  
endmodule
 
module RoundRawFNToRecFN_3 (
  input io_invalidExc,
  input io_infiniteExc,
  input io_in_isNaN,
  input io_in_isInf,
  input io_in_isZero,
  input io_in_sign,
  input [12:0] io_in_sExp,
  input [55:0] io_in_sig,
  input [2:0] io_roundingMode,
  input io_detectTininess,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundAnyRawFNToRecFN_io_invalidExc ;  
   wire roundAnyRawFNToRecFN_io_infiniteExc ;  
   wire roundAnyRawFNToRecFN_io_in_isNaN ;  
   wire roundAnyRawFNToRecFN_io_in_isInf ;  
   wire roundAnyRawFNToRecFN_io_in_isZero ;  
   wire roundAnyRawFNToRecFN_io_in_sign ;  
   wire [12:0] roundAnyRawFNToRecFN_io_in_sExp ;  
   wire [55:0] roundAnyRawFNToRecFN_io_in_sig ;  
   wire [2:0] roundAnyRawFNToRecFN_io_roundingMode ;  
   wire roundAnyRawFNToRecFN_io_detectTininess ;  
   wire [64:0] roundAnyRawFNToRecFN_io_out ;  
   wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags ;  
   wire [29:0] roundAnyRawFNToRecFN_io_covSum ;  
   wire roundAnyRawFNToRecFN_metaAssert ;  
   wire [29:0] RoundRawFNToRecFN_3_covSum ;  
   wire [29:0] roundAnyRawFNToRecFN_sum ;  
   wire roundAnyRawFNToRecFN_metaAssert_wire ;  
  RoundAnyRawFNToRecFN_6 roundAnyRawFNToRecFN(.io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),.io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),.io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),.io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),.io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),.io_in_sign(roundAnyRawFNToRecFN_io_in_sign),.io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),.io_in_sig(roundAnyRawFNToRecFN_io_in_sig),.io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),.io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),.io_out(roundAnyRawFNToRecFN_io_out),.io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags),.io_covSum(roundAnyRawFNToRecFN_io_covSum),.metaAssert(roundAnyRawFNToRecFN_metaAssert)); 
  assign io_out=roundAnyRawFNToRecFN_io_out; 
  assign io_exceptionFlags=roundAnyRawFNToRecFN_io_exceptionFlags; 
  assign roundAnyRawFNToRecFN_io_invalidExc=io_invalidExc; 
  assign roundAnyRawFNToRecFN_io_infiniteExc=io_infiniteExc; 
  assign roundAnyRawFNToRecFN_io_in_isNaN=io_in_isNaN; 
  assign roundAnyRawFNToRecFN_io_in_isInf=io_in_isInf; 
  assign roundAnyRawFNToRecFN_io_in_isZero=io_in_isZero; 
  assign roundAnyRawFNToRecFN_io_in_sign=io_in_sign; 
  assign roundAnyRawFNToRecFN_io_in_sExp=io_in_sExp; 
  assign roundAnyRawFNToRecFN_io_in_sig=io_in_sig; 
  assign roundAnyRawFNToRecFN_io_roundingMode=io_roundingMode; 
  assign roundAnyRawFNToRecFN_io_detectTininess=io_detectTininess; 
  assign RoundRawFNToRecFN_3_covSum=30'h0; 
  assign roundAnyRawFNToRecFN_sum=RoundRawFNToRecFN_3_covSum+roundAnyRawFNToRecFN_io_covSum; 
  assign io_covSum=roundAnyRawFNToRecFN_sum; 
  assign roundAnyRawFNToRecFN_metaAssert_wire=roundAnyRawFNToRecFN_metaAssert; 
  assign metaAssert=roundAnyRawFNToRecFN_metaAssert_wire; 
endmodule
 
module RVCExpander (
  input [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0] io_out_rd,
  output [4:0] io_out_rs1,
  output [4:0] io_out_rs2,
  output [4:0] io_out_rs3,
  output io_rvc,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire _io_out_s_opc_T_1 ;  
   wire [6:0] io_out_s_lo_lo ;  
   wire [3:0] io_out_s_hi_hi_hi ;  
   wire [1:0] io_out_s_hi_hi_lo ;  
   wire io_out_s_hi_lo ;  
   wire io_out_s_lo_hi ;  
   wire [2:0] io_out_s_lo_1 ;  
   wire [4:0] io_out_s_lo_hi_1 ;  
   wire [29:0] _io_out_s_T ;  
   wire [4:0] io_out_s_0_rs3 ;  
   wire [1:0] io_out_s_hi_hi_2 ;  
   wire [2:0] io_out_s_hi_lo_1 ;  
   wire [7:0] io_out_s_hi_hi_hi_2 ;  
   wire [2:0] io_out_s_lo_5 ;  
   wire [4:0] io_out_s_hi_hi_lo_1 ;  
   wire [27:0] _io_out_s_T_4 ;  
   wire [6:0] io_out_s_hi_hi_hi_3 ;  
   wire [26:0] _io_out_s_T_9 ;  
   wire [27:0] _io_out_s_T_14 ;  
   wire [1:0] io_out_s_hi_hi_hi_5 ;  
   wire [4:0] io_out_s_lo_hi_lo ;  
   wire [26:0] _io_out_s_T_21 ;  
   wire [2:0] io_out_s_hi_hi_hi_6 ;  
   wire [4:0] io_out_s_lo_hi_lo_1 ;  
   wire [27:0] _io_out_s_T_28 ;  
   wire [26:0] _io_out_s_T_35 ;  
   wire [27:0] _io_out_s_T_42 ;  
   wire [6:0] io_out_s_hi_20 ;  
   wire [4:0] io_out_s_lo_52 ;  
   wire [11:0] io_out_s_hi_hi_hi_9 ;  
   wire [4:0] io_out_s_hi_hi_lo_8 ;  
   wire [31:0] io_out_s_8_bits ;  
   wire _io_out_s_opc_T_3 ;  
   wire [6:0] io_out_s_lo_lo_1 ;  
   wire [31:0] io_out_s_9_bits ;  
   wire [31:0] io_out_s_10_bits ;  
   wire _io_out_s_opc_T_7 ;  
   wire [6:0] io_out_s_me_lo ;  
   wire [14:0] io_out_s_me_hi_hi ;  
   wire [31:0] _io_out_s_me_T_2 ;  
   wire [19:0] io_out_s_me_hi_hi_1 ;  
   wire [31:0] io_out_s_me_bits ;  
   wire _io_out_s_T_68 ;  
   wire _io_out_s_T_70 ;  
   wire _io_out_s_T_71 ;  
   wire [6:0] io_out_s_lo_lo_2 ;  
   wire [2:0] io_out_s_hi_hi_hi_12 ;  
   wire [1:0] io_out_s_hi_hi_lo_10 ;  
   wire io_out_s_lo_hi_hi ;  
   wire [31:0] io_out_s_res_bits ;  
   wire [31:0] io_out_s_11_bits ;  
   wire [4:0] io_out_s_11_rd ;  
   wire [4:0] io_out_s_11_rs2 ;  
   wire [4:0] io_out_s_11_rs3 ;  
   wire [25:0] _io_out_s_T_79 ;  
   wire [30:0] _GEN_0 ;  
   wire [30:0] _io_out_s_T_81 ;  
   wire [31:0] _io_out_s_T_84 ;  
   wire [2:0] _io_out_s_funct_T ;  
   wire _io_out_s_funct_T_1 ;  
   wire [2:0] _io_out_s_funct_T_2 ;  
   wire _io_out_s_funct_T_3 ;  
   wire [2:0] _io_out_s_funct_T_4 ;  
   wire _io_out_s_funct_T_5 ;  
   wire [2:0] _io_out_s_funct_T_6 ;  
   wire _io_out_s_funct_T_7 ;  
   wire [2:0] _io_out_s_funct_T_8 ;  
   wire _io_out_s_funct_T_9 ;  
   wire [2:0] _io_out_s_funct_T_10 ;  
   wire _io_out_s_funct_T_11 ;  
   wire [2:0] _io_out_s_funct_T_12 ;  
   wire _io_out_s_funct_T_13 ;  
   wire [2:0] io_out_s_hi_lo_17 ;  
   wire _io_out_s_sub_T_1 ;  
   wire [30:0] io_out_s_sub ;  
   wire [6:0] io_out_s_lo_lo_3 ;  
   wire [24:0] _io_out_s_T_85 ;  
   wire [30:0] _GEN_1 ;  
   wire [30:0] _io_out_s_T_86 ;  
   wire _io_out_s_T_88 ;  
   wire [30:0] _io_out_s_T_89 ;  
   wire _io_out_s_T_90 ;  
   wire [31:0] _io_out_s_T_91 ;  
   wire _io_out_s_T_92 ;  
   wire [31:0] io_out_s_12_bits ;  
   wire [9:0] io_out_s_hi_hi_hi_hi ;  
   wire io_out_s_hi_hi_hi_lo ;  
   wire [1:0] io_out_s_hi_hi_lo_16 ;  
   wire io_out_s_hi_lo_lo ;  
   wire io_out_s_lo_hi_lo_5 ;  
   wire [2:0] io_out_s_lo_lo_hi ;  
   wire [20:0] _io_out_s_T_100 ;  
   wire io_out_s_hi_hi_hi_19 ;  
   wire [9:0] io_out_s_hi_hi_lo_18 ;  
   wire io_out_s_hi_lo_21 ;  
   wire [7:0] io_out_s_lo_hi_hi_5 ;  
   wire [31:0] io_out_s_13_bits ;  
   wire [4:0] io_out_s_hi_hi_hi_23 ;  
   wire [12:0] _io_out_s_T_116 ;  
   wire io_out_s_hi_hi_hi_24 ;  
   wire [5:0] io_out_s_hi_hi_lo_23 ;  
   wire [3:0] io_out_s_lo_hi_lo_12 ;  
   wire io_out_s_lo_lo_hi_4 ;  
   wire [31:0] io_out_s_14_bits ;  
   wire [31:0] io_out_s_15_bits ;  
   wire [6:0] io_out_s_lo_lo_10 ;  
   wire [25:0] _io_out_s_T_145 ;  
   wire [28:0] _io_out_s_T_150 ;  
   wire [1:0] io_out_s_hi_hi_47 ;  
   wire [2:0] io_out_s_lo_hi_41 ;  
   wire [27:0] _io_out_s_T_154 ;  
   wire [28:0] _io_out_s_T_158 ;  
   wire [24:0] _io_out_s_mv_T ;  
   wire [24:0] _io_out_s_add_T ;  
   wire [24:0] io_out_s_jr ;  
   wire [17:0] io_out_s_reserved_hi ;  
   wire [24:0] io_out_s_reserved ;  
   wire [24:0] _io_out_s_jr_reserved_T_2 ;  
   wire _io_out_s_jr_mv_T_1 ;  
   wire [31:0] io_out_s_mv_bits ;  
   wire [31:0] io_out_s_jr_reserved_bits ;  
   wire [31:0] io_out_s_jr_mv_bits ;  
   wire [4:0] io_out_s_jr_mv_rd ;  
   wire [4:0] io_out_s_jr_mv_rs1 ;  
   wire [4:0] io_out_s_jr_mv_rs2 ;  
   wire [4:0] io_out_s_jr_mv_rs3 ;  
   wire [24:0] io_out_s_jalr ;  
   wire [24:0] _io_out_s_ebreak_T ;  
   wire [24:0] io_out_s_ebreak ;  
   wire [24:0] _io_out_s_jalr_ebreak_T_2 ;  
   wire [31:0] io_out_s_add_bits ;  
   wire [31:0] io_out_s_jalr_ebreak_bits ;  
   wire [31:0] io_out_s_jalr_add_bits ;  
   wire [4:0] io_out_s_jalr_add_rd ;  
   wire [4:0] io_out_s_jalr_add_rs1 ;  
   wire [31:0] io_out_s_20_bits ;  
   wire [4:0] io_out_s_20_rd ;  
   wire [4:0] io_out_s_20_rs1 ;  
   wire [4:0] io_out_s_20_rs2 ;  
   wire [4:0] io_out_s_20_rs3 ;  
   wire [8:0] _io_out_s_T_163 ;  
   wire [3:0] io_out_s_hi_hi_hi_37 ;  
   wire [4:0] io_out_s_lo_hi_lo_19 ;  
   wire [28:0] _io_out_s_T_165 ;  
   wire [1:0] io_out_s_hi_hi_54 ;  
   wire [3:0] io_out_s_hi_lo_38 ;  
   wire [7:0] _io_out_s_T_169 ;  
   wire [2:0] io_out_s_hi_hi_hi_38 ;  
   wire [4:0] io_out_s_lo_hi_lo_20 ;  
   wire [27:0] _io_out_s_T_171 ;  
   wire [28:0] _io_out_s_T_177 ;  
   wire [4:0] io_out_s_24_rs1 ;  
   wire [4:0] io_out_s_24_rs2 ;  
   wire [2:0] io_out_lo ;  
   wire [4:0] _io_out_T ;  
   wire _io_out_T_1 ;  
   wire [31:0] io_out_s_1_bits ;  
   wire [31:0] io_out_s_0_bits ;  
   wire [31:0] _io_out_T_2_bits ;  
   wire [4:0] _io_out_T_2_rd ;  
   wire [4:0] _io_out_T_2_rs1 ;  
   wire [4:0] _io_out_T_2_rs3 ;  
   wire _io_out_T_3 ;  
   wire [31:0] io_out_s_2_bits ;  
   wire [31:0] _io_out_T_4_bits ;  
   wire [4:0] _io_out_T_4_rd ;  
   wire [4:0] _io_out_T_4_rs1 ;  
   wire [4:0] _io_out_T_4_rs3 ;  
   wire _io_out_T_5 ;  
   wire [31:0] io_out_s_3_bits ;  
   wire [31:0] _io_out_T_6_bits ;  
   wire [4:0] _io_out_T_6_rd ;  
   wire [4:0] _io_out_T_6_rs1 ;  
   wire [4:0] _io_out_T_6_rs3 ;  
   wire _io_out_T_7 ;  
   wire [31:0] io_out_s_4_bits ;  
   wire [31:0] _io_out_T_8_bits ;  
   wire [4:0] _io_out_T_8_rd ;  
   wire [4:0] _io_out_T_8_rs1 ;  
   wire [4:0] _io_out_T_8_rs3 ;  
   wire _io_out_T_9 ;  
   wire [31:0] io_out_s_5_bits ;  
   wire [31:0] _io_out_T_10_bits ;  
   wire [4:0] _io_out_T_10_rd ;  
   wire [4:0] _io_out_T_10_rs1 ;  
   wire [4:0] _io_out_T_10_rs3 ;  
   wire _io_out_T_11 ;  
   wire [31:0] io_out_s_6_bits ;  
   wire [31:0] _io_out_T_12_bits ;  
   wire [4:0] _io_out_T_12_rd ;  
   wire [4:0] _io_out_T_12_rs1 ;  
   wire [4:0] _io_out_T_12_rs3 ;  
   wire _io_out_T_13 ;  
   wire [31:0] io_out_s_7_bits ;  
   wire [31:0] _io_out_T_14_bits ;  
   wire [4:0] _io_out_T_14_rd ;  
   wire [4:0] _io_out_T_14_rs1 ;  
   wire [4:0] _io_out_T_14_rs3 ;  
   wire _io_out_T_15 ;  
   wire [31:0] _io_out_T_16_bits ;  
   wire [4:0] _io_out_T_16_rd ;  
   wire [4:0] _io_out_T_16_rs1 ;  
   wire [4:0] _io_out_T_16_rs2 ;  
   wire [4:0] _io_out_T_16_rs3 ;  
   wire _io_out_T_17 ;  
   wire [31:0] _io_out_T_18_bits ;  
   wire [4:0] _io_out_T_18_rd ;  
   wire [4:0] _io_out_T_18_rs1 ;  
   wire [4:0] _io_out_T_18_rs2 ;  
   wire [4:0] _io_out_T_18_rs3 ;  
   wire _io_out_T_19 ;  
   wire [31:0] _io_out_T_20_bits ;  
   wire [4:0] _io_out_T_20_rd ;  
   wire [4:0] _io_out_T_20_rs1 ;  
   wire [4:0] _io_out_T_20_rs2 ;  
   wire [4:0] _io_out_T_20_rs3 ;  
   wire _io_out_T_21 ;  
   wire [31:0] _io_out_T_22_bits ;  
   wire [4:0] _io_out_T_22_rd ;  
   wire [4:0] _io_out_T_22_rs1 ;  
   wire [4:0] _io_out_T_22_rs2 ;  
   wire [4:0] _io_out_T_22_rs3 ;  
   wire _io_out_T_23 ;  
   wire [31:0] _io_out_T_24_bits ;  
   wire [4:0] _io_out_T_24_rd ;  
   wire [4:0] _io_out_T_24_rs1 ;  
   wire [4:0] _io_out_T_24_rs2 ;  
   wire [4:0] _io_out_T_24_rs3 ;  
   wire _io_out_T_25 ;  
   wire [31:0] _io_out_T_26_bits ;  
   wire [4:0] _io_out_T_26_rd ;  
   wire [4:0] _io_out_T_26_rs1 ;  
   wire [4:0] _io_out_T_26_rs2 ;  
   wire [4:0] _io_out_T_26_rs3 ;  
   wire _io_out_T_27 ;  
   wire [31:0] _io_out_T_28_bits ;  
   wire [4:0] _io_out_T_28_rd ;  
   wire [4:0] _io_out_T_28_rs1 ;  
   wire [4:0] _io_out_T_28_rs2 ;  
   wire [4:0] _io_out_T_28_rs3 ;  
   wire _io_out_T_29 ;  
   wire [31:0] _io_out_T_30_bits ;  
   wire [4:0] _io_out_T_30_rd ;  
   wire [4:0] _io_out_T_30_rs1 ;  
   wire [4:0] _io_out_T_30_rs2 ;  
   wire [4:0] _io_out_T_30_rs3 ;  
   wire _io_out_T_31 ;  
   wire [31:0] io_out_s_16_bits ;  
   wire [31:0] _io_out_T_32_bits ;  
   wire [4:0] _io_out_T_32_rd ;  
   wire [4:0] _io_out_T_32_rs1 ;  
   wire [4:0] _io_out_T_32_rs2 ;  
   wire [4:0] _io_out_T_32_rs3 ;  
   wire _io_out_T_33 ;  
   wire [31:0] io_out_s_17_bits ;  
   wire [31:0] _io_out_T_34_bits ;  
   wire [4:0] _io_out_T_34_rd ;  
   wire [4:0] _io_out_T_34_rs1 ;  
   wire [4:0] _io_out_T_34_rs2 ;  
   wire [4:0] _io_out_T_34_rs3 ;  
   wire _io_out_T_35 ;  
   wire [31:0] io_out_s_18_bits ;  
   wire [31:0] _io_out_T_36_bits ;  
   wire [4:0] _io_out_T_36_rd ;  
   wire [4:0] _io_out_T_36_rs1 ;  
   wire [4:0] _io_out_T_36_rs2 ;  
   wire [4:0] _io_out_T_36_rs3 ;  
   wire _io_out_T_37 ;  
   wire [31:0] io_out_s_19_bits ;  
   wire [31:0] _io_out_T_38_bits ;  
   wire [4:0] _io_out_T_38_rd ;  
   wire [4:0] _io_out_T_38_rs1 ;  
   wire [4:0] _io_out_T_38_rs2 ;  
   wire [4:0] _io_out_T_38_rs3 ;  
   wire _io_out_T_39 ;  
   wire [31:0] _io_out_T_40_bits ;  
   wire [4:0] _io_out_T_40_rd ;  
   wire [4:0] _io_out_T_40_rs1 ;  
   wire [4:0] _io_out_T_40_rs2 ;  
   wire [4:0] _io_out_T_40_rs3 ;  
   wire _io_out_T_41 ;  
   wire [31:0] io_out_s_21_bits ;  
   wire [31:0] _io_out_T_42_bits ;  
   wire [4:0] _io_out_T_42_rd ;  
   wire [4:0] _io_out_T_42_rs1 ;  
   wire [4:0] _io_out_T_42_rs2 ;  
   wire [4:0] _io_out_T_42_rs3 ;  
   wire _io_out_T_43 ;  
   wire [31:0] io_out_s_22_bits ;  
   wire [31:0] _io_out_T_44_bits ;  
   wire [4:0] _io_out_T_44_rd ;  
   wire [4:0] _io_out_T_44_rs1 ;  
   wire [4:0] _io_out_T_44_rs2 ;  
   wire [4:0] _io_out_T_44_rs3 ;  
   wire _io_out_T_45 ;  
   wire [31:0] io_out_s_23_bits ;  
   wire [31:0] _io_out_T_46_bits ;  
   wire [4:0] _io_out_T_46_rd ;  
   wire [4:0] _io_out_T_46_rs1 ;  
   wire [4:0] _io_out_T_46_rs2 ;  
   wire [4:0] _io_out_T_46_rs3 ;  
   wire _io_out_T_47 ;  
   wire [31:0] _io_out_T_48_bits ;  
   wire [4:0] _io_out_T_48_rd ;  
   wire [4:0] _io_out_T_48_rs1 ;  
   wire [4:0] _io_out_T_48_rs2 ;  
   wire [4:0] _io_out_T_48_rs3 ;  
   wire _io_out_T_49 ;  
   wire [31:0] _io_out_T_50_bits ;  
   wire [4:0] _io_out_T_50_rd ;  
   wire [4:0] _io_out_T_50_rs1 ;  
   wire [4:0] _io_out_T_50_rs2 ;  
   wire [4:0] _io_out_T_50_rs3 ;  
   wire _io_out_T_51 ;  
   wire [31:0] _io_out_T_52_bits ;  
   wire [4:0] _io_out_T_52_rd ;  
   wire [4:0] _io_out_T_52_rs1 ;  
   wire [4:0] _io_out_T_52_rs2 ;  
   wire [4:0] _io_out_T_52_rs3 ;  
   wire _io_out_T_53 ;  
   wire [31:0] _io_out_T_54_bits ;  
   wire [4:0] _io_out_T_54_rd ;  
   wire [4:0] _io_out_T_54_rs1 ;  
   wire [4:0] _io_out_T_54_rs2 ;  
   wire [4:0] _io_out_T_54_rs3 ;  
   wire _io_out_T_55 ;  
   wire [31:0] _io_out_T_56_bits ;  
   wire [4:0] _io_out_T_56_rd ;  
   wire [4:0] _io_out_T_56_rs1 ;  
   wire [4:0] _io_out_T_56_rs2 ;  
   wire [4:0] _io_out_T_56_rs3 ;  
   wire _io_out_T_57 ;  
   wire [31:0] _io_out_T_58_bits ;  
   wire [4:0] _io_out_T_58_rd ;  
   wire [4:0] _io_out_T_58_rs1 ;  
   wire [4:0] _io_out_T_58_rs2 ;  
   wire [4:0] _io_out_T_58_rs3 ;  
   wire _io_out_T_59 ;  
   wire [31:0] _io_out_T_60_bits ;  
   wire [4:0] _io_out_T_60_rd ;  
   wire [4:0] _io_out_T_60_rs1 ;  
   wire [4:0] _io_out_T_60_rs2 ;  
   wire [4:0] _io_out_T_60_rs3 ;  
   wire _io_out_T_61 ;  
   wire [29:0] RVCExpander_covSum ;  
  assign _io_out_s_opc_T_1=|io_in[12:5]; 
  assign io_out_s_lo_lo=_io_out_s_opc_T_1 ? 7'h13:7'h1f; 
  assign io_out_s_hi_hi_hi=io_in[10:7]; 
  assign io_out_s_hi_hi_lo=io_in[12:11]; 
  assign io_out_s_hi_lo=io_in[5]; 
  assign io_out_s_lo_hi=io_in[6]; 
  assign io_out_s_lo_1=io_in[4:2]; 
  assign io_out_s_lo_hi_1={2'h1,io_out_s_lo_1}; 
  assign _io_out_s_T={io_out_s_hi_hi_hi,io_out_s_hi_hi_lo,io_out_s_hi_lo,io_out_s_lo_hi,2'h0,5'h2,3'h0,2'h1,io_out_s_lo_1,io_out_s_lo_lo}; 
  assign io_out_s_0_rs3=io_in[31:27]; 
  assign io_out_s_hi_hi_2=io_in[6:5]; 
  assign io_out_s_hi_lo_1=io_in[12:10]; 
  assign io_out_s_hi_hi_hi_2={io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0}; 
  assign io_out_s_lo_5=io_in[9:7]; 
  assign io_out_s_hi_hi_lo_1={2'h1,io_out_s_lo_5}; 
  assign _io_out_s_T_4={io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0,2'h1,io_out_s_lo_5,3'h3,2'h1,io_out_s_lo_1,7'h7}; 
  assign io_out_s_hi_hi_hi_3={io_out_s_hi_lo,io_out_s_hi_lo_1,io_out_s_lo_hi,2'h0}; 
  assign _io_out_s_T_9={io_out_s_hi_lo,io_out_s_hi_lo_1,io_out_s_lo_hi,2'h0,2'h1,io_out_s_lo_5,3'h2,2'h1,io_out_s_lo_1,7'h3}; 
  assign _io_out_s_T_14={io_out_s_hi_hi_2,io_out_s_hi_lo_1,3'h0,2'h1,io_out_s_lo_5,3'h3,2'h1,io_out_s_lo_1,7'h3}; 
  assign io_out_s_hi_hi_hi_5=io_out_s_hi_hi_hi_3[6:5]; 
  assign io_out_s_lo_hi_lo=io_out_s_hi_hi_hi_3[4:0]; 
  assign _io_out_s_T_21={io_out_s_hi_hi_hi_5,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h2,io_out_s_lo_hi_lo,7'h3f}; 
  assign io_out_s_hi_hi_hi_6=io_out_s_hi_hi_hi_2[7:5]; 
  assign io_out_s_lo_hi_lo_1=io_out_s_hi_hi_hi_2[4:0]; 
  assign _io_out_s_T_28={io_out_s_hi_hi_hi_6,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h3,io_out_s_lo_hi_lo_1,7'h27}; 
  assign _io_out_s_T_35={io_out_s_hi_hi_hi_5,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h2,io_out_s_lo_hi_lo,7'h23}; 
  assign _io_out_s_T_42={io_out_s_hi_hi_hi_6,2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,3'h3,io_out_s_lo_hi_lo_1,7'h23}; 
  assign io_out_s_hi_20=io_in[12] ? 7'h7f:7'h0; 
  assign io_out_s_lo_52=io_in[6:2]; 
  assign io_out_s_hi_hi_hi_9={io_out_s_hi_20,io_out_s_lo_52}; 
  assign io_out_s_hi_hi_lo_8=io_in[11:7]; 
  assign io_out_s_8_bits={io_out_s_hi_20,io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,7'h13}; 
  assign _io_out_s_opc_T_3=|io_out_s_hi_hi_lo_8; 
  assign io_out_s_lo_lo_1=_io_out_s_opc_T_3 ? 7'h1b:7'h1f; 
  assign io_out_s_9_bits={io_out_s_hi_20,io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_1}; 
  assign io_out_s_10_bits={io_out_s_hi_20,io_out_s_lo_52,5'h0,3'h0,io_out_s_hi_hi_lo_8,7'h13}; 
  assign _io_out_s_opc_T_7=|io_out_s_hi_hi_hi_9; 
  assign io_out_s_me_lo=_io_out_s_opc_T_7 ? 7'h37:7'h3f; 
  assign io_out_s_me_hi_hi=io_in[12] ? 15'h7fff:15'h0; 
  assign _io_out_s_me_T_2={io_out_s_me_hi_hi,io_out_s_lo_52,12'h0}; 
  assign io_out_s_me_hi_hi_1=_io_out_s_me_T_2[31:12]; 
  assign io_out_s_me_bits={io_out_s_me_hi_hi_1,io_out_s_hi_hi_lo_8,io_out_s_me_lo}; 
  assign _io_out_s_T_68=io_out_s_hi_hi_lo_8==5'h0; 
  assign _io_out_s_T_70=io_out_s_hi_hi_lo_8==5'h2; 
  assign _io_out_s_T_71=_io_out_s_T_68|_io_out_s_T_70; 
  assign io_out_s_lo_lo_2=_io_out_s_opc_T_7 ? 7'h13:7'h1f; 
  assign io_out_s_hi_hi_hi_12=io_in[12] ? 3'h7:3'h0; 
  assign io_out_s_hi_hi_lo_10=io_in[4:3]; 
  assign io_out_s_lo_hi_hi=io_in[2]; 
  assign io_out_s_res_bits={io_out_s_hi_hi_hi_12,io_out_s_hi_hi_lo_10,io_out_s_hi_lo,io_out_s_lo_hi_hi,io_out_s_lo_hi,4'h0,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_2}; 
  assign io_out_s_11_bits=_io_out_s_T_71 ? io_out_s_res_bits:io_out_s_me_bits; 
  assign io_out_s_11_rd=_io_out_s_T_71 ? io_out_s_hi_hi_lo_8:io_out_s_hi_hi_lo_8; 
  assign io_out_s_11_rs2=_io_out_s_T_71 ? io_out_s_lo_hi_1:io_out_s_lo_hi_1; 
  assign io_out_s_11_rs3=_io_out_s_T_71 ? io_out_s_0_rs3:io_out_s_0_rs3; 
  assign _io_out_s_T_79={io_in[12],io_out_s_lo_52,2'h1,io_out_s_lo_5,3'h5,2'h1,io_out_s_lo_5,7'h13}; 
  assign _GEN_0={5'b0,_io_out_s_T_79}; 
  assign _io_out_s_T_81=_GEN_0|31'h40000000; 
  assign _io_out_s_T_84={io_out_s_hi_20,io_out_s_lo_52,2'h1,io_out_s_lo_5,3'h7,2'h1,io_out_s_lo_5,7'h13}; 
  assign _io_out_s_funct_T={io_in[12],io_out_s_hi_hi_2}; 
  assign _io_out_s_funct_T_1=_io_out_s_funct_T==3'h1; 
  assign _io_out_s_funct_T_2=_io_out_s_funct_T_1 ? 3'h4:3'h0; 
  assign _io_out_s_funct_T_3=_io_out_s_funct_T==3'h2; 
  assign _io_out_s_funct_T_4=_io_out_s_funct_T_3 ? 3'h6:_io_out_s_funct_T_2; 
  assign _io_out_s_funct_T_5=_io_out_s_funct_T==3'h3; 
  assign _io_out_s_funct_T_6=_io_out_s_funct_T_5 ? 3'h7:_io_out_s_funct_T_4; 
  assign _io_out_s_funct_T_7=_io_out_s_funct_T==3'h4; 
  assign _io_out_s_funct_T_8=_io_out_s_funct_T_7 ? 3'h0:_io_out_s_funct_T_6; 
  assign _io_out_s_funct_T_9=_io_out_s_funct_T==3'h5; 
  assign _io_out_s_funct_T_10=_io_out_s_funct_T_9 ? 3'h0:_io_out_s_funct_T_8; 
  assign _io_out_s_funct_T_11=_io_out_s_funct_T==3'h6; 
  assign _io_out_s_funct_T_12=_io_out_s_funct_T_11 ? 3'h2:_io_out_s_funct_T_10; 
  assign _io_out_s_funct_T_13=_io_out_s_funct_T==3'h7; 
  assign io_out_s_hi_lo_17=_io_out_s_funct_T_13 ? 3'h3:_io_out_s_funct_T_12; 
  assign _io_out_s_sub_T_1=io_out_s_hi_hi_2==2'h0; 
  assign io_out_s_sub=_io_out_s_sub_T_1 ? 31'h40000000:31'h0; 
  assign io_out_s_lo_lo_3=io_in[12] ? 7'h3b:7'h33; 
  assign _io_out_s_T_85={2'h1,io_out_s_lo_1,2'h1,io_out_s_lo_5,io_out_s_hi_lo_17,2'h1,io_out_s_lo_5,io_out_s_lo_lo_3}; 
  assign _GEN_1={6'b0,_io_out_s_T_85}; 
  assign _io_out_s_T_86=_GEN_1|io_out_s_sub; 
  assign _io_out_s_T_88=io_in[11:10]==2'h1; 
  assign _io_out_s_T_89=_io_out_s_T_88 ? _io_out_s_T_81:{5'b0,_io_out_s_T_79}; 
  assign _io_out_s_T_90=io_in[11:10]==2'h2; 
  assign _io_out_s_T_91=_io_out_s_T_90 ? _io_out_s_T_84:{1'b0,_io_out_s_T_89}; 
  assign _io_out_s_T_92=io_in[11:10]==2'h3; 
  assign io_out_s_12_bits=_io_out_s_T_92 ? {1'b0,_io_out_s_T_86}:_io_out_s_T_91; 
  assign io_out_s_hi_hi_hi_hi=io_in[12] ? 10'h3ff:10'h0; 
  assign io_out_s_hi_hi_hi_lo=io_in[8]; 
  assign io_out_s_hi_hi_lo_16=io_in[10:9]; 
  assign io_out_s_hi_lo_lo=io_in[7]; 
  assign io_out_s_lo_hi_lo_5=io_in[11]; 
  assign io_out_s_lo_lo_hi=io_in[5:3]; 
  assign _io_out_s_T_100={io_out_s_hi_hi_hi_hi,io_out_s_hi_hi_hi_lo,io_out_s_hi_hi_lo_16,io_out_s_lo_hi,io_out_s_hi_lo_lo,io_out_s_lo_hi_hi,io_out_s_lo_hi_lo_5,io_out_s_lo_lo_hi,1'h0}; 
  assign io_out_s_hi_hi_hi_19=_io_out_s_T_100[20]; 
  assign io_out_s_hi_hi_lo_18=_io_out_s_T_100[10:1]; 
  assign io_out_s_hi_lo_21=_io_out_s_T_100[11]; 
  assign io_out_s_lo_hi_hi_5=_io_out_s_T_100[19:12]; 
  assign io_out_s_13_bits={io_out_s_hi_hi_hi_19,io_out_s_hi_hi_lo_18,io_out_s_hi_lo_21,io_out_s_lo_hi_hi_5,5'h0,7'h6f}; 
  assign io_out_s_hi_hi_hi_23=io_in[12] ? 5'h1f:5'h0; 
  assign _io_out_s_T_116={io_out_s_hi_hi_hi_23,io_out_s_hi_hi_2,io_out_s_lo_hi_hi,io_in[11:10],io_out_s_hi_hi_lo_10,1'h0}; 
  assign io_out_s_hi_hi_hi_24=_io_out_s_T_116[12]; 
  assign io_out_s_hi_hi_lo_23=_io_out_s_T_116[10:5]; 
  assign io_out_s_lo_hi_lo_12=_io_out_s_T_116[4:1]; 
  assign io_out_s_lo_lo_hi_4=_io_out_s_T_116[11]; 
  assign io_out_s_14_bits={io_out_s_hi_hi_hi_24,io_out_s_hi_hi_lo_23,5'h0,2'h1,io_out_s_lo_5,3'h0,io_out_s_lo_hi_lo_12,io_out_s_lo_lo_hi_4,7'h63}; 
  assign io_out_s_15_bits={io_out_s_hi_hi_hi_24,io_out_s_hi_hi_lo_23,5'h0,2'h1,io_out_s_lo_5,3'h1,io_out_s_lo_hi_lo_12,io_out_s_lo_lo_hi_4,7'h63}; 
  assign io_out_s_lo_lo_10=_io_out_s_opc_T_3 ? 7'h3:7'h1f; 
  assign _io_out_s_T_145={io_in[12],io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h1,io_out_s_hi_hi_lo_8,7'h13}; 
  assign _io_out_s_T_150={io_out_s_lo_1,io_in[12],io_out_s_hi_hi_2,3'h0,5'h2,3'h3,io_out_s_hi_hi_lo_8,7'h7}; 
  assign io_out_s_hi_hi_47=io_in[3:2]; 
  assign io_out_s_lo_hi_41=io_in[6:4]; 
  assign _io_out_s_T_154={io_out_s_hi_hi_47,io_in[12],io_out_s_lo_hi_41,2'h0,5'h2,3'h2,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_10}; 
  assign _io_out_s_T_158={io_out_s_lo_1,io_in[12],io_out_s_hi_hi_2,3'h0,5'h2,3'h3,io_out_s_hi_hi_lo_8,io_out_s_lo_lo_10}; 
  assign _io_out_s_mv_T={io_out_s_lo_52,5'h0,3'h0,io_out_s_hi_hi_lo_8,7'h33}; 
  assign _io_out_s_add_T={io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,io_out_s_hi_hi_lo_8,7'h33}; 
  assign io_out_s_jr={io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,12'h67}; 
  assign io_out_s_reserved_hi=io_out_s_jr[24:7]; 
  assign io_out_s_reserved={io_out_s_reserved_hi,7'h1f}; 
  assign _io_out_s_jr_reserved_T_2=_io_out_s_opc_T_3 ? io_out_s_jr:io_out_s_reserved; 
  assign _io_out_s_jr_mv_T_1=|io_out_s_lo_52; 
  assign io_out_s_mv_bits={7'b0,_io_out_s_mv_T}; 
  assign io_out_s_jr_reserved_bits={7'b0,_io_out_s_jr_reserved_T_2}; 
  assign io_out_s_jr_mv_bits=_io_out_s_jr_mv_T_1 ? io_out_s_mv_bits:io_out_s_jr_reserved_bits; 
  assign io_out_s_jr_mv_rd=_io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8:5'h0; 
  assign io_out_s_jr_mv_rs1=_io_out_s_jr_mv_T_1 ? 5'h0:io_out_s_hi_hi_lo_8; 
  assign io_out_s_jr_mv_rs2=_io_out_s_jr_mv_T_1 ? io_out_s_lo_52:io_out_s_lo_52; 
  assign io_out_s_jr_mv_rs3=_io_out_s_jr_mv_T_1 ? io_out_s_0_rs3:io_out_s_0_rs3; 
  assign io_out_s_jalr={io_out_s_lo_52,io_out_s_hi_hi_lo_8,3'h0,12'he7}; 
  assign _io_out_s_ebreak_T={io_out_s_reserved_hi,7'h73}; 
  assign io_out_s_ebreak=_io_out_s_ebreak_T|25'h100000; 
  assign _io_out_s_jalr_ebreak_T_2=_io_out_s_opc_T_3 ? io_out_s_jalr:io_out_s_ebreak; 
  assign io_out_s_add_bits={7'b0,_io_out_s_add_T}; 
  assign io_out_s_jalr_ebreak_bits={7'b0,_io_out_s_jalr_ebreak_T_2}; 
  assign io_out_s_jalr_add_bits=_io_out_s_jr_mv_T_1 ? io_out_s_add_bits:io_out_s_jalr_ebreak_bits; 
  assign io_out_s_jalr_add_rd=_io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8:5'h1; 
  assign io_out_s_jalr_add_rs1=_io_out_s_jr_mv_T_1 ? io_out_s_hi_hi_lo_8:io_out_s_hi_hi_lo_8; 
  assign io_out_s_20_bits=io_in[12] ? io_out_s_jalr_add_bits:io_out_s_jr_mv_bits; 
  assign io_out_s_20_rd=io_in[12] ? io_out_s_jalr_add_rd:io_out_s_jr_mv_rd; 
  assign io_out_s_20_rs1=io_in[12] ? io_out_s_jalr_add_rs1:io_out_s_jr_mv_rs1; 
  assign io_out_s_20_rs2=io_in[12] ? io_out_s_jr_mv_rs2:io_out_s_jr_mv_rs2; 
  assign io_out_s_20_rs3=io_in[12] ? io_out_s_jr_mv_rs3:io_out_s_jr_mv_rs3; 
  assign _io_out_s_T_163={io_out_s_lo_5,io_out_s_hi_lo_1,3'h0}; 
  assign io_out_s_hi_hi_hi_37=_io_out_s_T_163[8:5]; 
  assign io_out_s_lo_hi_lo_19=_io_out_s_T_163[4:0]; 
  assign _io_out_s_T_165={io_out_s_hi_hi_hi_37,io_out_s_lo_52,5'h2,3'h3,io_out_s_lo_hi_lo_19,7'h27}; 
  assign io_out_s_hi_hi_54=io_in[8:7]; 
  assign io_out_s_hi_lo_38=io_in[12:9]; 
  assign _io_out_s_T_169={io_out_s_hi_hi_54,io_out_s_hi_lo_38,2'h0}; 
  assign io_out_s_hi_hi_hi_38=_io_out_s_T_169[7:5]; 
  assign io_out_s_lo_hi_lo_20=_io_out_s_T_169[4:0]; 
  assign _io_out_s_T_171={io_out_s_hi_hi_hi_38,io_out_s_lo_52,5'h2,3'h2,io_out_s_lo_hi_lo_20,7'h23}; 
  assign _io_out_s_T_177={io_out_s_hi_hi_hi_37,io_out_s_lo_52,5'h2,3'h3,io_out_s_lo_hi_lo_19,7'h23}; 
  assign io_out_s_24_rs1=io_in[19:15]; 
  assign io_out_s_24_rs2=io_in[24:20]; 
  assign io_out_lo=io_in[15:13]; 
  assign _io_out_T={io_in[1:0],io_out_lo}; 
  assign _io_out_T_1=_io_out_T==5'h1; 
  assign io_out_s_1_bits={4'b0,_io_out_s_T_4}; 
  assign io_out_s_0_bits={2'b0,_io_out_s_T}; 
  assign _io_out_T_2_bits=_io_out_T_1 ? io_out_s_1_bits:io_out_s_0_bits; 
  assign _io_out_T_2_rd=_io_out_T_1 ? io_out_s_lo_hi_1:io_out_s_lo_hi_1; 
  assign _io_out_T_2_rs1=_io_out_T_1 ? io_out_s_hi_hi_lo_1:5'h2; 
  assign _io_out_T_2_rs3=_io_out_T_1 ? io_out_s_0_rs3:io_out_s_0_rs3; 
  assign _io_out_T_3=_io_out_T==5'h2; 
  assign io_out_s_2_bits={5'b0,_io_out_s_T_9}; 
  assign _io_out_T_4_bits=_io_out_T_3 ? io_out_s_2_bits:_io_out_T_2_bits; 
  assign _io_out_T_4_rd=_io_out_T_3 ? io_out_s_lo_hi_1:_io_out_T_2_rd; 
  assign _io_out_T_4_rs1=_io_out_T_3 ? io_out_s_hi_hi_lo_1:_io_out_T_2_rs1; 
  assign _io_out_T_4_rs3=_io_out_T_3 ? io_out_s_0_rs3:_io_out_T_2_rs3; 
  assign _io_out_T_5=_io_out_T==5'h3; 
  assign io_out_s_3_bits={4'b0,_io_out_s_T_14}; 
  assign _io_out_T_6_bits=_io_out_T_5 ? io_out_s_3_bits:_io_out_T_4_bits; 
  assign _io_out_T_6_rd=_io_out_T_5 ? io_out_s_lo_hi_1:_io_out_T_4_rd; 
  assign _io_out_T_6_rs1=_io_out_T_5 ? io_out_s_hi_hi_lo_1:_io_out_T_4_rs1; 
  assign _io_out_T_6_rs3=_io_out_T_5 ? io_out_s_0_rs3:_io_out_T_4_rs3; 
  assign _io_out_T_7=_io_out_T==5'h4; 
  assign io_out_s_4_bits={5'b0,_io_out_s_T_21}; 
  assign _io_out_T_8_bits=_io_out_T_7 ? io_out_s_4_bits:_io_out_T_6_bits; 
  assign _io_out_T_8_rd=_io_out_T_7 ? io_out_s_lo_hi_1:_io_out_T_6_rd; 
  assign _io_out_T_8_rs1=_io_out_T_7 ? io_out_s_hi_hi_lo_1:_io_out_T_6_rs1; 
  assign _io_out_T_8_rs3=_io_out_T_7 ? io_out_s_0_rs3:_io_out_T_6_rs3; 
  assign _io_out_T_9=_io_out_T==5'h5; 
  assign io_out_s_5_bits={4'b0,_io_out_s_T_28}; 
  assign _io_out_T_10_bits=_io_out_T_9 ? io_out_s_5_bits:_io_out_T_8_bits; 
  assign _io_out_T_10_rd=_io_out_T_9 ? io_out_s_lo_hi_1:_io_out_T_8_rd; 
  assign _io_out_T_10_rs1=_io_out_T_9 ? io_out_s_hi_hi_lo_1:_io_out_T_8_rs1; 
  assign _io_out_T_10_rs3=_io_out_T_9 ? io_out_s_0_rs3:_io_out_T_8_rs3; 
  assign _io_out_T_11=_io_out_T==5'h6; 
  assign io_out_s_6_bits={5'b0,_io_out_s_T_35}; 
  assign _io_out_T_12_bits=_io_out_T_11 ? io_out_s_6_bits:_io_out_T_10_bits; 
  assign _io_out_T_12_rd=_io_out_T_11 ? io_out_s_lo_hi_1:_io_out_T_10_rd; 
  assign _io_out_T_12_rs1=_io_out_T_11 ? io_out_s_hi_hi_lo_1:_io_out_T_10_rs1; 
  assign _io_out_T_12_rs3=_io_out_T_11 ? io_out_s_0_rs3:_io_out_T_10_rs3; 
  assign _io_out_T_13=_io_out_T==5'h7; 
  assign io_out_s_7_bits={4'b0,_io_out_s_T_42}; 
  assign _io_out_T_14_bits=_io_out_T_13 ? io_out_s_7_bits:_io_out_T_12_bits; 
  assign _io_out_T_14_rd=_io_out_T_13 ? io_out_s_lo_hi_1:_io_out_T_12_rd; 
  assign _io_out_T_14_rs1=_io_out_T_13 ? io_out_s_hi_hi_lo_1:_io_out_T_12_rs1; 
  assign _io_out_T_14_rs3=_io_out_T_13 ? io_out_s_0_rs3:_io_out_T_12_rs3; 
  assign _io_out_T_15=_io_out_T==5'h8; 
  assign _io_out_T_16_bits=_io_out_T_15 ? io_out_s_8_bits:_io_out_T_14_bits; 
  assign _io_out_T_16_rd=_io_out_T_15 ? io_out_s_hi_hi_lo_8:_io_out_T_14_rd; 
  assign _io_out_T_16_rs1=_io_out_T_15 ? io_out_s_hi_hi_lo_8:_io_out_T_14_rs1; 
  assign _io_out_T_16_rs2=_io_out_T_15 ? io_out_s_lo_hi_1:_io_out_T_14_rd; 
  assign _io_out_T_16_rs3=_io_out_T_15 ? io_out_s_0_rs3:_io_out_T_14_rs3; 
  assign _io_out_T_17=_io_out_T==5'h9; 
  assign _io_out_T_18_bits=_io_out_T_17 ? io_out_s_9_bits:_io_out_T_16_bits; 
  assign _io_out_T_18_rd=_io_out_T_17 ? io_out_s_hi_hi_lo_8:_io_out_T_16_rd; 
  assign _io_out_T_18_rs1=_io_out_T_17 ? io_out_s_hi_hi_lo_8:_io_out_T_16_rs1; 
  assign _io_out_T_18_rs2=_io_out_T_17 ? io_out_s_lo_hi_1:_io_out_T_16_rs2; 
  assign _io_out_T_18_rs3=_io_out_T_17 ? io_out_s_0_rs3:_io_out_T_16_rs3; 
  assign _io_out_T_19=_io_out_T==5'ha; 
  assign _io_out_T_20_bits=_io_out_T_19 ? io_out_s_10_bits:_io_out_T_18_bits; 
  assign _io_out_T_20_rd=_io_out_T_19 ? io_out_s_hi_hi_lo_8:_io_out_T_18_rd; 
  assign _io_out_T_20_rs1=_io_out_T_19 ? 5'h0:_io_out_T_18_rs1; 
  assign _io_out_T_20_rs2=_io_out_T_19 ? io_out_s_lo_hi_1:_io_out_T_18_rs2; 
  assign _io_out_T_20_rs3=_io_out_T_19 ? io_out_s_0_rs3:_io_out_T_18_rs3; 
  assign _io_out_T_21=_io_out_T==5'hb; 
  assign _io_out_T_22_bits=_io_out_T_21 ? io_out_s_11_bits:_io_out_T_20_bits; 
  assign _io_out_T_22_rd=_io_out_T_21 ? io_out_s_11_rd:_io_out_T_20_rd; 
  assign _io_out_T_22_rs1=_io_out_T_21 ? io_out_s_11_rd:_io_out_T_20_rs1; 
  assign _io_out_T_22_rs2=_io_out_T_21 ? io_out_s_11_rs2:_io_out_T_20_rs2; 
  assign _io_out_T_22_rs3=_io_out_T_21 ? io_out_s_11_rs3:_io_out_T_20_rs3; 
  assign _io_out_T_23=_io_out_T==5'hc; 
  assign _io_out_T_24_bits=_io_out_T_23 ? io_out_s_12_bits:_io_out_T_22_bits; 
  assign _io_out_T_24_rd=_io_out_T_23 ? io_out_s_hi_hi_lo_1:_io_out_T_22_rd; 
  assign _io_out_T_24_rs1=_io_out_T_23 ? io_out_s_hi_hi_lo_1:_io_out_T_22_rs1; 
  assign _io_out_T_24_rs2=_io_out_T_23 ? io_out_s_lo_hi_1:_io_out_T_22_rs2; 
  assign _io_out_T_24_rs3=_io_out_T_23 ? io_out_s_0_rs3:_io_out_T_22_rs3; 
  assign _io_out_T_25=_io_out_T==5'hd; 
  assign _io_out_T_26_bits=_io_out_T_25 ? io_out_s_13_bits:_io_out_T_24_bits; 
  assign _io_out_T_26_rd=_io_out_T_25 ? 5'h0:_io_out_T_24_rd; 
  assign _io_out_T_26_rs1=_io_out_T_25 ? io_out_s_hi_hi_lo_1:_io_out_T_24_rs1; 
  assign _io_out_T_26_rs2=_io_out_T_25 ? io_out_s_lo_hi_1:_io_out_T_24_rs2; 
  assign _io_out_T_26_rs3=_io_out_T_25 ? io_out_s_0_rs3:_io_out_T_24_rs3; 
  assign _io_out_T_27=_io_out_T==5'he; 
  assign _io_out_T_28_bits=_io_out_T_27 ? io_out_s_14_bits:_io_out_T_26_bits; 
  assign _io_out_T_28_rd=_io_out_T_27 ? io_out_s_hi_hi_lo_1:_io_out_T_26_rd; 
  assign _io_out_T_28_rs1=_io_out_T_27 ? io_out_s_hi_hi_lo_1:_io_out_T_26_rs1; 
  assign _io_out_T_28_rs2=_io_out_T_27 ? 5'h0:_io_out_T_26_rs2; 
  assign _io_out_T_28_rs3=_io_out_T_27 ? io_out_s_0_rs3:_io_out_T_26_rs3; 
  assign _io_out_T_29=_io_out_T==5'hf; 
  assign _io_out_T_30_bits=_io_out_T_29 ? io_out_s_15_bits:_io_out_T_28_bits; 
  assign _io_out_T_30_rd=_io_out_T_29 ? 5'h0:_io_out_T_28_rd; 
  assign _io_out_T_30_rs1=_io_out_T_29 ? io_out_s_hi_hi_lo_1:_io_out_T_28_rs1; 
  assign _io_out_T_30_rs2=_io_out_T_29 ? 5'h0:_io_out_T_28_rs2; 
  assign _io_out_T_30_rs3=_io_out_T_29 ? io_out_s_0_rs3:_io_out_T_28_rs3; 
  assign _io_out_T_31=_io_out_T==5'h10; 
  assign io_out_s_16_bits={6'b0,_io_out_s_T_145}; 
  assign _io_out_T_32_bits=_io_out_T_31 ? io_out_s_16_bits:_io_out_T_30_bits; 
  assign _io_out_T_32_rd=_io_out_T_31 ? io_out_s_hi_hi_lo_8:_io_out_T_30_rd; 
  assign _io_out_T_32_rs1=_io_out_T_31 ? io_out_s_hi_hi_lo_8:_io_out_T_30_rs1; 
  assign _io_out_T_32_rs2=_io_out_T_31 ? io_out_s_lo_52:_io_out_T_30_rs2; 
  assign _io_out_T_32_rs3=_io_out_T_31 ? io_out_s_0_rs3:_io_out_T_30_rs3; 
  assign _io_out_T_33=_io_out_T==5'h11; 
  assign io_out_s_17_bits={3'b0,_io_out_s_T_150}; 
  assign _io_out_T_34_bits=_io_out_T_33 ? io_out_s_17_bits:_io_out_T_32_bits; 
  assign _io_out_T_34_rd=_io_out_T_33 ? io_out_s_hi_hi_lo_8:_io_out_T_32_rd; 
  assign _io_out_T_34_rs1=_io_out_T_33 ? 5'h2:_io_out_T_32_rs1; 
  assign _io_out_T_34_rs2=_io_out_T_33 ? io_out_s_lo_52:_io_out_T_32_rs2; 
  assign _io_out_T_34_rs3=_io_out_T_33 ? io_out_s_0_rs3:_io_out_T_32_rs3; 
  assign _io_out_T_35=_io_out_T==5'h12; 
  assign io_out_s_18_bits={4'b0,_io_out_s_T_154}; 
  assign _io_out_T_36_bits=_io_out_T_35 ? io_out_s_18_bits:_io_out_T_34_bits; 
  assign _io_out_T_36_rd=_io_out_T_35 ? io_out_s_hi_hi_lo_8:_io_out_T_34_rd; 
  assign _io_out_T_36_rs1=_io_out_T_35 ? 5'h2:_io_out_T_34_rs1; 
  assign _io_out_T_36_rs2=_io_out_T_35 ? io_out_s_lo_52:_io_out_T_34_rs2; 
  assign _io_out_T_36_rs3=_io_out_T_35 ? io_out_s_0_rs3:_io_out_T_34_rs3; 
  assign _io_out_T_37=_io_out_T==5'h13; 
  assign io_out_s_19_bits={3'b0,_io_out_s_T_158}; 
  assign _io_out_T_38_bits=_io_out_T_37 ? io_out_s_19_bits:_io_out_T_36_bits; 
  assign _io_out_T_38_rd=_io_out_T_37 ? io_out_s_hi_hi_lo_8:_io_out_T_36_rd; 
  assign _io_out_T_38_rs1=_io_out_T_37 ? 5'h2:_io_out_T_36_rs1; 
  assign _io_out_T_38_rs2=_io_out_T_37 ? io_out_s_lo_52:_io_out_T_36_rs2; 
  assign _io_out_T_38_rs3=_io_out_T_37 ? io_out_s_0_rs3:_io_out_T_36_rs3; 
  assign _io_out_T_39=_io_out_T==5'h14; 
  assign _io_out_T_40_bits=_io_out_T_39 ? io_out_s_20_bits:_io_out_T_38_bits; 
  assign _io_out_T_40_rd=_io_out_T_39 ? io_out_s_20_rd:_io_out_T_38_rd; 
  assign _io_out_T_40_rs1=_io_out_T_39 ? io_out_s_20_rs1:_io_out_T_38_rs1; 
  assign _io_out_T_40_rs2=_io_out_T_39 ? io_out_s_20_rs2:_io_out_T_38_rs2; 
  assign _io_out_T_40_rs3=_io_out_T_39 ? io_out_s_20_rs3:_io_out_T_38_rs3; 
  assign _io_out_T_41=_io_out_T==5'h15; 
  assign io_out_s_21_bits={3'b0,_io_out_s_T_165}; 
  assign _io_out_T_42_bits=_io_out_T_41 ? io_out_s_21_bits:_io_out_T_40_bits; 
  assign _io_out_T_42_rd=_io_out_T_41 ? io_out_s_hi_hi_lo_8:_io_out_T_40_rd; 
  assign _io_out_T_42_rs1=_io_out_T_41 ? 5'h2:_io_out_T_40_rs1; 
  assign _io_out_T_42_rs2=_io_out_T_41 ? io_out_s_lo_52:_io_out_T_40_rs2; 
  assign _io_out_T_42_rs3=_io_out_T_41 ? io_out_s_0_rs3:_io_out_T_40_rs3; 
  assign _io_out_T_43=_io_out_T==5'h16; 
  assign io_out_s_22_bits={4'b0,_io_out_s_T_171}; 
  assign _io_out_T_44_bits=_io_out_T_43 ? io_out_s_22_bits:_io_out_T_42_bits; 
  assign _io_out_T_44_rd=_io_out_T_43 ? io_out_s_hi_hi_lo_8:_io_out_T_42_rd; 
  assign _io_out_T_44_rs1=_io_out_T_43 ? 5'h2:_io_out_T_42_rs1; 
  assign _io_out_T_44_rs2=_io_out_T_43 ? io_out_s_lo_52:_io_out_T_42_rs2; 
  assign _io_out_T_44_rs3=_io_out_T_43 ? io_out_s_0_rs3:_io_out_T_42_rs3; 
  assign _io_out_T_45=_io_out_T==5'h17; 
  assign io_out_s_23_bits={3'b0,_io_out_s_T_177}; 
  assign _io_out_T_46_bits=_io_out_T_45 ? io_out_s_23_bits:_io_out_T_44_bits; 
  assign _io_out_T_46_rd=_io_out_T_45 ? io_out_s_hi_hi_lo_8:_io_out_T_44_rd; 
  assign _io_out_T_46_rs1=_io_out_T_45 ? 5'h2:_io_out_T_44_rs1; 
  assign _io_out_T_46_rs2=_io_out_T_45 ? io_out_s_lo_52:_io_out_T_44_rs2; 
  assign _io_out_T_46_rs3=_io_out_T_45 ? io_out_s_0_rs3:_io_out_T_44_rs3; 
  assign _io_out_T_47=_io_out_T==5'h18; 
  assign _io_out_T_48_bits=_io_out_T_47 ? io_in:_io_out_T_46_bits; 
  assign _io_out_T_48_rd=_io_out_T_47 ? io_out_s_hi_hi_lo_8:_io_out_T_46_rd; 
  assign _io_out_T_48_rs1=_io_out_T_47 ? io_out_s_24_rs1:_io_out_T_46_rs1; 
  assign _io_out_T_48_rs2=_io_out_T_47 ? io_out_s_24_rs2:_io_out_T_46_rs2; 
  assign _io_out_T_48_rs3=_io_out_T_47 ? io_out_s_0_rs3:_io_out_T_46_rs3; 
  assign _io_out_T_49=_io_out_T==5'h19; 
  assign _io_out_T_50_bits=_io_out_T_49 ? io_in:_io_out_T_48_bits; 
  assign _io_out_T_50_rd=_io_out_T_49 ? io_out_s_hi_hi_lo_8:_io_out_T_48_rd; 
  assign _io_out_T_50_rs1=_io_out_T_49 ? io_out_s_24_rs1:_io_out_T_48_rs1; 
  assign _io_out_T_50_rs2=_io_out_T_49 ? io_out_s_24_rs2:_io_out_T_48_rs2; 
  assign _io_out_T_50_rs3=_io_out_T_49 ? io_out_s_0_rs3:_io_out_T_48_rs3; 
  assign _io_out_T_51=_io_out_T==5'h1a; 
  assign _io_out_T_52_bits=_io_out_T_51 ? io_in:_io_out_T_50_bits; 
  assign _io_out_T_52_rd=_io_out_T_51 ? io_out_s_hi_hi_lo_8:_io_out_T_50_rd; 
  assign _io_out_T_52_rs1=_io_out_T_51 ? io_out_s_24_rs1:_io_out_T_50_rs1; 
  assign _io_out_T_52_rs2=_io_out_T_51 ? io_out_s_24_rs2:_io_out_T_50_rs2; 
  assign _io_out_T_52_rs3=_io_out_T_51 ? io_out_s_0_rs3:_io_out_T_50_rs3; 
  assign _io_out_T_53=_io_out_T==5'h1b; 
  assign _io_out_T_54_bits=_io_out_T_53 ? io_in:_io_out_T_52_bits; 
  assign _io_out_T_54_rd=_io_out_T_53 ? io_out_s_hi_hi_lo_8:_io_out_T_52_rd; 
  assign _io_out_T_54_rs1=_io_out_T_53 ? io_out_s_24_rs1:_io_out_T_52_rs1; 
  assign _io_out_T_54_rs2=_io_out_T_53 ? io_out_s_24_rs2:_io_out_T_52_rs2; 
  assign _io_out_T_54_rs3=_io_out_T_53 ? io_out_s_0_rs3:_io_out_T_52_rs3; 
  assign _io_out_T_55=_io_out_T==5'h1c; 
  assign _io_out_T_56_bits=_io_out_T_55 ? io_in:_io_out_T_54_bits; 
  assign _io_out_T_56_rd=_io_out_T_55 ? io_out_s_hi_hi_lo_8:_io_out_T_54_rd; 
  assign _io_out_T_56_rs1=_io_out_T_55 ? io_out_s_24_rs1:_io_out_T_54_rs1; 
  assign _io_out_T_56_rs2=_io_out_T_55 ? io_out_s_24_rs2:_io_out_T_54_rs2; 
  assign _io_out_T_56_rs3=_io_out_T_55 ? io_out_s_0_rs3:_io_out_T_54_rs3; 
  assign _io_out_T_57=_io_out_T==5'h1d; 
  assign _io_out_T_58_bits=_io_out_T_57 ? io_in:_io_out_T_56_bits; 
  assign _io_out_T_58_rd=_io_out_T_57 ? io_out_s_hi_hi_lo_8:_io_out_T_56_rd; 
  assign _io_out_T_58_rs1=_io_out_T_57 ? io_out_s_24_rs1:_io_out_T_56_rs1; 
  assign _io_out_T_58_rs2=_io_out_T_57 ? io_out_s_24_rs2:_io_out_T_56_rs2; 
  assign _io_out_T_58_rs3=_io_out_T_57 ? io_out_s_0_rs3:_io_out_T_56_rs3; 
  assign _io_out_T_59=_io_out_T==5'h1e; 
  assign _io_out_T_60_bits=_io_out_T_59 ? io_in:_io_out_T_58_bits; 
  assign _io_out_T_60_rd=_io_out_T_59 ? io_out_s_hi_hi_lo_8:_io_out_T_58_rd; 
  assign _io_out_T_60_rs1=_io_out_T_59 ? io_out_s_24_rs1:_io_out_T_58_rs1; 
  assign _io_out_T_60_rs2=_io_out_T_59 ? io_out_s_24_rs2:_io_out_T_58_rs2; 
  assign _io_out_T_60_rs3=_io_out_T_59 ? io_out_s_0_rs3:_io_out_T_58_rs3; 
  assign _io_out_T_61=_io_out_T==5'h1f; 
  assign io_out_bits=_io_out_T_61 ? io_in:_io_out_T_60_bits; 
  assign io_out_rd=_io_out_T_61 ? io_out_s_hi_hi_lo_8:_io_out_T_60_rd; 
  assign io_out_rs1=_io_out_T_61 ? io_out_s_24_rs1:_io_out_T_60_rs1; 
  assign io_out_rs2=_io_out_T_61 ? io_out_s_24_rs2:_io_out_T_60_rs2; 
  assign io_out_rs3=_io_out_T_61 ? io_out_s_0_rs3:_io_out_T_60_rs3; 
  assign io_rvc=io_in[1:0]!=2'h3; 
  assign RVCExpander_covSum=30'h0; 
  assign io_covSum=RVCExpander_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module MulAddRecFNToRaw_preMul (
  input [1:0] io_op,
  input [32:0] io_a,
  input [32:0] io_b,
  input [32:0] io_c,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output io_toPostMul_isSigNaNAny,
  output io_toPostMul_isNaNAOrB,
  output io_toPostMul_isInfA,
  output io_toPostMul_isZeroA,
  output io_toPostMul_isInfB,
  output io_toPostMul_isZeroB,
  output io_toPostMul_signProd,
  output io_toPostMul_isNaNC,
  output io_toPostMul_isInfC,
  output io_toPostMul_isZeroC,
  output [9:0] io_toPostMul_sExpSum,
  output io_toPostMul_doSubMags,
  output io_toPostMul_CIsDominant,
  output [4:0] io_toPostMul_CDom_CAlignDist,
  output [25:0] io_toPostMul_highAlignedSigC,
  output io_toPostMul_bit0AlignedSigC,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [8:0] rawA_exp ;  
   wire rawA_isZero ;  
   wire rawA_isSpecial ;  
   wire rawA__isNaN ;  
   wire rawA__sign ;  
   wire [9:0] rawA__sExp ;  
   wire rawA_out_sig_hi_lo ;  
   wire [22:0] rawA_out_sig_lo ;  
   wire [24:0] rawA__sig ;  
   wire [8:0] rawB_exp ;  
   wire rawB_isZero ;  
   wire rawB_isSpecial ;  
   wire rawB__isNaN ;  
   wire rawB__sign ;  
   wire [9:0] rawB__sExp ;  
   wire rawB_out_sig_hi_lo ;  
   wire [22:0] rawB_out_sig_lo ;  
   wire [24:0] rawB__sig ;  
   wire [8:0] rawC_exp ;  
   wire rawC_isZero ;  
   wire rawC_isSpecial ;  
   wire rawC__isNaN ;  
   wire rawC__sign ;  
   wire [9:0] rawC__sExp ;  
   wire rawC_out_sig_hi_lo ;  
   wire [22:0] rawC_out_sig_lo ;  
   wire [24:0] rawC__sig ;  
   wire _signProd_T ;  
   wire signProd ;  
   wire [10:0] _sExpAlignedProd_T ;  
   wire [10:0] sExpAlignedProd ;  
   wire _doSubMags_T ;  
   wire doSubMags ;  
   wire [10:0] _GEN_0 ;  
   wire [10:0] sNatCAlignDist ;  
   wire [9:0] posNatCAlignDist ;  
   wire _isMinCAlign_T ;  
   wire _isMinCAlign_T_1 ;  
   wire isMinCAlign ;  
   wire _CIsDominant_T_1 ;  
   wire _CIsDominant_T_2 ;  
   wire CIsDominant ;  
   wire _CAlignDist_T ;  
   wire [6:0] _CAlignDist_T_2 ;  
   wire [6:0] CAlignDist ;  
   wire [24:0] mainAlignedSigC_hi ;  
   wire [52:0] mainAlignedSigC_lo ;  
   wire [77:0] _mainAlignedSigC_T_3 ;  
   wire [77:0] mainAlignedSigC ;  
   wire [26:0] _reduced4CExtra_T ;  
   wire reduced4CExtra_reducedVec_0 ;  
   wire reduced4CExtra_reducedVec_1 ;  
   wire reduced4CExtra_reducedVec_2 ;  
   wire reduced4CExtra_reducedVec_3 ;  
   wire reduced4CExtra_reducedVec_4 ;  
   wire reduced4CExtra_reducedVec_5 ;  
   wire reduced4CExtra_reducedVec_6 ;  
   wire [6:0] _reduced4CExtra_T_1 ;  
   wire [32:0] reduced4CExtra_shift ;  
   wire reduced4CExtra_hi_1 ;  
   wire reduced4CExtra_lo_1 ;  
   wire reduced4CExtra_hi_3 ;  
   wire reduced4CExtra_lo_2 ;  
   wire reduced4CExtra_hi_5 ;  
   wire reduced4CExtra_lo_4 ;  
   wire [5:0] _reduced4CExtra_T_8 ;  
   wire [6:0] _GEN_1 ;  
   wire [6:0] _reduced4CExtra_T_9 ;  
   wire reduced4CExtra ;  
   wire _alignedSigC_T_2 ;  
   wire _alignedSigC_T_4 ;  
   wire _alignedSigC_T_6 ;  
   wire _alignedSigC_T_7 ;  
   wire alignedSigC_lo ;  
   wire [74:0] alignedSigC_hi ;  
   wire [75:0] alignedSigC ;  
   wire _io_toPostMul_isSigNaNAny_T_2 ;  
   wire _io_toPostMul_isSigNaNAny_T_5 ;  
   wire _io_toPostMul_isSigNaNAny_T_6 ;  
   wire _io_toPostMul_isSigNaNAny_T_9 ;  
   wire [10:0] _io_toPostMul_sExpSum_T_2 ;  
   wire [10:0] _io_toPostMul_sExpSum_T_3 ;  
   wire [29:0] MulAddRecFNToRaw_preMul_covSum ;  
  assign rawA_exp=io_a[31:23]; 
  assign rawA_isZero=rawA_exp[8:6]==3'h0; 
  assign rawA_isSpecial=rawA_exp[8:7]==2'h3; 
  assign rawA__isNaN=rawA_isSpecial&rawA_exp[6]; 
  assign rawA__sign=io_a[32]; 
  assign rawA__sExp={1'b0,$signed(rawA_exp)}; 
  assign rawA_out_sig_hi_lo=~rawA_isZero; 
  assign rawA_out_sig_lo=io_a[22:0]; 
  assign rawA__sig={1'h0,rawA_out_sig_hi_lo,rawA_out_sig_lo}; 
  assign rawB_exp=io_b[31:23]; 
  assign rawB_isZero=rawB_exp[8:6]==3'h0; 
  assign rawB_isSpecial=rawB_exp[8:7]==2'h3; 
  assign rawB__isNaN=rawB_isSpecial&rawB_exp[6]; 
  assign rawB__sign=io_b[32]; 
  assign rawB__sExp={1'b0,$signed(rawB_exp)}; 
  assign rawB_out_sig_hi_lo=~rawB_isZero; 
  assign rawB_out_sig_lo=io_b[22:0]; 
  assign rawB__sig={1'h0,rawB_out_sig_hi_lo,rawB_out_sig_lo}; 
  assign rawC_exp=io_c[31:23]; 
  assign rawC_isZero=rawC_exp[8:6]==3'h0; 
  assign rawC_isSpecial=rawC_exp[8:7]==2'h3; 
  assign rawC__isNaN=rawC_isSpecial&rawC_exp[6]; 
  assign rawC__sign=io_c[32]; 
  assign rawC__sExp={1'b0,$signed(rawC_exp)}; 
  assign rawC_out_sig_hi_lo=~rawC_isZero; 
  assign rawC_out_sig_lo=io_c[22:0]; 
  assign rawC__sig={1'h0,rawC_out_sig_hi_lo,rawC_out_sig_lo}; 
  assign _signProd_T=rawA__sign^rawB__sign; 
  assign signProd=_signProd_T^io_op[1]; 
  assign _sExpAlignedProd_T=$signed(rawA__sExp)+$signed(rawB__sExp); 
  assign sExpAlignedProd=$signed(_sExpAlignedProd_T)+-11'she5; 
  assign _doSubMags_T=signProd^rawC__sign; 
  assign doSubMags=_doSubMags_T^io_op[0]; 
  assign _GEN_0={{1{rawC__sExp[9]}},rawC__sExp}; 
  assign sNatCAlignDist=$signed(sExpAlignedProd)-$signed(_GEN_0); 
  assign posNatCAlignDist=sNatCAlignDist[9:0]; 
  assign _isMinCAlign_T=rawA_isZero|rawB_isZero; 
  assign _isMinCAlign_T_1=$signed(sNatCAlignDist)<11'sh0; 
  assign isMinCAlign=_isMinCAlign_T|_isMinCAlign_T_1; 
  assign _CIsDominant_T_1=posNatCAlignDist<=10'h18; 
  assign _CIsDominant_T_2=isMinCAlign|_CIsDominant_T_1; 
  assign CIsDominant=rawC_out_sig_hi_lo&_CIsDominant_T_2; 
  assign _CAlignDist_T=posNatCAlignDist<10'h4a; 
  assign _CAlignDist_T_2=_CAlignDist_T ? posNatCAlignDist[6:0]:7'h4a; 
  assign CAlignDist=isMinCAlign ? 7'h0:_CAlignDist_T_2; 
  assign mainAlignedSigC_hi=doSubMags ? ~rawC__sig:rawC__sig; 
  assign mainAlignedSigC_lo=doSubMags ? 53'h1fffffffffffff:53'h0; 
  assign _mainAlignedSigC_T_3={mainAlignedSigC_hi,mainAlignedSigC_lo}; 
  assign mainAlignedSigC=$signed(_mainAlignedSigC_T_3)>>>CAlignDist; 
  assign _reduced4CExtra_T={rawC__sig,2'h0}; 
  assign reduced4CExtra_reducedVec_0=|_reduced4CExtra_T[3:0]; 
  assign reduced4CExtra_reducedVec_1=|_reduced4CExtra_T[7:4]; 
  assign reduced4CExtra_reducedVec_2=|_reduced4CExtra_T[11:8]; 
  assign reduced4CExtra_reducedVec_3=|_reduced4CExtra_T[15:12]; 
  assign reduced4CExtra_reducedVec_4=|_reduced4CExtra_T[19:16]; 
  assign reduced4CExtra_reducedVec_5=|_reduced4CExtra_T[23:20]; 
  assign reduced4CExtra_reducedVec_6=|_reduced4CExtra_T[26:24]; 
  assign _reduced4CExtra_T_1={reduced4CExtra_reducedVec_6,reduced4CExtra_reducedVec_5,reduced4CExtra_reducedVec_4,reduced4CExtra_reducedVec_3,reduced4CExtra_reducedVec_2,reduced4CExtra_reducedVec_1,reduced4CExtra_reducedVec_0}; 
  assign reduced4CExtra_shift=-33'sh100000000>>>CAlignDist[6:2]; 
  assign reduced4CExtra_hi_1=reduced4CExtra_shift[14]; 
  assign reduced4CExtra_lo_1=reduced4CExtra_shift[15]; 
  assign reduced4CExtra_hi_3=reduced4CExtra_shift[16]; 
  assign reduced4CExtra_lo_2=reduced4CExtra_shift[17]; 
  assign reduced4CExtra_hi_5=reduced4CExtra_shift[18]; 
  assign reduced4CExtra_lo_4=reduced4CExtra_shift[19]; 
  assign _reduced4CExtra_T_8={reduced4CExtra_hi_1,reduced4CExtra_lo_1,reduced4CExtra_hi_3,reduced4CExtra_lo_2,reduced4CExtra_hi_5,reduced4CExtra_lo_4}; 
  assign _GEN_1={1'b0,_reduced4CExtra_T_8}; 
  assign _reduced4CExtra_T_9=_reduced4CExtra_T_1&_GEN_1; 
  assign reduced4CExtra=|_reduced4CExtra_T_9; 
  assign _alignedSigC_T_2=&mainAlignedSigC[2:0]; 
  assign _alignedSigC_T_4=_alignedSigC_T_2&~reduced4CExtra; 
  assign _alignedSigC_T_6=|mainAlignedSigC[2:0]; 
  assign _alignedSigC_T_7=_alignedSigC_T_6|reduced4CExtra; 
  assign alignedSigC_lo=doSubMags ? _alignedSigC_T_4:_alignedSigC_T_7; 
  assign alignedSigC_hi=mainAlignedSigC[77:3]; 
  assign alignedSigC={alignedSigC_hi,alignedSigC_lo}; 
  assign _io_toPostMul_isSigNaNAny_T_2=rawA__isNaN&~rawA__sig[22]; 
  assign _io_toPostMul_isSigNaNAny_T_5=rawB__isNaN&~rawB__sig[22]; 
  assign _io_toPostMul_isSigNaNAny_T_6=_io_toPostMul_isSigNaNAny_T_2|_io_toPostMul_isSigNaNAny_T_5; 
  assign _io_toPostMul_isSigNaNAny_T_9=rawC__isNaN&~rawC__sig[22]; 
  assign _io_toPostMul_sExpSum_T_2=$signed(sExpAlignedProd)-11'sh18; 
  assign _io_toPostMul_sExpSum_T_3=CIsDominant ? $signed({{1{rawC__sExp[9]}},rawC__sExp}):$signed(_io_toPostMul_sExpSum_T_2); 
  assign io_mulAddA=rawA__sig[23:0]; 
  assign io_mulAddB=rawB__sig[23:0]; 
  assign io_mulAddC=alignedSigC[48:1]; 
  assign io_toPostMul_isSigNaNAny=_io_toPostMul_isSigNaNAny_T_6|_io_toPostMul_isSigNaNAny_T_9; 
  assign io_toPostMul_isNaNAOrB=rawA__isNaN|rawB__isNaN; 
  assign io_toPostMul_isInfA=rawA_isSpecial&~rawA_exp[6]; 
  assign io_toPostMul_isZeroA=rawA_exp[8:6]==3'h0; 
  assign io_toPostMul_isInfB=rawB_isSpecial&~rawB_exp[6]; 
  assign io_toPostMul_isZeroB=rawB_exp[8:6]==3'h0; 
  assign io_toPostMul_signProd=_signProd_T^io_op[1]; 
  assign io_toPostMul_isNaNC=rawC_isSpecial&rawC_exp[6]; 
  assign io_toPostMul_isInfC=rawC_isSpecial&~rawC_exp[6]; 
  assign io_toPostMul_isZeroC=rawC_exp[8:6]==3'h0; 
  assign io_toPostMul_sExpSum=_io_toPostMul_sExpSum_T_3[9:0]; 
  assign io_toPostMul_doSubMags=_doSubMags_T^io_op[0]; 
  assign io_toPostMul_CIsDominant=rawC_out_sig_hi_lo&_CIsDominant_T_2; 
  assign io_toPostMul_CDom_CAlignDist=CAlignDist[4:0]; 
  assign io_toPostMul_highAlignedSigC=alignedSigC[74:49]; 
  assign io_toPostMul_bit0AlignedSigC=alignedSigC[0]; 
  assign MulAddRecFNToRaw_preMul_covSum=30'h0; 
  assign io_covSum=MulAddRecFNToRaw_preMul_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module MulAddRecFNToRaw_postMul (
  input io_fromPreMul_isSigNaNAny,
  input io_fromPreMul_isNaNAOrB,
  input io_fromPreMul_isInfA,
  input io_fromPreMul_isZeroA,
  input io_fromPreMul_isInfB,
  input io_fromPreMul_isZeroB,
  input io_fromPreMul_signProd,
  input io_fromPreMul_isNaNC,
  input io_fromPreMul_isInfC,
  input io_fromPreMul_isZeroC,
  input [9:0] io_fromPreMul_sExpSum,
  input io_fromPreMul_doSubMags,
  input io_fromPreMul_CIsDominant,
  input [4:0] io_fromPreMul_CDom_CAlignDist,
  input [25:0] io_fromPreMul_highAlignedSigC,
  input io_fromPreMul_bit0AlignedSigC,
  input [48:0] io_mulAddResult,
  input [2:0] io_roundingMode,
  output io_invalidExc,
  output io_rawOut_isNaN,
  output io_rawOut_isInf,
  output io_rawOut_isZero,
  output io_rawOut_sign,
  output [9:0] io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundingMode_min ;  
   wire CDom_sign ;  
   wire [25:0] _sigSum_T_2 ;  
   wire [25:0] sigSum_hi_hi ;  
   wire [47:0] sigSum_hi_lo ;  
   wire [74:0] sigSum ;  
   wire [1:0] _CDom_sExp_T ;  
   wire [9:0] _GEN_0 ;  
   wire [9:0] CDom_sExp ;  
   wire [1:0] CDom_absSigSum_hi_lo ;  
   wire [46:0] CDom_absSigSum_lo ;  
   wire [49:0] _CDom_absSigSum_T_2 ;  
   wire [49:0] CDom_absSigSum ;  
   wire _CDom_absSigSumExtra_T_2 ;  
   wire _CDom_absSigSumExtra_T_4 ;  
   wire CDom_absSigSumExtra ;  
   wire [80:0] _GEN_1 ;  
   wire [80:0] _CDom_mainSig_T ;  
   wire [28:0] CDom_mainSig ;  
   wire [26:0] _CDom_reduced4SigExtra_T_1 ;  
   wire CDom_reduced4SigExtra_reducedVec_0 ;  
   wire CDom_reduced4SigExtra_reducedVec_1 ;  
   wire CDom_reduced4SigExtra_reducedVec_2 ;  
   wire CDom_reduced4SigExtra_reducedVec_3 ;  
   wire CDom_reduced4SigExtra_reducedVec_4 ;  
   wire CDom_reduced4SigExtra_reducedVec_5 ;  
   wire CDom_reduced4SigExtra_reducedVec_6 ;  
   wire [6:0] _CDom_reduced4SigExtra_T_2 ;  
   wire [8:0] CDom_reduced4SigExtra_shift ;  
   wire CDom_reduced4SigExtra_hi_1 ;  
   wire CDom_reduced4SigExtra_lo_1 ;  
   wire CDom_reduced4SigExtra_hi_3 ;  
   wire CDom_reduced4SigExtra_lo_2 ;  
   wire CDom_reduced4SigExtra_hi_5 ;  
   wire CDom_reduced4SigExtra_lo_4 ;  
   wire [5:0] _CDom_reduced4SigExtra_T_10 ;  
   wire [6:0] _GEN_2 ;  
   wire [6:0] _CDom_reduced4SigExtra_T_11 ;  
   wire CDom_reduced4SigExtra ;  
   wire [25:0] CDom_sig_hi ;  
   wire _CDom_sig_T_1 ;  
   wire _CDom_sig_T_2 ;  
   wire CDom_sig_lo ;  
   wire [26:0] CDom_sig ;  
   wire notCDom_signSigSum ;  
   wire [50:0] _GEN_3 ;  
   wire [50:0] _notCDom_absSigSum_T_4 ;  
   wire [50:0] notCDom_absSigSum ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_0 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_1 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_2 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_3 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_4 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_5 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_6 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_7 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_8 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_9 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_10 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_11 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_12 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_13 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_14 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_15 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_16 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_17 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_18 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_19 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_20 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_21 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_22 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_23 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_24 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_25 ;  
   wire [5:0] notCDom_reduced2AbsSigSum_lo_lo ;  
   wire [12:0] notCDom_reduced2AbsSigSum_lo ;  
   wire [5:0] notCDom_reduced2AbsSigSum_hi_lo ;  
   wire [25:0] notCDom_reduced2AbsSigSum ;  
   wire [4:0] _notCDom_normDistReduced2_T_26 ;  
   wire [4:0] _notCDom_normDistReduced2_T_27 ;  
   wire [4:0] _notCDom_normDistReduced2_T_28 ;  
   wire [4:0] _notCDom_normDistReduced2_T_29 ;  
   wire [4:0] _notCDom_normDistReduced2_T_30 ;  
   wire [4:0] _notCDom_normDistReduced2_T_31 ;  
   wire [4:0] _notCDom_normDistReduced2_T_32 ;  
   wire [4:0] _notCDom_normDistReduced2_T_33 ;  
   wire [4:0] _notCDom_normDistReduced2_T_34 ;  
   wire [4:0] _notCDom_normDistReduced2_T_35 ;  
   wire [4:0] _notCDom_normDistReduced2_T_36 ;  
   wire [4:0] _notCDom_normDistReduced2_T_37 ;  
   wire [4:0] _notCDom_normDistReduced2_T_38 ;  
   wire [4:0] _notCDom_normDistReduced2_T_39 ;  
   wire [4:0] _notCDom_normDistReduced2_T_40 ;  
   wire [4:0] _notCDom_normDistReduced2_T_41 ;  
   wire [4:0] _notCDom_normDistReduced2_T_42 ;  
   wire [4:0] _notCDom_normDistReduced2_T_43 ;  
   wire [4:0] _notCDom_normDistReduced2_T_44 ;  
   wire [4:0] _notCDom_normDistReduced2_T_45 ;  
   wire [4:0] _notCDom_normDistReduced2_T_46 ;  
   wire [4:0] _notCDom_normDistReduced2_T_47 ;  
   wire [4:0] _notCDom_normDistReduced2_T_48 ;  
   wire [4:0] _notCDom_normDistReduced2_T_49 ;  
   wire [4:0] notCDom_normDistReduced2 ;  
   wire [5:0] notCDom_nearNormDist ;  
   wire [6:0] _notCDom_sExp_T ;  
   wire [9:0] _GEN_4 ;  
   wire [9:0] notCDom_sExp ;  
   wire [113:0] _GEN_5 ;  
   wire [113:0] _notCDom_mainSig_T ;  
   wire [28:0] notCDom_mainSig ;  
   wire notCDom_reduced4SigExtra_reducedVec_0 ;  
   wire notCDom_reduced4SigExtra_reducedVec_1 ;  
   wire notCDom_reduced4SigExtra_reducedVec_2 ;  
   wire notCDom_reduced4SigExtra_reducedVec_3 ;  
   wire notCDom_reduced4SigExtra_reducedVec_4 ;  
   wire notCDom_reduced4SigExtra_reducedVec_5 ;  
   wire notCDom_reduced4SigExtra_reducedVec_6 ;  
   wire [6:0] _notCDom_reduced4SigExtra_T_2 ;  
   wire [16:0] notCDom_reduced4SigExtra_shift ;  
   wire notCDom_reduced4SigExtra_hi_1 ;  
   wire notCDom_reduced4SigExtra_lo_1 ;  
   wire notCDom_reduced4SigExtra_hi_3 ;  
   wire notCDom_reduced4SigExtra_lo_2 ;  
   wire notCDom_reduced4SigExtra_hi_5 ;  
   wire notCDom_reduced4SigExtra_lo_4 ;  
   wire [5:0] _notCDom_reduced4SigExtra_T_10 ;  
   wire [6:0] _GEN_6 ;  
   wire [6:0] _notCDom_reduced4SigExtra_T_11 ;  
   wire notCDom_reduced4SigExtra ;  
   wire [25:0] notCDom_sig_hi ;  
   wire _notCDom_sig_T_1 ;  
   wire notCDom_sig_lo ;  
   wire [26:0] notCDom_sig ;  
   wire notCDom_completeCancellation ;  
   wire _notCDom_sign_T ;  
   wire notCDom_sign ;  
   wire notNaN_isInfProd ;  
   wire notNaN_isInfOut ;  
   wire _notNaN_addZeros_T ;  
   wire notNaN_addZeros ;  
   wire _io_invalidExc_T ;  
   wire _io_invalidExc_T_1 ;  
   wire _io_invalidExc_T_2 ;  
   wire _io_invalidExc_T_3 ;  
   wire _io_invalidExc_T_6 ;  
   wire _io_invalidExc_T_7 ;  
   wire _io_invalidExc_T_8 ;  
   wire _io_rawOut_isZero_T_1 ;  
   wire _io_rawOut_sign_T ;  
   wire _io_rawOut_sign_T_1 ;  
   wire _io_rawOut_sign_T_2 ;  
   wire _io_rawOut_sign_T_4 ;  
   wire _io_rawOut_sign_T_5 ;  
   wire _io_rawOut_sign_T_6 ;  
   wire _io_rawOut_sign_T_7 ;  
   wire _io_rawOut_sign_T_8 ;  
   wire _io_rawOut_sign_T_9 ;  
   wire _io_rawOut_sign_T_10 ;  
   wire _io_rawOut_sign_T_11 ;  
   wire _io_rawOut_sign_T_14 ;  
   wire _io_rawOut_sign_T_15 ;  
   wire _io_rawOut_sign_T_16 ;  
   wire [29:0] MulAddRecFNToRaw_postMul_covSum ;  
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign CDom_sign=io_fromPreMul_signProd^io_fromPreMul_doSubMags; 
  assign _sigSum_T_2=io_fromPreMul_highAlignedSigC+26'h1; 
  assign sigSum_hi_hi=io_mulAddResult[48] ? _sigSum_T_2:io_fromPreMul_highAlignedSigC; 
  assign sigSum_hi_lo=io_mulAddResult[47:0]; 
  assign sigSum={sigSum_hi_hi,sigSum_hi_lo,io_fromPreMul_bit0AlignedSigC}; 
  assign _CDom_sExp_T={1'b0,$signed(io_fromPreMul_doSubMags)}; 
  assign _GEN_0={{8{_CDom_sExp_T[1]}},_CDom_sExp_T}; 
  assign CDom_sExp=$signed(io_fromPreMul_sExpSum)-$signed(_GEN_0); 
  assign CDom_absSigSum_hi_lo=io_fromPreMul_highAlignedSigC[25:24]; 
  assign CDom_absSigSum_lo=sigSum[72:26]; 
  assign _CDom_absSigSum_T_2={1'h0,CDom_absSigSum_hi_lo,CDom_absSigSum_lo}; 
  assign CDom_absSigSum=io_fromPreMul_doSubMags ? ~sigSum[74:25]:_CDom_absSigSum_T_2; 
  assign _CDom_absSigSumExtra_T_2=|(~sigSum[24:1]); 
  assign _CDom_absSigSumExtra_T_4=|sigSum[25:1]; 
  assign CDom_absSigSumExtra=io_fromPreMul_doSubMags ? _CDom_absSigSumExtra_T_2:_CDom_absSigSumExtra_T_4; 
  assign _GEN_1={31'b0,CDom_absSigSum}; 
  assign _CDom_mainSig_T=_GEN_1<<io_fromPreMul_CDom_CAlignDist; 
  assign CDom_mainSig=_CDom_mainSig_T[49:21]; 
  assign _CDom_reduced4SigExtra_T_1={CDom_absSigSum[23:0],3'h0}; 
  assign CDom_reduced4SigExtra_reducedVec_0=|_CDom_reduced4SigExtra_T_1[3:0]; 
  assign CDom_reduced4SigExtra_reducedVec_1=|_CDom_reduced4SigExtra_T_1[7:4]; 
  assign CDom_reduced4SigExtra_reducedVec_2=|_CDom_reduced4SigExtra_T_1[11:8]; 
  assign CDom_reduced4SigExtra_reducedVec_3=|_CDom_reduced4SigExtra_T_1[15:12]; 
  assign CDom_reduced4SigExtra_reducedVec_4=|_CDom_reduced4SigExtra_T_1[19:16]; 
  assign CDom_reduced4SigExtra_reducedVec_5=|_CDom_reduced4SigExtra_T_1[23:20]; 
  assign CDom_reduced4SigExtra_reducedVec_6=|_CDom_reduced4SigExtra_T_1[26:24]; 
  assign _CDom_reduced4SigExtra_T_2={CDom_reduced4SigExtra_reducedVec_6,CDom_reduced4SigExtra_reducedVec_5,CDom_reduced4SigExtra_reducedVec_4,CDom_reduced4SigExtra_reducedVec_3,CDom_reduced4SigExtra_reducedVec_2,CDom_reduced4SigExtra_reducedVec_1,CDom_reduced4SigExtra_reducedVec_0}; 
  assign CDom_reduced4SigExtra_shift=-9'sh100>>>~io_fromPreMul_CDom_CAlignDist[4:2]; 
  assign CDom_reduced4SigExtra_hi_1=CDom_reduced4SigExtra_shift[1]; 
  assign CDom_reduced4SigExtra_lo_1=CDom_reduced4SigExtra_shift[2]; 
  assign CDom_reduced4SigExtra_hi_3=CDom_reduced4SigExtra_shift[3]; 
  assign CDom_reduced4SigExtra_lo_2=CDom_reduced4SigExtra_shift[4]; 
  assign CDom_reduced4SigExtra_hi_5=CDom_reduced4SigExtra_shift[5]; 
  assign CDom_reduced4SigExtra_lo_4=CDom_reduced4SigExtra_shift[6]; 
  assign _CDom_reduced4SigExtra_T_10={CDom_reduced4SigExtra_hi_1,CDom_reduced4SigExtra_lo_1,CDom_reduced4SigExtra_hi_3,CDom_reduced4SigExtra_lo_2,CDom_reduced4SigExtra_hi_5,CDom_reduced4SigExtra_lo_4}; 
  assign _GEN_2={1'b0,_CDom_reduced4SigExtra_T_10}; 
  assign _CDom_reduced4SigExtra_T_11=_CDom_reduced4SigExtra_T_2&_GEN_2; 
  assign CDom_reduced4SigExtra=|_CDom_reduced4SigExtra_T_11; 
  assign CDom_sig_hi=CDom_mainSig[28:3]; 
  assign _CDom_sig_T_1=|CDom_mainSig[2:0]; 
  assign _CDom_sig_T_2=_CDom_sig_T_1|CDom_reduced4SigExtra; 
  assign CDom_sig_lo=_CDom_sig_T_2|CDom_absSigSumExtra; 
  assign CDom_sig={CDom_sig_hi,CDom_sig_lo}; 
  assign notCDom_signSigSum=sigSum[51]; 
  assign _GEN_3={50'b0,io_fromPreMul_doSubMags}; 
  assign _notCDom_absSigSum_T_4=sigSum[50:0]+_GEN_3; 
  assign notCDom_absSigSum=notCDom_signSigSum ? ~sigSum[50:0]:_notCDom_absSigSum_T_4; 
  assign notCDom_reduced2AbsSigSum_reducedVec_0=|notCDom_absSigSum[1:0]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_1=|notCDom_absSigSum[3:2]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_2=|notCDom_absSigSum[5:4]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_3=|notCDom_absSigSum[7:6]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_4=|notCDom_absSigSum[9:8]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_5=|notCDom_absSigSum[11:10]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_6=|notCDom_absSigSum[13:12]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_7=|notCDom_absSigSum[15:14]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_8=|notCDom_absSigSum[17:16]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_9=|notCDom_absSigSum[19:18]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_10=|notCDom_absSigSum[21:20]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_11=|notCDom_absSigSum[23:22]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_12=|notCDom_absSigSum[25:24]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_13=|notCDom_absSigSum[27:26]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_14=|notCDom_absSigSum[29:28]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_15=|notCDom_absSigSum[31:30]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_16=|notCDom_absSigSum[33:32]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_17=|notCDom_absSigSum[35:34]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_18=|notCDom_absSigSum[37:36]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_19=|notCDom_absSigSum[39:38]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_20=|notCDom_absSigSum[41:40]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_21=|notCDom_absSigSum[43:42]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_22=|notCDom_absSigSum[45:44]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_23=|notCDom_absSigSum[47:46]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_24=|notCDom_absSigSum[49:48]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_25=|notCDom_absSigSum[50]; 
  assign notCDom_reduced2AbsSigSum_lo_lo={notCDom_reduced2AbsSigSum_reducedVec_5,notCDom_reduced2AbsSigSum_reducedVec_4,notCDom_reduced2AbsSigSum_reducedVec_3,notCDom_reduced2AbsSigSum_reducedVec_2,notCDom_reduced2AbsSigSum_reducedVec_1,notCDom_reduced2AbsSigSum_reducedVec_0}; 
  assign notCDom_reduced2AbsSigSum_lo={notCDom_reduced2AbsSigSum_reducedVec_12,notCDom_reduced2AbsSigSum_reducedVec_11,notCDom_reduced2AbsSigSum_reducedVec_10,notCDom_reduced2AbsSigSum_reducedVec_9,notCDom_reduced2AbsSigSum_reducedVec_8,notCDom_reduced2AbsSigSum_reducedVec_7,notCDom_reduced2AbsSigSum_reducedVec_6,notCDom_reduced2AbsSigSum_lo_lo}; 
  assign notCDom_reduced2AbsSigSum_hi_lo={notCDom_reduced2AbsSigSum_reducedVec_18,notCDom_reduced2AbsSigSum_reducedVec_17,notCDom_reduced2AbsSigSum_reducedVec_16,notCDom_reduced2AbsSigSum_reducedVec_15,notCDom_reduced2AbsSigSum_reducedVec_14,notCDom_reduced2AbsSigSum_reducedVec_13}; 
  assign notCDom_reduced2AbsSigSum={notCDom_reduced2AbsSigSum_reducedVec_25,notCDom_reduced2AbsSigSum_reducedVec_24,notCDom_reduced2AbsSigSum_reducedVec_23,notCDom_reduced2AbsSigSum_reducedVec_22,notCDom_reduced2AbsSigSum_reducedVec_21,notCDom_reduced2AbsSigSum_reducedVec_20,notCDom_reduced2AbsSigSum_reducedVec_19,notCDom_reduced2AbsSigSum_hi_lo,notCDom_reduced2AbsSigSum_lo}; 
  assign _notCDom_normDistReduced2_T_26=notCDom_reduced2AbsSigSum[1] ? 5'h18:5'h19; 
  assign _notCDom_normDistReduced2_T_27=notCDom_reduced2AbsSigSum[2] ? 5'h17:_notCDom_normDistReduced2_T_26; 
  assign _notCDom_normDistReduced2_T_28=notCDom_reduced2AbsSigSum[3] ? 5'h16:_notCDom_normDistReduced2_T_27; 
  assign _notCDom_normDistReduced2_T_29=notCDom_reduced2AbsSigSum[4] ? 5'h15:_notCDom_normDistReduced2_T_28; 
  assign _notCDom_normDistReduced2_T_30=notCDom_reduced2AbsSigSum[5] ? 5'h14:_notCDom_normDistReduced2_T_29; 
  assign _notCDom_normDistReduced2_T_31=notCDom_reduced2AbsSigSum[6] ? 5'h13:_notCDom_normDistReduced2_T_30; 
  assign _notCDom_normDistReduced2_T_32=notCDom_reduced2AbsSigSum[7] ? 5'h12:_notCDom_normDistReduced2_T_31; 
  assign _notCDom_normDistReduced2_T_33=notCDom_reduced2AbsSigSum[8] ? 5'h11:_notCDom_normDistReduced2_T_32; 
  assign _notCDom_normDistReduced2_T_34=notCDom_reduced2AbsSigSum[9] ? 5'h10:_notCDom_normDistReduced2_T_33; 
  assign _notCDom_normDistReduced2_T_35=notCDom_reduced2AbsSigSum[10] ? 5'hf:_notCDom_normDistReduced2_T_34; 
  assign _notCDom_normDistReduced2_T_36=notCDom_reduced2AbsSigSum[11] ? 5'he:_notCDom_normDistReduced2_T_35; 
  assign _notCDom_normDistReduced2_T_37=notCDom_reduced2AbsSigSum[12] ? 5'hd:_notCDom_normDistReduced2_T_36; 
  assign _notCDom_normDistReduced2_T_38=notCDom_reduced2AbsSigSum[13] ? 5'hc:_notCDom_normDistReduced2_T_37; 
  assign _notCDom_normDistReduced2_T_39=notCDom_reduced2AbsSigSum[14] ? 5'hb:_notCDom_normDistReduced2_T_38; 
  assign _notCDom_normDistReduced2_T_40=notCDom_reduced2AbsSigSum[15] ? 5'ha:_notCDom_normDistReduced2_T_39; 
  assign _notCDom_normDistReduced2_T_41=notCDom_reduced2AbsSigSum[16] ? 5'h9:_notCDom_normDistReduced2_T_40; 
  assign _notCDom_normDistReduced2_T_42=notCDom_reduced2AbsSigSum[17] ? 5'h8:_notCDom_normDistReduced2_T_41; 
  assign _notCDom_normDistReduced2_T_43=notCDom_reduced2AbsSigSum[18] ? 5'h7:_notCDom_normDistReduced2_T_42; 
  assign _notCDom_normDistReduced2_T_44=notCDom_reduced2AbsSigSum[19] ? 5'h6:_notCDom_normDistReduced2_T_43; 
  assign _notCDom_normDistReduced2_T_45=notCDom_reduced2AbsSigSum[20] ? 5'h5:_notCDom_normDistReduced2_T_44; 
  assign _notCDom_normDistReduced2_T_46=notCDom_reduced2AbsSigSum[21] ? 5'h4:_notCDom_normDistReduced2_T_45; 
  assign _notCDom_normDistReduced2_T_47=notCDom_reduced2AbsSigSum[22] ? 5'h3:_notCDom_normDistReduced2_T_46; 
  assign _notCDom_normDistReduced2_T_48=notCDom_reduced2AbsSigSum[23] ? 5'h2:_notCDom_normDistReduced2_T_47; 
  assign _notCDom_normDistReduced2_T_49=notCDom_reduced2AbsSigSum[24] ? 5'h1:_notCDom_normDistReduced2_T_48; 
  assign notCDom_normDistReduced2=notCDom_reduced2AbsSigSum[25] ? 5'h0:_notCDom_normDistReduced2_T_49; 
  assign notCDom_nearNormDist={notCDom_normDistReduced2,1'h0}; 
  assign _notCDom_sExp_T={1'b0,$signed(notCDom_nearNormDist)}; 
  assign _GEN_4={{3{_notCDom_sExp_T[6]}},_notCDom_sExp_T}; 
  assign notCDom_sExp=$signed(io_fromPreMul_sExpSum)-$signed(_GEN_4); 
  assign _GEN_5={63'b0,notCDom_absSigSum}; 
  assign _notCDom_mainSig_T=_GEN_5<<notCDom_nearNormDist; 
  assign notCDom_mainSig=_notCDom_mainSig_T[51:23]; 
  assign notCDom_reduced4SigExtra_reducedVec_0=|notCDom_reduced2AbsSigSum[1:0]; 
  assign notCDom_reduced4SigExtra_reducedVec_1=|notCDom_reduced2AbsSigSum[3:2]; 
  assign notCDom_reduced4SigExtra_reducedVec_2=|notCDom_reduced2AbsSigSum[5:4]; 
  assign notCDom_reduced4SigExtra_reducedVec_3=|notCDom_reduced2AbsSigSum[7:6]; 
  assign notCDom_reduced4SigExtra_reducedVec_4=|notCDom_reduced2AbsSigSum[9:8]; 
  assign notCDom_reduced4SigExtra_reducedVec_5=|notCDom_reduced2AbsSigSum[11:10]; 
  assign notCDom_reduced4SigExtra_reducedVec_6=|notCDom_reduced2AbsSigSum[12]; 
  assign _notCDom_reduced4SigExtra_T_2={notCDom_reduced4SigExtra_reducedVec_6,notCDom_reduced4SigExtra_reducedVec_5,notCDom_reduced4SigExtra_reducedVec_4,notCDom_reduced4SigExtra_reducedVec_3,notCDom_reduced4SigExtra_reducedVec_2,notCDom_reduced4SigExtra_reducedVec_1,notCDom_reduced4SigExtra_reducedVec_0}; 
  assign notCDom_reduced4SigExtra_shift=-17'sh10000>>>~notCDom_normDistReduced2[4:1]; 
  assign notCDom_reduced4SigExtra_hi_1=notCDom_reduced4SigExtra_shift[1]; 
  assign notCDom_reduced4SigExtra_lo_1=notCDom_reduced4SigExtra_shift[2]; 
  assign notCDom_reduced4SigExtra_hi_3=notCDom_reduced4SigExtra_shift[3]; 
  assign notCDom_reduced4SigExtra_lo_2=notCDom_reduced4SigExtra_shift[4]; 
  assign notCDom_reduced4SigExtra_hi_5=notCDom_reduced4SigExtra_shift[5]; 
  assign notCDom_reduced4SigExtra_lo_4=notCDom_reduced4SigExtra_shift[6]; 
  assign _notCDom_reduced4SigExtra_T_10={notCDom_reduced4SigExtra_hi_1,notCDom_reduced4SigExtra_lo_1,notCDom_reduced4SigExtra_hi_3,notCDom_reduced4SigExtra_lo_2,notCDom_reduced4SigExtra_hi_5,notCDom_reduced4SigExtra_lo_4}; 
  assign _GEN_6={1'b0,_notCDom_reduced4SigExtra_T_10}; 
  assign _notCDom_reduced4SigExtra_T_11=_notCDom_reduced4SigExtra_T_2&_GEN_6; 
  assign notCDom_reduced4SigExtra=|_notCDom_reduced4SigExtra_T_11; 
  assign notCDom_sig_hi=notCDom_mainSig[28:3]; 
  assign _notCDom_sig_T_1=|notCDom_mainSig[2:0]; 
  assign notCDom_sig_lo=_notCDom_sig_T_1|notCDom_reduced4SigExtra; 
  assign notCDom_sig={notCDom_sig_hi,notCDom_sig_lo}; 
  assign notCDom_completeCancellation=notCDom_sig[26:25]==2'h0; 
  assign _notCDom_sign_T=io_fromPreMul_signProd^notCDom_signSigSum; 
  assign notCDom_sign=notCDom_completeCancellation ? roundingMode_min:_notCDom_sign_T; 
  assign notNaN_isInfProd=io_fromPreMul_isInfA|io_fromPreMul_isInfB; 
  assign notNaN_isInfOut=notNaN_isInfProd|io_fromPreMul_isInfC; 
  assign _notNaN_addZeros_T=io_fromPreMul_isZeroA|io_fromPreMul_isZeroB; 
  assign notNaN_addZeros=_notNaN_addZeros_T&io_fromPreMul_isZeroC; 
  assign _io_invalidExc_T=io_fromPreMul_isInfA&io_fromPreMul_isZeroB; 
  assign _io_invalidExc_T_1=io_fromPreMul_isSigNaNAny|_io_invalidExc_T; 
  assign _io_invalidExc_T_2=io_fromPreMul_isZeroA&io_fromPreMul_isInfB; 
  assign _io_invalidExc_T_3=_io_invalidExc_T_1|_io_invalidExc_T_2; 
  assign _io_invalidExc_T_6=~io_fromPreMul_isNaNAOrB&notNaN_isInfProd; 
  assign _io_invalidExc_T_7=_io_invalidExc_T_6&io_fromPreMul_isInfC; 
  assign _io_invalidExc_T_8=_io_invalidExc_T_7&io_fromPreMul_doSubMags; 
  assign _io_rawOut_isZero_T_1=~io_fromPreMul_CIsDominant&notCDom_completeCancellation; 
  assign _io_rawOut_sign_T=notNaN_isInfProd&io_fromPreMul_signProd; 
  assign _io_rawOut_sign_T_1=io_fromPreMul_isInfC&CDom_sign; 
  assign _io_rawOut_sign_T_2=_io_rawOut_sign_T|_io_rawOut_sign_T_1; 
  assign _io_rawOut_sign_T_4=notNaN_addZeros&~roundingMode_min; 
  assign _io_rawOut_sign_T_5=_io_rawOut_sign_T_4&io_fromPreMul_signProd; 
  assign _io_rawOut_sign_T_6=_io_rawOut_sign_T_5&CDom_sign; 
  assign _io_rawOut_sign_T_7=_io_rawOut_sign_T_2|_io_rawOut_sign_T_6; 
  assign _io_rawOut_sign_T_8=notNaN_addZeros&roundingMode_min; 
  assign _io_rawOut_sign_T_9=io_fromPreMul_signProd|CDom_sign; 
  assign _io_rawOut_sign_T_10=_io_rawOut_sign_T_8&_io_rawOut_sign_T_9; 
  assign _io_rawOut_sign_T_11=_io_rawOut_sign_T_7|_io_rawOut_sign_T_10; 
  assign _io_rawOut_sign_T_14=~notNaN_isInfOut&~notNaN_addZeros; 
  assign _io_rawOut_sign_T_15=io_fromPreMul_CIsDominant ? CDom_sign:notCDom_sign; 
  assign _io_rawOut_sign_T_16=_io_rawOut_sign_T_14&_io_rawOut_sign_T_15; 
  assign io_invalidExc=_io_invalidExc_T_3|_io_invalidExc_T_8; 
  assign io_rawOut_isNaN=io_fromPreMul_isNaNAOrB|io_fromPreMul_isNaNC; 
  assign io_rawOut_isInf=notNaN_isInfProd|io_fromPreMul_isInfC; 
  assign io_rawOut_isZero=notNaN_addZeros|_io_rawOut_isZero_T_1; 
  assign io_rawOut_sign=_io_rawOut_sign_T_11|_io_rawOut_sign_T_16; 
  assign io_rawOut_sExp=io_fromPreMul_CIsDominant ? $signed(CDom_sExp):$signed(notCDom_sExp); 
  assign io_rawOut_sig=io_fromPreMul_CIsDominant ? CDom_sig:notCDom_sig; 
  assign MulAddRecFNToRaw_postMul_covSum=30'h0; 
  assign io_covSum=MulAddRecFNToRaw_postMul_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module RoundAnyRawFNToRecFN_1 (
  input io_in_isZero,
  input io_in_sign,
  input [8:0] io_in_sExp,
  input [64:0] io_in_sig,
  input [2:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundingMode_near_even ;  
   wire roundingMode_min ;  
   wire roundingMode_max ;  
   wire roundingMode_near_maxMag ;  
   wire roundingMode_odd ;  
   wire _roundMagUp_T ;  
   wire _roundMagUp_T_2 ;  
   wire roundMagUp ;  
   wire [9:0] _sAdjustedExp_T ;  
   wire [9:0] sAdjustedExp ;  
   wire [25:0] adjustedSig_hi ;  
   wire adjustedSig_lo ;  
   wire [26:0] adjustedSig ;  
   wire [26:0] _roundPosBit_T ;  
   wire roundPosBit ;  
   wire [26:0] _anyRoundExtra_T ;  
   wire anyRoundExtra ;  
   wire anyRound ;  
   wire _roundIncr_T ;  
   wire _roundIncr_T_1 ;  
   wire _roundIncr_T_2 ;  
   wire roundIncr ;  
   wire [26:0] _roundedSig_T ;  
   wire [25:0] _roundedSig_T_2 ;  
   wire _roundedSig_T_3 ;  
   wire _roundedSig_T_5 ;  
   wire [25:0] _roundedSig_T_7 ;  
   wire [25:0] _roundedSig_T_9 ;  
   wire [26:0] _roundedSig_T_11 ;  
   wire _roundedSig_T_13 ;  
   wire [25:0] _roundedSig_T_15 ;  
   wire [25:0] _GEN_0 ;  
   wire [25:0] _roundedSig_T_16 ;  
   wire [25:0] roundedSig ;  
   wire [2:0] _sRoundedExp_T_1 ;  
   wire [9:0] _GEN_1 ;  
   wire [10:0] sRoundedExp ;  
   wire [8:0] common_expOut ;  
   wire [22:0] common_fractOut ;  
   wire commonCase ;  
   wire inexact ;  
   wire [8:0] _expOut_T_1 ;  
   wire [8:0] expOut ;  
   wire [22:0] fractOut ;  
   wire [9:0] io_out_hi ;  
   wire [1:0] io_exceptionFlags_lo ;  
   wire [29:0] RoundAnyRawFNToRecFN_1_covSum ;  
  assign roundingMode_near_even=io_roundingMode==3'h0; 
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign roundingMode_max=io_roundingMode==3'h3; 
  assign roundingMode_near_maxMag=io_roundingMode==3'h4; 
  assign roundingMode_odd=io_roundingMode==3'h6; 
  assign _roundMagUp_T=roundingMode_min&io_in_sign; 
  assign _roundMagUp_T_2=roundingMode_max&~io_in_sign; 
  assign roundMagUp=_roundMagUp_T|_roundMagUp_T_2; 
  assign _sAdjustedExp_T=$signed(io_in_sExp)+9'sh80; 
  assign sAdjustedExp={1'b0,$signed(_sAdjustedExp_T[8:0])}; 
  assign adjustedSig_hi=io_in_sig[64:39]; 
  assign adjustedSig_lo=|io_in_sig[38:0]; 
  assign adjustedSig={adjustedSig_hi,adjustedSig_lo}; 
  assign _roundPosBit_T=adjustedSig&27'h2; 
  assign roundPosBit=|_roundPosBit_T; 
  assign _anyRoundExtra_T=adjustedSig&27'h1; 
  assign anyRoundExtra=|_anyRoundExtra_T; 
  assign anyRound=roundPosBit|anyRoundExtra; 
  assign _roundIncr_T=roundingMode_near_even|roundingMode_near_maxMag; 
  assign _roundIncr_T_1=_roundIncr_T&roundPosBit; 
  assign _roundIncr_T_2=roundMagUp&anyRound; 
  assign roundIncr=_roundIncr_T_1|_roundIncr_T_2; 
  assign _roundedSig_T=adjustedSig|27'h3; 
  assign _roundedSig_T_2=_roundedSig_T[26:2]+25'h1; 
  assign _roundedSig_T_3=roundingMode_near_even&roundPosBit; 
  assign _roundedSig_T_5=_roundedSig_T_3&~anyRoundExtra; 
  assign _roundedSig_T_7=_roundedSig_T_5 ? 26'h1:26'h0; 
  assign _roundedSig_T_9=_roundedSig_T_2&~_roundedSig_T_7; 
  assign _roundedSig_T_11=adjustedSig&27'h7fffffc; 
  assign _roundedSig_T_13=roundingMode_odd&anyRound; 
  assign _roundedSig_T_15=_roundedSig_T_13 ? 26'h1:26'h0; 
  assign _GEN_0={1'b0,_roundedSig_T_11[26:2]}; 
  assign _roundedSig_T_16=_GEN_0|_roundedSig_T_15; 
  assign roundedSig=roundIncr ? _roundedSig_T_9:_roundedSig_T_16; 
  assign _sRoundedExp_T_1={1'b0,$signed(roundedSig[25:24])}; 
  assign _GEN_1={{7{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; 
  assign sRoundedExp=$signed(sAdjustedExp)+$signed(_GEN_1); 
  assign common_expOut=sRoundedExp[8:0]; 
  assign common_fractOut=roundedSig[22:0]; 
  assign commonCase=~io_in_isZero; 
  assign inexact=commonCase&anyRound; 
  assign _expOut_T_1=io_in_isZero ? 9'h1c0:9'h0; 
  assign expOut=common_expOut&~_expOut_T_1; 
  assign fractOut=io_in_isZero ? 23'h0:common_fractOut; 
  assign io_out_hi={io_in_sign,expOut}; 
  assign io_exceptionFlags_lo={1'h0,inexact}; 
  assign io_out={io_out_hi,fractOut}; 
  assign io_exceptionFlags={3'h0,io_exceptionFlags_lo}; 
  assign RoundAnyRawFNToRecFN_1_covSum=30'h0; 
  assign io_covSum=RoundAnyRawFNToRecFN_1_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module RoundAnyRawFNToRecFN_2 (
  input io_in_isZero,
  input io_in_sign,
  input [8:0] io_in_sExp,
  input [64:0] io_in_sig,
  input [2:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundingMode_near_even ;  
   wire roundingMode_min ;  
   wire roundingMode_max ;  
   wire roundingMode_near_maxMag ;  
   wire roundingMode_odd ;  
   wire _roundMagUp_T ;  
   wire _roundMagUp_T_2 ;  
   wire roundMagUp ;  
   wire [11:0] _GEN_0 ;  
   wire [12:0] _sAdjustedExp_T ;  
   wire [12:0] sAdjustedExp ;  
   wire [54:0] adjustedSig_hi ;  
   wire adjustedSig_lo ;  
   wire [55:0] adjustedSig ;  
   wire [55:0] _roundPosBit_T ;  
   wire roundPosBit ;  
   wire [55:0] _anyRoundExtra_T ;  
   wire anyRoundExtra ;  
   wire anyRound ;  
   wire _roundIncr_T ;  
   wire _roundIncr_T_1 ;  
   wire _roundIncr_T_2 ;  
   wire roundIncr ;  
   wire [55:0] _roundedSig_T ;  
   wire [54:0] _roundedSig_T_2 ;  
   wire _roundedSig_T_3 ;  
   wire _roundedSig_T_5 ;  
   wire [54:0] _roundedSig_T_7 ;  
   wire [54:0] _roundedSig_T_9 ;  
   wire [55:0] _roundedSig_T_11 ;  
   wire _roundedSig_T_13 ;  
   wire [54:0] _roundedSig_T_15 ;  
   wire [54:0] _GEN_1 ;  
   wire [54:0] _roundedSig_T_16 ;  
   wire [54:0] roundedSig ;  
   wire [2:0] _sRoundedExp_T_1 ;  
   wire [12:0] _GEN_2 ;  
   wire [13:0] sRoundedExp ;  
   wire [11:0] common_expOut ;  
   wire [51:0] common_fractOut ;  
   wire commonCase ;  
   wire inexact ;  
   wire [11:0] _expOut_T_1 ;  
   wire [11:0] expOut ;  
   wire [51:0] fractOut ;  
   wire [12:0] io_out_hi ;  
   wire [1:0] io_exceptionFlags_lo ;  
   wire [29:0] RoundAnyRawFNToRecFN_2_covSum ;  
  assign roundingMode_near_even=io_roundingMode==3'h0; 
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign roundingMode_max=io_roundingMode==3'h3; 
  assign roundingMode_near_maxMag=io_roundingMode==3'h4; 
  assign roundingMode_odd=io_roundingMode==3'h6; 
  assign _roundMagUp_T=roundingMode_min&io_in_sign; 
  assign _roundMagUp_T_2=roundingMode_max&~io_in_sign; 
  assign roundMagUp=_roundMagUp_T|_roundMagUp_T_2; 
  assign _GEN_0={{3{io_in_sExp[8]}},io_in_sExp}; 
  assign _sAdjustedExp_T=$signed(_GEN_0)+12'sh780; 
  assign sAdjustedExp={1'b0,$signed(_sAdjustedExp_T[11:0])}; 
  assign adjustedSig_hi=io_in_sig[64:10]; 
  assign adjustedSig_lo=|io_in_sig[9:0]; 
  assign adjustedSig={adjustedSig_hi,adjustedSig_lo}; 
  assign _roundPosBit_T=adjustedSig&56'h2; 
  assign roundPosBit=|_roundPosBit_T; 
  assign _anyRoundExtra_T=adjustedSig&56'h1; 
  assign anyRoundExtra=|_anyRoundExtra_T; 
  assign anyRound=roundPosBit|anyRoundExtra; 
  assign _roundIncr_T=roundingMode_near_even|roundingMode_near_maxMag; 
  assign _roundIncr_T_1=_roundIncr_T&roundPosBit; 
  assign _roundIncr_T_2=roundMagUp&anyRound; 
  assign roundIncr=_roundIncr_T_1|_roundIncr_T_2; 
  assign _roundedSig_T=adjustedSig|56'h3; 
  assign _roundedSig_T_2=_roundedSig_T[55:2]+54'h1; 
  assign _roundedSig_T_3=roundingMode_near_even&roundPosBit; 
  assign _roundedSig_T_5=_roundedSig_T_3&~anyRoundExtra; 
  assign _roundedSig_T_7=_roundedSig_T_5 ? 55'h1:55'h0; 
  assign _roundedSig_T_9=_roundedSig_T_2&~_roundedSig_T_7; 
  assign _roundedSig_T_11=adjustedSig&56'hfffffffffffffc; 
  assign _roundedSig_T_13=roundingMode_odd&anyRound; 
  assign _roundedSig_T_15=_roundedSig_T_13 ? 55'h1:55'h0; 
  assign _GEN_1={1'b0,_roundedSig_T_11[55:2]}; 
  assign _roundedSig_T_16=_GEN_1|_roundedSig_T_15; 
  assign roundedSig=roundIncr ? _roundedSig_T_9:_roundedSig_T_16; 
  assign _sRoundedExp_T_1={1'b0,$signed(roundedSig[54:53])}; 
  assign _GEN_2={{10{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; 
  assign sRoundedExp=$signed(sAdjustedExp)+$signed(_GEN_2); 
  assign common_expOut=sRoundedExp[11:0]; 
  assign common_fractOut=roundedSig[51:0]; 
  assign commonCase=~io_in_isZero; 
  assign inexact=commonCase&anyRound; 
  assign _expOut_T_1=io_in_isZero ? 12'he00:12'h0; 
  assign expOut=common_expOut&~_expOut_T_1; 
  assign fractOut=io_in_isZero ? 52'h0:common_fractOut; 
  assign io_out_hi={io_in_sign,expOut}; 
  assign io_exceptionFlags_lo={1'h0,inexact}; 
  assign io_out={io_out_hi,fractOut}; 
  assign io_exceptionFlags={3'h0,io_exceptionFlags_lo}; 
  assign RoundAnyRawFNToRecFN_2_covSum=30'h0; 
  assign io_covSum=RoundAnyRawFNToRecFN_2_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module RoundAnyRawFNToRecFN_3 (
  input io_invalidExc,
  input io_in_isNaN,
  input io_in_isInf,
  input io_in_isZero,
  input io_in_sign,
  input [12:0] io_in_sExp,
  input [53:0] io_in_sig,
  input [2:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundingMode_near_even ;  
   wire roundingMode_min ;  
   wire roundingMode_max ;  
   wire roundingMode_near_maxMag ;  
   wire roundingMode_odd ;  
   wire _roundMagUp_T ;  
   wire _roundMagUp_T_2 ;  
   wire roundMagUp ;  
   wire [13:0] sAdjustedExp ;  
   wire [25:0] adjustedSig_hi ;  
   wire adjustedSig_lo ;  
   wire [26:0] adjustedSig ;  
   wire roundMask_msb ;  
   wire [7:0] roundMask_lsbs ;  
   wire roundMask_msb_1 ;  
   wire [6:0] roundMask_lsbs_1 ;  
   wire roundMask_msb_2 ;  
   wire [5:0] roundMask_lsbs_2 ;  
   wire [64:0] roundMask_shift ;  
   wire [15:0] _roundMask_T_7 ;  
   wire [15:0] _roundMask_T_9 ;  
   wire [15:0] _roundMask_T_11 ;  
   wire [15:0] _roundMask_T_12 ;  
   wire [15:0] _GEN_0 ;  
   wire [15:0] _roundMask_T_17 ;  
   wire [15:0] _roundMask_T_19 ;  
   wire [15:0] _roundMask_T_21 ;  
   wire [15:0] _roundMask_T_22 ;  
   wire [15:0] _GEN_1 ;  
   wire [15:0] _roundMask_T_27 ;  
   wire [15:0] _roundMask_T_29 ;  
   wire [15:0] _roundMask_T_31 ;  
   wire [15:0] _roundMask_T_32 ;  
   wire [15:0] _GEN_2 ;  
   wire [15:0] _roundMask_T_37 ;  
   wire [15:0] _roundMask_T_39 ;  
   wire [15:0] _roundMask_T_41 ;  
   wire [15:0] roundMask_hi ;  
   wire roundMask_hi_1 ;  
   wire roundMask_lo ;  
   wire roundMask_hi_3 ;  
   wire roundMask_lo_1 ;  
   wire roundMask_hi_5 ;  
   wire roundMask_lo_3 ;  
   wire [21:0] _roundMask_T_47 ;  
   wire [21:0] _roundMask_T_49 ;  
   wire [21:0] roundMask_hi_6 ;  
   wire [24:0] _roundMask_T_50 ;  
   wire roundMask_hi_7 ;  
   wire roundMask_lo_6 ;  
   wire roundMask_lo_7 ;  
   wire [2:0] _roundMask_T_53 ;  
   wire [2:0] _roundMask_T_54 ;  
   wire [24:0] _roundMask_T_55 ;  
   wire [24:0] roundMask_hi_9 ;  
   wire [26:0] roundMask ;  
   wire [25:0] shiftedRoundMask_lo ;  
   wire [26:0] shiftedRoundMask ;  
   wire [26:0] roundPosMask ;  
   wire [26:0] _roundPosBit_T ;  
   wire roundPosBit ;  
   wire [26:0] _anyRoundExtra_T ;  
   wire anyRoundExtra ;  
   wire anyRound ;  
   wire _roundIncr_T ;  
   wire _roundIncr_T_1 ;  
   wire _roundIncr_T_2 ;  
   wire roundIncr ;  
   wire [26:0] _roundedSig_T ;  
   wire [25:0] _roundedSig_T_2 ;  
   wire _roundedSig_T_3 ;  
   wire _roundedSig_T_5 ;  
   wire [25:0] _roundedSig_T_7 ;  
   wire [25:0] _roundedSig_T_9 ;  
   wire [26:0] _roundedSig_T_11 ;  
   wire _roundedSig_T_13 ;  
   wire [25:0] _roundedSig_T_15 ;  
   wire [25:0] _GEN_3 ;  
   wire [25:0] _roundedSig_T_16 ;  
   wire [25:0] roundedSig ;  
   wire [2:0] _sRoundedExp_T_1 ;  
   wire [13:0] _GEN_4 ;  
   wire [14:0] sRoundedExp ;  
   wire [8:0] common_expOut ;  
   wire [22:0] common_fractOut ;  
   wire [7:0] _common_overflow_T ;  
   wire common_overflow ;  
   wire common_totalUnderflow ;  
   wire unboundedRange_roundPosBit ;  
   wire unboundedRange_anyRound ;  
   wire _unboundedRange_roundIncr_T_1 ;  
   wire _unboundedRange_roundIncr_T_2 ;  
   wire unboundedRange_roundIncr ;  
   wire roundCarry ;  
   wire [5:0] _common_underflow_T ;  
   wire _common_underflow_T_1 ;  
   wire _common_underflow_T_2 ;  
   wire _common_underflow_T_6 ;  
   wire _common_underflow_T_13 ;  
   wire _common_underflow_T_14 ;  
   wire _common_underflow_T_15 ;  
   wire _common_underflow_T_17 ;  
   wire common_underflow ;  
   wire common_inexact ;  
   wire isNaNOut ;  
   wire _commonCase_T_2 ;  
   wire commonCase ;  
   wire overflow ;  
   wire underflow ;  
   wire _inexact_T ;  
   wire inexact ;  
   wire overflow_roundMagUp ;  
   wire _pegMinNonzeroMagOut_T ;  
   wire _pegMinNonzeroMagOut_T_1 ;  
   wire pegMinNonzeroMagOut ;  
   wire pegMaxFiniteMagOut ;  
   wire _notNaN_isInfOut_T ;  
   wire notNaN_isInfOut ;  
   wire signOut ;  
   wire _expOut_T ;  
   wire [8:0] _expOut_T_1 ;  
   wire [8:0] _expOut_T_3 ;  
   wire [8:0] _expOut_T_5 ;  
   wire [8:0] _expOut_T_7 ;  
   wire [8:0] _expOut_T_8 ;  
   wire [8:0] _expOut_T_10 ;  
   wire [8:0] _expOut_T_11 ;  
   wire [8:0] _expOut_T_13 ;  
   wire [8:0] _expOut_T_14 ;  
   wire [8:0] _expOut_T_15 ;  
   wire [8:0] _expOut_T_16 ;  
   wire [8:0] _expOut_T_17 ;  
   wire [8:0] _expOut_T_18 ;  
   wire [8:0] _expOut_T_19 ;  
   wire [8:0] _expOut_T_20 ;  
   wire [8:0] expOut ;  
   wire _fractOut_T ;  
   wire _fractOut_T_1 ;  
   wire [22:0] _fractOut_T_2 ;  
   wire [22:0] _fractOut_T_3 ;  
   wire [22:0] _fractOut_T_5 ;  
   wire [22:0] fractOut ;  
   wire [9:0] io_out_hi ;  
   wire [1:0] io_exceptionFlags_lo ;  
   wire [2:0] io_exceptionFlags_hi ;  
   wire [29:0] RoundAnyRawFNToRecFN_3_covSum ;  
  assign roundingMode_near_even=io_roundingMode==3'h0; 
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign roundingMode_max=io_roundingMode==3'h3; 
  assign roundingMode_near_maxMag=io_roundingMode==3'h4; 
  assign roundingMode_odd=io_roundingMode==3'h6; 
  assign _roundMagUp_T=roundingMode_min&io_in_sign; 
  assign _roundMagUp_T_2=roundingMode_max&~io_in_sign; 
  assign roundMagUp=_roundMagUp_T|_roundMagUp_T_2; 
  assign sAdjustedExp=$signed(io_in_sExp)+$signed(-13'sh700); 
  assign adjustedSig_hi=io_in_sig[53:28]; 
  assign adjustedSig_lo=|io_in_sig[27:0]; 
  assign adjustedSig={adjustedSig_hi,adjustedSig_lo}; 
  assign roundMask_msb=~sAdjustedExp[8]; 
  assign roundMask_lsbs=~sAdjustedExp[7:0]; 
  assign roundMask_msb_1=roundMask_lsbs[7]; 
  assign roundMask_lsbs_1=roundMask_lsbs[6:0]; 
  assign roundMask_msb_2=roundMask_lsbs_1[6]; 
  assign roundMask_lsbs_2=roundMask_lsbs_1[5:0]; 
  assign roundMask_shift=-65'sh10000000000000000>>>roundMask_lsbs_2; 
  assign _roundMask_T_7={8'b0,roundMask_shift[57:50]}; 
  assign _roundMask_T_9={roundMask_shift[49:42],8'h0}; 
  assign _roundMask_T_11=_roundMask_T_9&16'hff00; 
  assign _roundMask_T_12=_roundMask_T_7|_roundMask_T_11; 
  assign _GEN_0={4'b0,_roundMask_T_12[15:4]}; 
  assign _roundMask_T_17=_GEN_0&16'hf0f; 
  assign _roundMask_T_19={_roundMask_T_12[11:0],4'h0}; 
  assign _roundMask_T_21=_roundMask_T_19&16'hf0f0; 
  assign _roundMask_T_22=_roundMask_T_17|_roundMask_T_21; 
  assign _GEN_1={2'b0,_roundMask_T_22[15:2]}; 
  assign _roundMask_T_27=_GEN_1&16'h3333; 
  assign _roundMask_T_29={_roundMask_T_22[13:0],2'h0}; 
  assign _roundMask_T_31=_roundMask_T_29&16'hcccc; 
  assign _roundMask_T_32=_roundMask_T_27|_roundMask_T_31; 
  assign _GEN_2={1'b0,_roundMask_T_32[15:1]}; 
  assign _roundMask_T_37=_GEN_2&16'h5555; 
  assign _roundMask_T_39={_roundMask_T_32[14:0],1'h0}; 
  assign _roundMask_T_41=_roundMask_T_39&16'haaaa; 
  assign roundMask_hi=_roundMask_T_37|_roundMask_T_41; 
  assign roundMask_hi_1=roundMask_shift[58]; 
  assign roundMask_lo=roundMask_shift[59]; 
  assign roundMask_hi_3=roundMask_shift[60]; 
  assign roundMask_lo_1=roundMask_shift[61]; 
  assign roundMask_hi_5=roundMask_shift[62]; 
  assign roundMask_lo_3=roundMask_shift[63]; 
  assign _roundMask_T_47={roundMask_hi,roundMask_hi_1,roundMask_lo,roundMask_hi_3,roundMask_lo_1,roundMask_hi_5,roundMask_lo_3}; 
  assign _roundMask_T_49=roundMask_msb_2 ? 22'h0:~_roundMask_T_47; 
  assign roundMask_hi_6=~_roundMask_T_49; 
  assign _roundMask_T_50={roundMask_hi_6,3'h7}; 
  assign roundMask_hi_7=roundMask_shift[0]; 
  assign roundMask_lo_6=roundMask_shift[1]; 
  assign roundMask_lo_7=roundMask_shift[2]; 
  assign _roundMask_T_53={roundMask_hi_7,roundMask_lo_6,roundMask_lo_7}; 
  assign _roundMask_T_54=roundMask_msb_2 ? _roundMask_T_53:3'h0; 
  assign _roundMask_T_55=roundMask_msb_1 ? _roundMask_T_50:{22'b0,_roundMask_T_54}; 
  assign roundMask_hi_9=roundMask_msb ? _roundMask_T_55:25'h0; 
  assign roundMask={roundMask_hi_9,2'h3}; 
  assign shiftedRoundMask_lo=roundMask[26:1]; 
  assign shiftedRoundMask={1'h0,shiftedRoundMask_lo}; 
  assign roundPosMask=~shiftedRoundMask&roundMask; 
  assign _roundPosBit_T=adjustedSig&roundPosMask; 
  assign roundPosBit=|_roundPosBit_T; 
  assign _anyRoundExtra_T=adjustedSig&shiftedRoundMask; 
  assign anyRoundExtra=|_anyRoundExtra_T; 
  assign anyRound=roundPosBit|anyRoundExtra; 
  assign _roundIncr_T=roundingMode_near_even|roundingMode_near_maxMag; 
  assign _roundIncr_T_1=_roundIncr_T&roundPosBit; 
  assign _roundIncr_T_2=roundMagUp&anyRound; 
  assign roundIncr=_roundIncr_T_1|_roundIncr_T_2; 
  assign _roundedSig_T=adjustedSig|roundMask; 
  assign _roundedSig_T_2=_roundedSig_T[26:2]+25'h1; 
  assign _roundedSig_T_3=roundingMode_near_even&roundPosBit; 
  assign _roundedSig_T_5=_roundedSig_T_3&~anyRoundExtra; 
  assign _roundedSig_T_7=_roundedSig_T_5 ? shiftedRoundMask_lo:26'h0; 
  assign _roundedSig_T_9=_roundedSig_T_2&~_roundedSig_T_7; 
  assign _roundedSig_T_11=adjustedSig&~roundMask; 
  assign _roundedSig_T_13=roundingMode_odd&anyRound; 
  assign _roundedSig_T_15=_roundedSig_T_13 ? roundPosMask[26:1]:26'h0; 
  assign _GEN_3={1'b0,_roundedSig_T_11[26:2]}; 
  assign _roundedSig_T_16=_GEN_3|_roundedSig_T_15; 
  assign roundedSig=roundIncr ? _roundedSig_T_9:_roundedSig_T_16; 
  assign _sRoundedExp_T_1={1'b0,$signed(roundedSig[25:24])}; 
  assign _GEN_4={{11{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; 
  assign sRoundedExp=$signed(sAdjustedExp)+$signed(_GEN_4); 
  assign common_expOut=sRoundedExp[8:0]; 
  assign common_fractOut=roundedSig[22:0]; 
  assign _common_overflow_T=sRoundedExp[14:7]; 
  assign common_overflow=$signed(_common_overflow_T)>=8'sh3; 
  assign common_totalUnderflow=$signed(sRoundedExp)<15'sh6b; 
  assign unboundedRange_roundPosBit=adjustedSig[1]; 
  assign unboundedRange_anyRound=|adjustedSig[1:0]; 
  assign _unboundedRange_roundIncr_T_1=_roundIncr_T&unboundedRange_roundPosBit; 
  assign _unboundedRange_roundIncr_T_2=roundMagUp&unboundedRange_anyRound; 
  assign unboundedRange_roundIncr=_unboundedRange_roundIncr_T_1|_unboundedRange_roundIncr_T_2; 
  assign roundCarry=roundedSig[24]; 
  assign _common_underflow_T=sAdjustedExp[13:8]; 
  assign _common_underflow_T_1=$signed(_common_underflow_T)<=6'sh0; 
  assign _common_underflow_T_2=anyRound&_common_underflow_T_1; 
  assign _common_underflow_T_6=_common_underflow_T_2&roundMask[2]; 
  assign _common_underflow_T_13=~roundMask[3]&roundCarry; 
  assign _common_underflow_T_14=_common_underflow_T_13&roundPosBit; 
  assign _common_underflow_T_15=_common_underflow_T_14&unboundedRange_roundIncr; 
  assign _common_underflow_T_17=_common_underflow_T_6&~_common_underflow_T_15; 
  assign common_underflow=common_totalUnderflow|_common_underflow_T_17; 
  assign common_inexact=common_totalUnderflow|anyRound; 
  assign isNaNOut=io_invalidExc|io_in_isNaN; 
  assign _commonCase_T_2=~isNaNOut&~io_in_isInf; 
  assign commonCase=_commonCase_T_2&~io_in_isZero; 
  assign overflow=commonCase&common_overflow; 
  assign underflow=commonCase&common_underflow; 
  assign _inexact_T=commonCase&common_inexact; 
  assign inexact=overflow|_inexact_T; 
  assign overflow_roundMagUp=_roundIncr_T|roundMagUp; 
  assign _pegMinNonzeroMagOut_T=commonCase&common_totalUnderflow; 
  assign _pegMinNonzeroMagOut_T_1=roundMagUp|roundingMode_odd; 
  assign pegMinNonzeroMagOut=_pegMinNonzeroMagOut_T&_pegMinNonzeroMagOut_T_1; 
  assign pegMaxFiniteMagOut=overflow&~overflow_roundMagUp; 
  assign _notNaN_isInfOut_T=overflow&overflow_roundMagUp; 
  assign notNaN_isInfOut=io_in_isInf|_notNaN_isInfOut_T; 
  assign signOut=isNaNOut ? 1'h0:io_in_sign; 
  assign _expOut_T=io_in_isZero|common_totalUnderflow; 
  assign _expOut_T_1=_expOut_T ? 9'h1c0:9'h0; 
  assign _expOut_T_3=common_expOut&~_expOut_T_1; 
  assign _expOut_T_5=pegMinNonzeroMagOut ? 9'h194:9'h0; 
  assign _expOut_T_7=_expOut_T_3&~_expOut_T_5; 
  assign _expOut_T_8=pegMaxFiniteMagOut ? 9'h80:9'h0; 
  assign _expOut_T_10=_expOut_T_7&~_expOut_T_8; 
  assign _expOut_T_11=notNaN_isInfOut ? 9'h40:9'h0; 
  assign _expOut_T_13=_expOut_T_10&~_expOut_T_11; 
  assign _expOut_T_14=pegMinNonzeroMagOut ? 9'h6b:9'h0; 
  assign _expOut_T_15=_expOut_T_13|_expOut_T_14; 
  assign _expOut_T_16=pegMaxFiniteMagOut ? 9'h17f:9'h0; 
  assign _expOut_T_17=_expOut_T_15|_expOut_T_16; 
  assign _expOut_T_18=notNaN_isInfOut ? 9'h180:9'h0; 
  assign _expOut_T_19=_expOut_T_17|_expOut_T_18; 
  assign _expOut_T_20=isNaNOut ? 9'h1c0:9'h0; 
  assign expOut=_expOut_T_19|_expOut_T_20; 
  assign _fractOut_T=isNaNOut|io_in_isZero; 
  assign _fractOut_T_1=_fractOut_T|common_totalUnderflow; 
  assign _fractOut_T_2=isNaNOut ? 23'h400000:23'h0; 
  assign _fractOut_T_3=_fractOut_T_1 ? _fractOut_T_2:common_fractOut; 
  assign _fractOut_T_5=pegMaxFiniteMagOut ? 23'h7fffff:23'h0; 
  assign fractOut=_fractOut_T_3|_fractOut_T_5; 
  assign io_out_hi={signOut,expOut}; 
  assign io_exceptionFlags_lo={underflow,inexact}; 
  assign io_exceptionFlags_hi={io_invalidExc,1'h0,overflow}; 
  assign io_out={io_out_hi,fractOut}; 
  assign io_exceptionFlags={io_exceptionFlags_hi,io_exceptionFlags_lo}; 
  assign RoundAnyRawFNToRecFN_3_covSum=30'h0; 
  assign io_covSum=RoundAnyRawFNToRecFN_3_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module MulAddRecFNToRaw_preMul_1 (
  input [1:0] io_op,
  input [64:0] io_a,
  input [64:0] io_b,
  input [64:0] io_c,
  output [52:0] io_mulAddA,
  output [52:0] io_mulAddB,
  output [105:0] io_mulAddC,
  output io_toPostMul_isSigNaNAny,
  output io_toPostMul_isNaNAOrB,
  output io_toPostMul_isInfA,
  output io_toPostMul_isZeroA,
  output io_toPostMul_isInfB,
  output io_toPostMul_isZeroB,
  output io_toPostMul_signProd,
  output io_toPostMul_isNaNC,
  output io_toPostMul_isInfC,
  output io_toPostMul_isZeroC,
  output [12:0] io_toPostMul_sExpSum,
  output io_toPostMul_doSubMags,
  output io_toPostMul_CIsDominant,
  output [5:0] io_toPostMul_CDom_CAlignDist,
  output [54:0] io_toPostMul_highAlignedSigC,
  output io_toPostMul_bit0AlignedSigC,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire [11:0] rawA_exp ;  
   wire rawA_isZero ;  
   wire rawA_isSpecial ;  
   wire rawA__isNaN ;  
   wire rawA__sign ;  
   wire [12:0] rawA__sExp ;  
   wire rawA_out_sig_hi_lo ;  
   wire [51:0] rawA_out_sig_lo ;  
   wire [53:0] rawA__sig ;  
   wire [11:0] rawB_exp ;  
   wire rawB_isZero ;  
   wire rawB_isSpecial ;  
   wire rawB__isNaN ;  
   wire rawB__sign ;  
   wire [12:0] rawB__sExp ;  
   wire rawB_out_sig_hi_lo ;  
   wire [51:0] rawB_out_sig_lo ;  
   wire [53:0] rawB__sig ;  
   wire [11:0] rawC_exp ;  
   wire rawC_isZero ;  
   wire rawC_isSpecial ;  
   wire rawC__isNaN ;  
   wire rawC__sign ;  
   wire [12:0] rawC__sExp ;  
   wire rawC_out_sig_hi_lo ;  
   wire [51:0] rawC_out_sig_lo ;  
   wire [53:0] rawC__sig ;  
   wire _signProd_T ;  
   wire signProd ;  
   wire [13:0] _sExpAlignedProd_T ;  
   wire [13:0] sExpAlignedProd ;  
   wire _doSubMags_T ;  
   wire doSubMags ;  
   wire [13:0] _GEN_0 ;  
   wire [13:0] sNatCAlignDist ;  
   wire [12:0] posNatCAlignDist ;  
   wire _isMinCAlign_T ;  
   wire _isMinCAlign_T_1 ;  
   wire isMinCAlign ;  
   wire _CIsDominant_T_1 ;  
   wire _CIsDominant_T_2 ;  
   wire CIsDominant ;  
   wire _CAlignDist_T ;  
   wire [7:0] _CAlignDist_T_2 ;  
   wire [7:0] CAlignDist ;  
   wire [53:0] mainAlignedSigC_hi ;  
   wire [110:0] mainAlignedSigC_lo ;  
   wire [164:0] _mainAlignedSigC_T_3 ;  
   wire [164:0] mainAlignedSigC ;  
   wire reduced4CExtra_reducedVec_0 ;  
   wire reduced4CExtra_reducedVec_1 ;  
   wire reduced4CExtra_reducedVec_2 ;  
   wire reduced4CExtra_reducedVec_3 ;  
   wire reduced4CExtra_reducedVec_4 ;  
   wire reduced4CExtra_reducedVec_5 ;  
   wire reduced4CExtra_reducedVec_6 ;  
   wire reduced4CExtra_reducedVec_7 ;  
   wire reduced4CExtra_reducedVec_8 ;  
   wire reduced4CExtra_reducedVec_9 ;  
   wire reduced4CExtra_reducedVec_10 ;  
   wire reduced4CExtra_reducedVec_11 ;  
   wire reduced4CExtra_reducedVec_12 ;  
   wire reduced4CExtra_reducedVec_13 ;  
   wire [6:0] reduced4CExtra_lo ;  
   wire [13:0] _reduced4CExtra_T_1 ;  
   wire [64:0] reduced4CExtra_shift ;  
   wire [7:0] _reduced4CExtra_T_8 ;  
   wire [7:0] _reduced4CExtra_T_10 ;  
   wire [7:0] _reduced4CExtra_T_12 ;  
   wire [7:0] _reduced4CExtra_T_13 ;  
   wire [7:0] _GEN_1 ;  
   wire [7:0] _reduced4CExtra_T_18 ;  
   wire [7:0] _reduced4CExtra_T_20 ;  
   wire [7:0] _reduced4CExtra_T_22 ;  
   wire [7:0] _reduced4CExtra_T_23 ;  
   wire [7:0] _GEN_2 ;  
   wire [7:0] _reduced4CExtra_T_28 ;  
   wire [7:0] _reduced4CExtra_T_30 ;  
   wire [7:0] _reduced4CExtra_T_32 ;  
   wire [7:0] reduced4CExtra_hi_1 ;  
   wire reduced4CExtra_hi_2 ;  
   wire reduced4CExtra_lo_1 ;  
   wire reduced4CExtra_hi_4 ;  
   wire reduced4CExtra_lo_2 ;  
   wire reduced4CExtra_lo_4 ;  
   wire [12:0] _reduced4CExtra_T_37 ;  
   wire [13:0] _GEN_3 ;  
   wire [13:0] _reduced4CExtra_T_38 ;  
   wire reduced4CExtra ;  
   wire _alignedSigC_T_2 ;  
   wire _alignedSigC_T_4 ;  
   wire _alignedSigC_T_6 ;  
   wire _alignedSigC_T_7 ;  
   wire alignedSigC_lo ;  
   wire [161:0] alignedSigC_hi ;  
   wire [162:0] alignedSigC ;  
   wire _io_toPostMul_isSigNaNAny_T_2 ;  
   wire _io_toPostMul_isSigNaNAny_T_5 ;  
   wire _io_toPostMul_isSigNaNAny_T_6 ;  
   wire _io_toPostMul_isSigNaNAny_T_9 ;  
   wire [13:0] _io_toPostMul_sExpSum_T_2 ;  
   wire [13:0] _io_toPostMul_sExpSum_T_3 ;  
   wire [29:0] MulAddRecFNToRaw_preMul_1_covSum ;  
  assign rawA_exp=io_a[63:52]; 
  assign rawA_isZero=rawA_exp[11:9]==3'h0; 
  assign rawA_isSpecial=rawA_exp[11:10]==2'h3; 
  assign rawA__isNaN=rawA_isSpecial&rawA_exp[9]; 
  assign rawA__sign=io_a[64]; 
  assign rawA__sExp={1'b0,$signed(rawA_exp)}; 
  assign rawA_out_sig_hi_lo=~rawA_isZero; 
  assign rawA_out_sig_lo=io_a[51:0]; 
  assign rawA__sig={1'h0,rawA_out_sig_hi_lo,rawA_out_sig_lo}; 
  assign rawB_exp=io_b[63:52]; 
  assign rawB_isZero=rawB_exp[11:9]==3'h0; 
  assign rawB_isSpecial=rawB_exp[11:10]==2'h3; 
  assign rawB__isNaN=rawB_isSpecial&rawB_exp[9]; 
  assign rawB__sign=io_b[64]; 
  assign rawB__sExp={1'b0,$signed(rawB_exp)}; 
  assign rawB_out_sig_hi_lo=~rawB_isZero; 
  assign rawB_out_sig_lo=io_b[51:0]; 
  assign rawB__sig={1'h0,rawB_out_sig_hi_lo,rawB_out_sig_lo}; 
  assign rawC_exp=io_c[63:52]; 
  assign rawC_isZero=rawC_exp[11:9]==3'h0; 
  assign rawC_isSpecial=rawC_exp[11:10]==2'h3; 
  assign rawC__isNaN=rawC_isSpecial&rawC_exp[9]; 
  assign rawC__sign=io_c[64]; 
  assign rawC__sExp={1'b0,$signed(rawC_exp)}; 
  assign rawC_out_sig_hi_lo=~rawC_isZero; 
  assign rawC_out_sig_lo=io_c[51:0]; 
  assign rawC__sig={1'h0,rawC_out_sig_hi_lo,rawC_out_sig_lo}; 
  assign _signProd_T=rawA__sign^rawB__sign; 
  assign signProd=_signProd_T^io_op[1]; 
  assign _sExpAlignedProd_T=$signed(rawA__sExp)+$signed(rawB__sExp); 
  assign sExpAlignedProd=$signed(_sExpAlignedProd_T)+-14'sh7c8; 
  assign _doSubMags_T=signProd^rawC__sign; 
  assign doSubMags=_doSubMags_T^io_op[0]; 
  assign _GEN_0={{1{rawC__sExp[12]}},rawC__sExp}; 
  assign sNatCAlignDist=$signed(sExpAlignedProd)-$signed(_GEN_0); 
  assign posNatCAlignDist=sNatCAlignDist[12:0]; 
  assign _isMinCAlign_T=rawA_isZero|rawB_isZero; 
  assign _isMinCAlign_T_1=$signed(sNatCAlignDist)<14'sh0; 
  assign isMinCAlign=_isMinCAlign_T|_isMinCAlign_T_1; 
  assign _CIsDominant_T_1=posNatCAlignDist<=13'h35; 
  assign _CIsDominant_T_2=isMinCAlign|_CIsDominant_T_1; 
  assign CIsDominant=rawC_out_sig_hi_lo&_CIsDominant_T_2; 
  assign _CAlignDist_T=posNatCAlignDist<13'ha1; 
  assign _CAlignDist_T_2=_CAlignDist_T ? posNatCAlignDist[7:0]:8'ha1; 
  assign CAlignDist=isMinCAlign ? 8'h0:_CAlignDist_T_2; 
  assign mainAlignedSigC_hi=doSubMags ? ~rawC__sig:rawC__sig; 
  assign mainAlignedSigC_lo=doSubMags ? 111'h7fffffffffffffffffffffffffff:111'h0; 
  assign _mainAlignedSigC_T_3={mainAlignedSigC_hi,mainAlignedSigC_lo}; 
  assign mainAlignedSigC=$signed(_mainAlignedSigC_T_3)>>>CAlignDist; 
  assign reduced4CExtra_reducedVec_0=|rawC__sig[3:0]; 
  assign reduced4CExtra_reducedVec_1=|rawC__sig[7:4]; 
  assign reduced4CExtra_reducedVec_2=|rawC__sig[11:8]; 
  assign reduced4CExtra_reducedVec_3=|rawC__sig[15:12]; 
  assign reduced4CExtra_reducedVec_4=|rawC__sig[19:16]; 
  assign reduced4CExtra_reducedVec_5=|rawC__sig[23:20]; 
  assign reduced4CExtra_reducedVec_6=|rawC__sig[27:24]; 
  assign reduced4CExtra_reducedVec_7=|rawC__sig[31:28]; 
  assign reduced4CExtra_reducedVec_8=|rawC__sig[35:32]; 
  assign reduced4CExtra_reducedVec_9=|rawC__sig[39:36]; 
  assign reduced4CExtra_reducedVec_10=|rawC__sig[43:40]; 
  assign reduced4CExtra_reducedVec_11=|rawC__sig[47:44]; 
  assign reduced4CExtra_reducedVec_12=|rawC__sig[51:48]; 
  assign reduced4CExtra_reducedVec_13=|rawC__sig[53:52]; 
  assign reduced4CExtra_lo={reduced4CExtra_reducedVec_6,reduced4CExtra_reducedVec_5,reduced4CExtra_reducedVec_4,reduced4CExtra_reducedVec_3,reduced4CExtra_reducedVec_2,reduced4CExtra_reducedVec_1,reduced4CExtra_reducedVec_0}; 
  assign _reduced4CExtra_T_1={reduced4CExtra_reducedVec_13,reduced4CExtra_reducedVec_12,reduced4CExtra_reducedVec_11,reduced4CExtra_reducedVec_10,reduced4CExtra_reducedVec_9,reduced4CExtra_reducedVec_8,reduced4CExtra_reducedVec_7,reduced4CExtra_lo}; 
  assign reduced4CExtra_shift=-65'sh10000000000000000>>>CAlignDist[7:2]; 
  assign _reduced4CExtra_T_8={4'b0,reduced4CExtra_shift[31:28]}; 
  assign _reduced4CExtra_T_10={reduced4CExtra_shift[27:24],4'h0}; 
  assign _reduced4CExtra_T_12=_reduced4CExtra_T_10&8'hf0; 
  assign _reduced4CExtra_T_13=_reduced4CExtra_T_8|_reduced4CExtra_T_12; 
  assign _GEN_1={2'b0,_reduced4CExtra_T_13[7:2]}; 
  assign _reduced4CExtra_T_18=_GEN_1&8'h33; 
  assign _reduced4CExtra_T_20={_reduced4CExtra_T_13[5:0],2'h0}; 
  assign _reduced4CExtra_T_22=_reduced4CExtra_T_20&8'hcc; 
  assign _reduced4CExtra_T_23=_reduced4CExtra_T_18|_reduced4CExtra_T_22; 
  assign _GEN_2={1'b0,_reduced4CExtra_T_23[7:1]}; 
  assign _reduced4CExtra_T_28=_GEN_2&8'h55; 
  assign _reduced4CExtra_T_30={_reduced4CExtra_T_23[6:0],1'h0}; 
  assign _reduced4CExtra_T_32=_reduced4CExtra_T_30&8'haa; 
  assign reduced4CExtra_hi_1=_reduced4CExtra_T_28|_reduced4CExtra_T_32; 
  assign reduced4CExtra_hi_2=reduced4CExtra_shift[32]; 
  assign reduced4CExtra_lo_1=reduced4CExtra_shift[33]; 
  assign reduced4CExtra_hi_4=reduced4CExtra_shift[34]; 
  assign reduced4CExtra_lo_2=reduced4CExtra_shift[35]; 
  assign reduced4CExtra_lo_4=reduced4CExtra_shift[36]; 
  assign _reduced4CExtra_T_37={reduced4CExtra_hi_1,reduced4CExtra_hi_2,reduced4CExtra_lo_1,reduced4CExtra_hi_4,reduced4CExtra_lo_2,reduced4CExtra_lo_4}; 
  assign _GEN_3={1'b0,_reduced4CExtra_T_37}; 
  assign _reduced4CExtra_T_38=_reduced4CExtra_T_1&_GEN_3; 
  assign reduced4CExtra=|_reduced4CExtra_T_38; 
  assign _alignedSigC_T_2=&mainAlignedSigC[2:0]; 
  assign _alignedSigC_T_4=_alignedSigC_T_2&~reduced4CExtra; 
  assign _alignedSigC_T_6=|mainAlignedSigC[2:0]; 
  assign _alignedSigC_T_7=_alignedSigC_T_6|reduced4CExtra; 
  assign alignedSigC_lo=doSubMags ? _alignedSigC_T_4:_alignedSigC_T_7; 
  assign alignedSigC_hi=mainAlignedSigC[164:3]; 
  assign alignedSigC={alignedSigC_hi,alignedSigC_lo}; 
  assign _io_toPostMul_isSigNaNAny_T_2=rawA__isNaN&~rawA__sig[51]; 
  assign _io_toPostMul_isSigNaNAny_T_5=rawB__isNaN&~rawB__sig[51]; 
  assign _io_toPostMul_isSigNaNAny_T_6=_io_toPostMul_isSigNaNAny_T_2|_io_toPostMul_isSigNaNAny_T_5; 
  assign _io_toPostMul_isSigNaNAny_T_9=rawC__isNaN&~rawC__sig[51]; 
  assign _io_toPostMul_sExpSum_T_2=$signed(sExpAlignedProd)-14'sh35; 
  assign _io_toPostMul_sExpSum_T_3=CIsDominant ? $signed({{1{rawC__sExp[12]}},rawC__sExp}):$signed(_io_toPostMul_sExpSum_T_2); 
  assign io_mulAddA=rawA__sig[52:0]; 
  assign io_mulAddB=rawB__sig[52:0]; 
  assign io_mulAddC=alignedSigC[106:1]; 
  assign io_toPostMul_isSigNaNAny=_io_toPostMul_isSigNaNAny_T_6|_io_toPostMul_isSigNaNAny_T_9; 
  assign io_toPostMul_isNaNAOrB=rawA__isNaN|rawB__isNaN; 
  assign io_toPostMul_isInfA=rawA_isSpecial&~rawA_exp[9]; 
  assign io_toPostMul_isZeroA=rawA_exp[11:9]==3'h0; 
  assign io_toPostMul_isInfB=rawB_isSpecial&~rawB_exp[9]; 
  assign io_toPostMul_isZeroB=rawB_exp[11:9]==3'h0; 
  assign io_toPostMul_signProd=_signProd_T^io_op[1]; 
  assign io_toPostMul_isNaNC=rawC_isSpecial&rawC_exp[9]; 
  assign io_toPostMul_isInfC=rawC_isSpecial&~rawC_exp[9]; 
  assign io_toPostMul_isZeroC=rawC_exp[11:9]==3'h0; 
  assign io_toPostMul_sExpSum=_io_toPostMul_sExpSum_T_3[12:0]; 
  assign io_toPostMul_doSubMags=_doSubMags_T^io_op[0]; 
  assign io_toPostMul_CIsDominant=rawC_out_sig_hi_lo&_CIsDominant_T_2; 
  assign io_toPostMul_CDom_CAlignDist=CAlignDist[5:0]; 
  assign io_toPostMul_highAlignedSigC=alignedSigC[161:107]; 
  assign io_toPostMul_bit0AlignedSigC=alignedSigC[0]; 
  assign MulAddRecFNToRaw_preMul_1_covSum=30'h0; 
  assign io_covSum=MulAddRecFNToRaw_preMul_1_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module MulAddRecFNToRaw_postMul_1 (
  input io_fromPreMul_isSigNaNAny,
  input io_fromPreMul_isNaNAOrB,
  input io_fromPreMul_isInfA,
  input io_fromPreMul_isZeroA,
  input io_fromPreMul_isInfB,
  input io_fromPreMul_isZeroB,
  input io_fromPreMul_signProd,
  input io_fromPreMul_isNaNC,
  input io_fromPreMul_isInfC,
  input io_fromPreMul_isZeroC,
  input [12:0] io_fromPreMul_sExpSum,
  input io_fromPreMul_doSubMags,
  input io_fromPreMul_CIsDominant,
  input [5:0] io_fromPreMul_CDom_CAlignDist,
  input [54:0] io_fromPreMul_highAlignedSigC,
  input io_fromPreMul_bit0AlignedSigC,
  input [106:0] io_mulAddResult,
  input [2:0] io_roundingMode,
  output io_invalidExc,
  output io_rawOut_isNaN,
  output io_rawOut_isInf,
  output io_rawOut_isZero,
  output io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundingMode_min ;  
   wire CDom_sign ;  
   wire [54:0] _sigSum_T_2 ;  
   wire [54:0] sigSum_hi_hi ;  
   wire [105:0] sigSum_hi_lo ;  
   wire [161:0] sigSum ;  
   wire [1:0] _CDom_sExp_T ;  
   wire [12:0] _GEN_0 ;  
   wire [12:0] CDom_sExp ;  
   wire [1:0] CDom_absSigSum_hi_lo ;  
   wire [104:0] CDom_absSigSum_lo ;  
   wire [107:0] _CDom_absSigSum_T_2 ;  
   wire [107:0] CDom_absSigSum ;  
   wire _CDom_absSigSumExtra_T_2 ;  
   wire _CDom_absSigSumExtra_T_4 ;  
   wire CDom_absSigSumExtra ;  
   wire [170:0] _GEN_1 ;  
   wire [170:0] _CDom_mainSig_T ;  
   wire [57:0] CDom_mainSig ;  
   wire [54:0] _CDom_reduced4SigExtra_T_1 ;  
   wire CDom_reduced4SigExtra_reducedVec_0 ;  
   wire CDom_reduced4SigExtra_reducedVec_1 ;  
   wire CDom_reduced4SigExtra_reducedVec_2 ;  
   wire CDom_reduced4SigExtra_reducedVec_3 ;  
   wire CDom_reduced4SigExtra_reducedVec_4 ;  
   wire CDom_reduced4SigExtra_reducedVec_5 ;  
   wire CDom_reduced4SigExtra_reducedVec_6 ;  
   wire CDom_reduced4SigExtra_reducedVec_7 ;  
   wire CDom_reduced4SigExtra_reducedVec_8 ;  
   wire CDom_reduced4SigExtra_reducedVec_9 ;  
   wire CDom_reduced4SigExtra_reducedVec_10 ;  
   wire CDom_reduced4SigExtra_reducedVec_11 ;  
   wire CDom_reduced4SigExtra_reducedVec_12 ;  
   wire CDom_reduced4SigExtra_reducedVec_13 ;  
   wire [6:0] CDom_reduced4SigExtra_lo ;  
   wire [13:0] _CDom_reduced4SigExtra_T_2 ;  
   wire [16:0] CDom_reduced4SigExtra_shift ;  
   wire [7:0] _CDom_reduced4SigExtra_T_10 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_12 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_14 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_15 ;  
   wire [7:0] _GEN_2 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_20 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_22 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_24 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_25 ;  
   wire [7:0] _GEN_3 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_30 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_32 ;  
   wire [7:0] _CDom_reduced4SigExtra_T_34 ;  
   wire [7:0] CDom_reduced4SigExtra_hi_1 ;  
   wire CDom_reduced4SigExtra_hi_2 ;  
   wire CDom_reduced4SigExtra_lo_1 ;  
   wire CDom_reduced4SigExtra_hi_4 ;  
   wire CDom_reduced4SigExtra_lo_2 ;  
   wire CDom_reduced4SigExtra_lo_4 ;  
   wire [12:0] _CDom_reduced4SigExtra_T_39 ;  
   wire [13:0] _GEN_4 ;  
   wire [13:0] _CDom_reduced4SigExtra_T_40 ;  
   wire CDom_reduced4SigExtra ;  
   wire [54:0] CDom_sig_hi ;  
   wire _CDom_sig_T_1 ;  
   wire _CDom_sig_T_2 ;  
   wire CDom_sig_lo ;  
   wire [55:0] CDom_sig ;  
   wire notCDom_signSigSum ;  
   wire [108:0] _GEN_5 ;  
   wire [108:0] _notCDom_absSigSum_T_4 ;  
   wire [108:0] notCDom_absSigSum ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_0 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_1 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_2 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_3 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_4 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_5 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_6 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_7 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_8 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_9 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_10 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_11 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_12 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_13 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_14 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_15 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_16 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_17 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_18 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_19 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_20 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_21 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_22 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_23 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_24 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_25 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_26 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_27 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_28 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_29 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_30 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_31 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_32 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_33 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_34 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_35 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_36 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_37 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_38 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_39 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_40 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_41 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_42 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_43 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_44 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_45 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_46 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_47 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_48 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_49 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_50 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_51 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_52 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_53 ;  
   wire notCDom_reduced2AbsSigSum_reducedVec_54 ;  
   wire [5:0] notCDom_reduced2AbsSigSum_lo_lo_lo ;  
   wire [12:0] notCDom_reduced2AbsSigSum_lo_lo ;  
   wire [6:0] notCDom_reduced2AbsSigSum_lo_hi_lo ;  
   wire [26:0] notCDom_reduced2AbsSigSum_lo ;  
   wire [6:0] notCDom_reduced2AbsSigSum_hi_lo_lo ;  
   wire [13:0] notCDom_reduced2AbsSigSum_hi_lo ;  
   wire [6:0] notCDom_reduced2AbsSigSum_hi_hi_lo ;  
   wire [54:0] notCDom_reduced2AbsSigSum ;  
   wire [5:0] _notCDom_normDistReduced2_T_55 ;  
   wire [5:0] _notCDom_normDistReduced2_T_56 ;  
   wire [5:0] _notCDom_normDistReduced2_T_57 ;  
   wire [5:0] _notCDom_normDistReduced2_T_58 ;  
   wire [5:0] _notCDom_normDistReduced2_T_59 ;  
   wire [5:0] _notCDom_normDistReduced2_T_60 ;  
   wire [5:0] _notCDom_normDistReduced2_T_61 ;  
   wire [5:0] _notCDom_normDistReduced2_T_62 ;  
   wire [5:0] _notCDom_normDistReduced2_T_63 ;  
   wire [5:0] _notCDom_normDistReduced2_T_64 ;  
   wire [5:0] _notCDom_normDistReduced2_T_65 ;  
   wire [5:0] _notCDom_normDistReduced2_T_66 ;  
   wire [5:0] _notCDom_normDistReduced2_T_67 ;  
   wire [5:0] _notCDom_normDistReduced2_T_68 ;  
   wire [5:0] _notCDom_normDistReduced2_T_69 ;  
   wire [5:0] _notCDom_normDistReduced2_T_70 ;  
   wire [5:0] _notCDom_normDistReduced2_T_71 ;  
   wire [5:0] _notCDom_normDistReduced2_T_72 ;  
   wire [5:0] _notCDom_normDistReduced2_T_73 ;  
   wire [5:0] _notCDom_normDistReduced2_T_74 ;  
   wire [5:0] _notCDom_normDistReduced2_T_75 ;  
   wire [5:0] _notCDom_normDistReduced2_T_76 ;  
   wire [5:0] _notCDom_normDistReduced2_T_77 ;  
   wire [5:0] _notCDom_normDistReduced2_T_78 ;  
   wire [5:0] _notCDom_normDistReduced2_T_79 ;  
   wire [5:0] _notCDom_normDistReduced2_T_80 ;  
   wire [5:0] _notCDom_normDistReduced2_T_81 ;  
   wire [5:0] _notCDom_normDistReduced2_T_82 ;  
   wire [5:0] _notCDom_normDistReduced2_T_83 ;  
   wire [5:0] _notCDom_normDistReduced2_T_84 ;  
   wire [5:0] _notCDom_normDistReduced2_T_85 ;  
   wire [5:0] _notCDom_normDistReduced2_T_86 ;  
   wire [5:0] _notCDom_normDistReduced2_T_87 ;  
   wire [5:0] _notCDom_normDistReduced2_T_88 ;  
   wire [5:0] _notCDom_normDistReduced2_T_89 ;  
   wire [5:0] _notCDom_normDistReduced2_T_90 ;  
   wire [5:0] _notCDom_normDistReduced2_T_91 ;  
   wire [5:0] _notCDom_normDistReduced2_T_92 ;  
   wire [5:0] _notCDom_normDistReduced2_T_93 ;  
   wire [5:0] _notCDom_normDistReduced2_T_94 ;  
   wire [5:0] _notCDom_normDistReduced2_T_95 ;  
   wire [5:0] _notCDom_normDistReduced2_T_96 ;  
   wire [5:0] _notCDom_normDistReduced2_T_97 ;  
   wire [5:0] _notCDom_normDistReduced2_T_98 ;  
   wire [5:0] _notCDom_normDistReduced2_T_99 ;  
   wire [5:0] _notCDom_normDistReduced2_T_100 ;  
   wire [5:0] _notCDom_normDistReduced2_T_101 ;  
   wire [5:0] _notCDom_normDistReduced2_T_102 ;  
   wire [5:0] _notCDom_normDistReduced2_T_103 ;  
   wire [5:0] _notCDom_normDistReduced2_T_104 ;  
   wire [5:0] _notCDom_normDistReduced2_T_105 ;  
   wire [5:0] _notCDom_normDistReduced2_T_106 ;  
   wire [5:0] _notCDom_normDistReduced2_T_107 ;  
   wire [5:0] notCDom_normDistReduced2 ;  
   wire [6:0] notCDom_nearNormDist ;  
   wire [7:0] _notCDom_sExp_T ;  
   wire [12:0] _GEN_6 ;  
   wire [12:0] notCDom_sExp ;  
   wire [235:0] _GEN_7 ;  
   wire [235:0] _notCDom_mainSig_T ;  
   wire [57:0] notCDom_mainSig ;  
   wire notCDom_reduced4SigExtra_reducedVec_0 ;  
   wire notCDom_reduced4SigExtra_reducedVec_1 ;  
   wire notCDom_reduced4SigExtra_reducedVec_2 ;  
   wire notCDom_reduced4SigExtra_reducedVec_3 ;  
   wire notCDom_reduced4SigExtra_reducedVec_4 ;  
   wire notCDom_reduced4SigExtra_reducedVec_5 ;  
   wire notCDom_reduced4SigExtra_reducedVec_6 ;  
   wire notCDom_reduced4SigExtra_reducedVec_7 ;  
   wire notCDom_reduced4SigExtra_reducedVec_8 ;  
   wire notCDom_reduced4SigExtra_reducedVec_9 ;  
   wire notCDom_reduced4SigExtra_reducedVec_10 ;  
   wire notCDom_reduced4SigExtra_reducedVec_11 ;  
   wire notCDom_reduced4SigExtra_reducedVec_12 ;  
   wire notCDom_reduced4SigExtra_reducedVec_13 ;  
   wire [6:0] notCDom_reduced4SigExtra_lo ;  
   wire [13:0] _notCDom_reduced4SigExtra_T_2 ;  
   wire [32:0] notCDom_reduced4SigExtra_shift ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_10 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_12 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_14 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_15 ;  
   wire [7:0] _GEN_8 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_20 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_22 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_24 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_25 ;  
   wire [7:0] _GEN_9 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_30 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_32 ;  
   wire [7:0] _notCDom_reduced4SigExtra_T_34 ;  
   wire [7:0] notCDom_reduced4SigExtra_hi_1 ;  
   wire notCDom_reduced4SigExtra_hi_2 ;  
   wire notCDom_reduced4SigExtra_lo_1 ;  
   wire notCDom_reduced4SigExtra_hi_4 ;  
   wire notCDom_reduced4SigExtra_lo_2 ;  
   wire notCDom_reduced4SigExtra_lo_4 ;  
   wire [12:0] _notCDom_reduced4SigExtra_T_39 ;  
   wire [13:0] _GEN_10 ;  
   wire [13:0] _notCDom_reduced4SigExtra_T_40 ;  
   wire notCDom_reduced4SigExtra ;  
   wire [54:0] notCDom_sig_hi ;  
   wire _notCDom_sig_T_1 ;  
   wire notCDom_sig_lo ;  
   wire [55:0] notCDom_sig ;  
   wire notCDom_completeCancellation ;  
   wire _notCDom_sign_T ;  
   wire notCDom_sign ;  
   wire notNaN_isInfProd ;  
   wire notNaN_isInfOut ;  
   wire _notNaN_addZeros_T ;  
   wire notNaN_addZeros ;  
   wire _io_invalidExc_T ;  
   wire _io_invalidExc_T_1 ;  
   wire _io_invalidExc_T_2 ;  
   wire _io_invalidExc_T_3 ;  
   wire _io_invalidExc_T_6 ;  
   wire _io_invalidExc_T_7 ;  
   wire _io_invalidExc_T_8 ;  
   wire _io_rawOut_isZero_T_1 ;  
   wire _io_rawOut_sign_T ;  
   wire _io_rawOut_sign_T_1 ;  
   wire _io_rawOut_sign_T_2 ;  
   wire _io_rawOut_sign_T_4 ;  
   wire _io_rawOut_sign_T_5 ;  
   wire _io_rawOut_sign_T_6 ;  
   wire _io_rawOut_sign_T_7 ;  
   wire _io_rawOut_sign_T_8 ;  
   wire _io_rawOut_sign_T_9 ;  
   wire _io_rawOut_sign_T_10 ;  
   wire _io_rawOut_sign_T_11 ;  
   wire _io_rawOut_sign_T_14 ;  
   wire _io_rawOut_sign_T_15 ;  
   wire _io_rawOut_sign_T_16 ;  
   wire [29:0] MulAddRecFNToRaw_postMul_1_covSum ;  
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign CDom_sign=io_fromPreMul_signProd^io_fromPreMul_doSubMags; 
  assign _sigSum_T_2=io_fromPreMul_highAlignedSigC+55'h1; 
  assign sigSum_hi_hi=io_mulAddResult[106] ? _sigSum_T_2:io_fromPreMul_highAlignedSigC; 
  assign sigSum_hi_lo=io_mulAddResult[105:0]; 
  assign sigSum={sigSum_hi_hi,sigSum_hi_lo,io_fromPreMul_bit0AlignedSigC}; 
  assign _CDom_sExp_T={1'b0,$signed(io_fromPreMul_doSubMags)}; 
  assign _GEN_0={{11{_CDom_sExp_T[1]}},_CDom_sExp_T}; 
  assign CDom_sExp=$signed(io_fromPreMul_sExpSum)-$signed(_GEN_0); 
  assign CDom_absSigSum_hi_lo=io_fromPreMul_highAlignedSigC[54:53]; 
  assign CDom_absSigSum_lo=sigSum[159:55]; 
  assign _CDom_absSigSum_T_2={1'h0,CDom_absSigSum_hi_lo,CDom_absSigSum_lo}; 
  assign CDom_absSigSum=io_fromPreMul_doSubMags ? ~sigSum[161:54]:_CDom_absSigSum_T_2; 
  assign _CDom_absSigSumExtra_T_2=|(~sigSum[53:1]); 
  assign _CDom_absSigSumExtra_T_4=|sigSum[54:1]; 
  assign CDom_absSigSumExtra=io_fromPreMul_doSubMags ? _CDom_absSigSumExtra_T_2:_CDom_absSigSumExtra_T_4; 
  assign _GEN_1={63'b0,CDom_absSigSum}; 
  assign _CDom_mainSig_T=_GEN_1<<io_fromPreMul_CDom_CAlignDist; 
  assign CDom_mainSig=_CDom_mainSig_T[107:50]; 
  assign _CDom_reduced4SigExtra_T_1={CDom_absSigSum[52:0],2'h0}; 
  assign CDom_reduced4SigExtra_reducedVec_0=|_CDom_reduced4SigExtra_T_1[3:0]; 
  assign CDom_reduced4SigExtra_reducedVec_1=|_CDom_reduced4SigExtra_T_1[7:4]; 
  assign CDom_reduced4SigExtra_reducedVec_2=|_CDom_reduced4SigExtra_T_1[11:8]; 
  assign CDom_reduced4SigExtra_reducedVec_3=|_CDom_reduced4SigExtra_T_1[15:12]; 
  assign CDom_reduced4SigExtra_reducedVec_4=|_CDom_reduced4SigExtra_T_1[19:16]; 
  assign CDom_reduced4SigExtra_reducedVec_5=|_CDom_reduced4SigExtra_T_1[23:20]; 
  assign CDom_reduced4SigExtra_reducedVec_6=|_CDom_reduced4SigExtra_T_1[27:24]; 
  assign CDom_reduced4SigExtra_reducedVec_7=|_CDom_reduced4SigExtra_T_1[31:28]; 
  assign CDom_reduced4SigExtra_reducedVec_8=|_CDom_reduced4SigExtra_T_1[35:32]; 
  assign CDom_reduced4SigExtra_reducedVec_9=|_CDom_reduced4SigExtra_T_1[39:36]; 
  assign CDom_reduced4SigExtra_reducedVec_10=|_CDom_reduced4SigExtra_T_1[43:40]; 
  assign CDom_reduced4SigExtra_reducedVec_11=|_CDom_reduced4SigExtra_T_1[47:44]; 
  assign CDom_reduced4SigExtra_reducedVec_12=|_CDom_reduced4SigExtra_T_1[51:48]; 
  assign CDom_reduced4SigExtra_reducedVec_13=|_CDom_reduced4SigExtra_T_1[54:52]; 
  assign CDom_reduced4SigExtra_lo={CDom_reduced4SigExtra_reducedVec_6,CDom_reduced4SigExtra_reducedVec_5,CDom_reduced4SigExtra_reducedVec_4,CDom_reduced4SigExtra_reducedVec_3,CDom_reduced4SigExtra_reducedVec_2,CDom_reduced4SigExtra_reducedVec_1,CDom_reduced4SigExtra_reducedVec_0}; 
  assign _CDom_reduced4SigExtra_T_2={CDom_reduced4SigExtra_reducedVec_13,CDom_reduced4SigExtra_reducedVec_12,CDom_reduced4SigExtra_reducedVec_11,CDom_reduced4SigExtra_reducedVec_10,CDom_reduced4SigExtra_reducedVec_9,CDom_reduced4SigExtra_reducedVec_8,CDom_reduced4SigExtra_reducedVec_7,CDom_reduced4SigExtra_lo}; 
  assign CDom_reduced4SigExtra_shift=-17'sh10000>>>~io_fromPreMul_CDom_CAlignDist[5:2]; 
  assign _CDom_reduced4SigExtra_T_10={4'b0,CDom_reduced4SigExtra_shift[8:5]}; 
  assign _CDom_reduced4SigExtra_T_12={CDom_reduced4SigExtra_shift[4:1],4'h0}; 
  assign _CDom_reduced4SigExtra_T_14=_CDom_reduced4SigExtra_T_12&8'hf0; 
  assign _CDom_reduced4SigExtra_T_15=_CDom_reduced4SigExtra_T_10|_CDom_reduced4SigExtra_T_14; 
  assign _GEN_2={2'b0,_CDom_reduced4SigExtra_T_15[7:2]}; 
  assign _CDom_reduced4SigExtra_T_20=_GEN_2&8'h33; 
  assign _CDom_reduced4SigExtra_T_22={_CDom_reduced4SigExtra_T_15[5:0],2'h0}; 
  assign _CDom_reduced4SigExtra_T_24=_CDom_reduced4SigExtra_T_22&8'hcc; 
  assign _CDom_reduced4SigExtra_T_25=_CDom_reduced4SigExtra_T_20|_CDom_reduced4SigExtra_T_24; 
  assign _GEN_3={1'b0,_CDom_reduced4SigExtra_T_25[7:1]}; 
  assign _CDom_reduced4SigExtra_T_30=_GEN_3&8'h55; 
  assign _CDom_reduced4SigExtra_T_32={_CDom_reduced4SigExtra_T_25[6:0],1'h0}; 
  assign _CDom_reduced4SigExtra_T_34=_CDom_reduced4SigExtra_T_32&8'haa; 
  assign CDom_reduced4SigExtra_hi_1=_CDom_reduced4SigExtra_T_30|_CDom_reduced4SigExtra_T_34; 
  assign CDom_reduced4SigExtra_hi_2=CDom_reduced4SigExtra_shift[9]; 
  assign CDom_reduced4SigExtra_lo_1=CDom_reduced4SigExtra_shift[10]; 
  assign CDom_reduced4SigExtra_hi_4=CDom_reduced4SigExtra_shift[11]; 
  assign CDom_reduced4SigExtra_lo_2=CDom_reduced4SigExtra_shift[12]; 
  assign CDom_reduced4SigExtra_lo_4=CDom_reduced4SigExtra_shift[13]; 
  assign _CDom_reduced4SigExtra_T_39={CDom_reduced4SigExtra_hi_1,CDom_reduced4SigExtra_hi_2,CDom_reduced4SigExtra_lo_1,CDom_reduced4SigExtra_hi_4,CDom_reduced4SigExtra_lo_2,CDom_reduced4SigExtra_lo_4}; 
  assign _GEN_4={1'b0,_CDom_reduced4SigExtra_T_39}; 
  assign _CDom_reduced4SigExtra_T_40=_CDom_reduced4SigExtra_T_2&_GEN_4; 
  assign CDom_reduced4SigExtra=|_CDom_reduced4SigExtra_T_40; 
  assign CDom_sig_hi=CDom_mainSig[57:3]; 
  assign _CDom_sig_T_1=|CDom_mainSig[2:0]; 
  assign _CDom_sig_T_2=_CDom_sig_T_1|CDom_reduced4SigExtra; 
  assign CDom_sig_lo=_CDom_sig_T_2|CDom_absSigSumExtra; 
  assign CDom_sig={CDom_sig_hi,CDom_sig_lo}; 
  assign notCDom_signSigSum=sigSum[109]; 
  assign _GEN_5={108'b0,io_fromPreMul_doSubMags}; 
  assign _notCDom_absSigSum_T_4=sigSum[108:0]+_GEN_5; 
  assign notCDom_absSigSum=notCDom_signSigSum ? ~sigSum[108:0]:_notCDom_absSigSum_T_4; 
  assign notCDom_reduced2AbsSigSum_reducedVec_0=|notCDom_absSigSum[1:0]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_1=|notCDom_absSigSum[3:2]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_2=|notCDom_absSigSum[5:4]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_3=|notCDom_absSigSum[7:6]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_4=|notCDom_absSigSum[9:8]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_5=|notCDom_absSigSum[11:10]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_6=|notCDom_absSigSum[13:12]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_7=|notCDom_absSigSum[15:14]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_8=|notCDom_absSigSum[17:16]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_9=|notCDom_absSigSum[19:18]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_10=|notCDom_absSigSum[21:20]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_11=|notCDom_absSigSum[23:22]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_12=|notCDom_absSigSum[25:24]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_13=|notCDom_absSigSum[27:26]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_14=|notCDom_absSigSum[29:28]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_15=|notCDom_absSigSum[31:30]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_16=|notCDom_absSigSum[33:32]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_17=|notCDom_absSigSum[35:34]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_18=|notCDom_absSigSum[37:36]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_19=|notCDom_absSigSum[39:38]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_20=|notCDom_absSigSum[41:40]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_21=|notCDom_absSigSum[43:42]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_22=|notCDom_absSigSum[45:44]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_23=|notCDom_absSigSum[47:46]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_24=|notCDom_absSigSum[49:48]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_25=|notCDom_absSigSum[51:50]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_26=|notCDom_absSigSum[53:52]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_27=|notCDom_absSigSum[55:54]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_28=|notCDom_absSigSum[57:56]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_29=|notCDom_absSigSum[59:58]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_30=|notCDom_absSigSum[61:60]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_31=|notCDom_absSigSum[63:62]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_32=|notCDom_absSigSum[65:64]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_33=|notCDom_absSigSum[67:66]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_34=|notCDom_absSigSum[69:68]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_35=|notCDom_absSigSum[71:70]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_36=|notCDom_absSigSum[73:72]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_37=|notCDom_absSigSum[75:74]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_38=|notCDom_absSigSum[77:76]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_39=|notCDom_absSigSum[79:78]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_40=|notCDom_absSigSum[81:80]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_41=|notCDom_absSigSum[83:82]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_42=|notCDom_absSigSum[85:84]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_43=|notCDom_absSigSum[87:86]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_44=|notCDom_absSigSum[89:88]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_45=|notCDom_absSigSum[91:90]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_46=|notCDom_absSigSum[93:92]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_47=|notCDom_absSigSum[95:94]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_48=|notCDom_absSigSum[97:96]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_49=|notCDom_absSigSum[99:98]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_50=|notCDom_absSigSum[101:100]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_51=|notCDom_absSigSum[103:102]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_52=|notCDom_absSigSum[105:104]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_53=|notCDom_absSigSum[107:106]; 
  assign notCDom_reduced2AbsSigSum_reducedVec_54=|notCDom_absSigSum[108]; 
  assign notCDom_reduced2AbsSigSum_lo_lo_lo={notCDom_reduced2AbsSigSum_reducedVec_5,notCDom_reduced2AbsSigSum_reducedVec_4,notCDom_reduced2AbsSigSum_reducedVec_3,notCDom_reduced2AbsSigSum_reducedVec_2,notCDom_reduced2AbsSigSum_reducedVec_1,notCDom_reduced2AbsSigSum_reducedVec_0}; 
  assign notCDom_reduced2AbsSigSum_lo_lo={notCDom_reduced2AbsSigSum_reducedVec_12,notCDom_reduced2AbsSigSum_reducedVec_11,notCDom_reduced2AbsSigSum_reducedVec_10,notCDom_reduced2AbsSigSum_reducedVec_9,notCDom_reduced2AbsSigSum_reducedVec_8,notCDom_reduced2AbsSigSum_reducedVec_7,notCDom_reduced2AbsSigSum_reducedVec_6,notCDom_reduced2AbsSigSum_lo_lo_lo}; 
  assign notCDom_reduced2AbsSigSum_lo_hi_lo={notCDom_reduced2AbsSigSum_reducedVec_19,notCDom_reduced2AbsSigSum_reducedVec_18,notCDom_reduced2AbsSigSum_reducedVec_17,notCDom_reduced2AbsSigSum_reducedVec_16,notCDom_reduced2AbsSigSum_reducedVec_15,notCDom_reduced2AbsSigSum_reducedVec_14,notCDom_reduced2AbsSigSum_reducedVec_13}; 
  assign notCDom_reduced2AbsSigSum_lo={notCDom_reduced2AbsSigSum_reducedVec_26,notCDom_reduced2AbsSigSum_reducedVec_25,notCDom_reduced2AbsSigSum_reducedVec_24,notCDom_reduced2AbsSigSum_reducedVec_23,notCDom_reduced2AbsSigSum_reducedVec_22,notCDom_reduced2AbsSigSum_reducedVec_21,notCDom_reduced2AbsSigSum_reducedVec_20,notCDom_reduced2AbsSigSum_lo_hi_lo,notCDom_reduced2AbsSigSum_lo_lo}; 
  assign notCDom_reduced2AbsSigSum_hi_lo_lo={notCDom_reduced2AbsSigSum_reducedVec_33,notCDom_reduced2AbsSigSum_reducedVec_32,notCDom_reduced2AbsSigSum_reducedVec_31,notCDom_reduced2AbsSigSum_reducedVec_30,notCDom_reduced2AbsSigSum_reducedVec_29,notCDom_reduced2AbsSigSum_reducedVec_28,notCDom_reduced2AbsSigSum_reducedVec_27}; 
  assign notCDom_reduced2AbsSigSum_hi_lo={notCDom_reduced2AbsSigSum_reducedVec_40,notCDom_reduced2AbsSigSum_reducedVec_39,notCDom_reduced2AbsSigSum_reducedVec_38,notCDom_reduced2AbsSigSum_reducedVec_37,notCDom_reduced2AbsSigSum_reducedVec_36,notCDom_reduced2AbsSigSum_reducedVec_35,notCDom_reduced2AbsSigSum_reducedVec_34,notCDom_reduced2AbsSigSum_hi_lo_lo}; 
  assign notCDom_reduced2AbsSigSum_hi_hi_lo={notCDom_reduced2AbsSigSum_reducedVec_47,notCDom_reduced2AbsSigSum_reducedVec_46,notCDom_reduced2AbsSigSum_reducedVec_45,notCDom_reduced2AbsSigSum_reducedVec_44,notCDom_reduced2AbsSigSum_reducedVec_43,notCDom_reduced2AbsSigSum_reducedVec_42,notCDom_reduced2AbsSigSum_reducedVec_41}; 
  assign notCDom_reduced2AbsSigSum={notCDom_reduced2AbsSigSum_reducedVec_54,notCDom_reduced2AbsSigSum_reducedVec_53,notCDom_reduced2AbsSigSum_reducedVec_52,notCDom_reduced2AbsSigSum_reducedVec_51,notCDom_reduced2AbsSigSum_reducedVec_50,notCDom_reduced2AbsSigSum_reducedVec_49,notCDom_reduced2AbsSigSum_reducedVec_48,notCDom_reduced2AbsSigSum_hi_hi_lo,notCDom_reduced2AbsSigSum_hi_lo,notCDom_reduced2AbsSigSum_lo}; 
  assign _notCDom_normDistReduced2_T_55=notCDom_reduced2AbsSigSum[1] ? 6'h35:6'h36; 
  assign _notCDom_normDistReduced2_T_56=notCDom_reduced2AbsSigSum[2] ? 6'h34:_notCDom_normDistReduced2_T_55; 
  assign _notCDom_normDistReduced2_T_57=notCDom_reduced2AbsSigSum[3] ? 6'h33:_notCDom_normDistReduced2_T_56; 
  assign _notCDom_normDistReduced2_T_58=notCDom_reduced2AbsSigSum[4] ? 6'h32:_notCDom_normDistReduced2_T_57; 
  assign _notCDom_normDistReduced2_T_59=notCDom_reduced2AbsSigSum[5] ? 6'h31:_notCDom_normDistReduced2_T_58; 
  assign _notCDom_normDistReduced2_T_60=notCDom_reduced2AbsSigSum[6] ? 6'h30:_notCDom_normDistReduced2_T_59; 
  assign _notCDom_normDistReduced2_T_61=notCDom_reduced2AbsSigSum[7] ? 6'h2f:_notCDom_normDistReduced2_T_60; 
  assign _notCDom_normDistReduced2_T_62=notCDom_reduced2AbsSigSum[8] ? 6'h2e:_notCDom_normDistReduced2_T_61; 
  assign _notCDom_normDistReduced2_T_63=notCDom_reduced2AbsSigSum[9] ? 6'h2d:_notCDom_normDistReduced2_T_62; 
  assign _notCDom_normDistReduced2_T_64=notCDom_reduced2AbsSigSum[10] ? 6'h2c:_notCDom_normDistReduced2_T_63; 
  assign _notCDom_normDistReduced2_T_65=notCDom_reduced2AbsSigSum[11] ? 6'h2b:_notCDom_normDistReduced2_T_64; 
  assign _notCDom_normDistReduced2_T_66=notCDom_reduced2AbsSigSum[12] ? 6'h2a:_notCDom_normDistReduced2_T_65; 
  assign _notCDom_normDistReduced2_T_67=notCDom_reduced2AbsSigSum[13] ? 6'h29:_notCDom_normDistReduced2_T_66; 
  assign _notCDom_normDistReduced2_T_68=notCDom_reduced2AbsSigSum[14] ? 6'h28:_notCDom_normDistReduced2_T_67; 
  assign _notCDom_normDistReduced2_T_69=notCDom_reduced2AbsSigSum[15] ? 6'h27:_notCDom_normDistReduced2_T_68; 
  assign _notCDom_normDistReduced2_T_70=notCDom_reduced2AbsSigSum[16] ? 6'h26:_notCDom_normDistReduced2_T_69; 
  assign _notCDom_normDistReduced2_T_71=notCDom_reduced2AbsSigSum[17] ? 6'h25:_notCDom_normDistReduced2_T_70; 
  assign _notCDom_normDistReduced2_T_72=notCDom_reduced2AbsSigSum[18] ? 6'h24:_notCDom_normDistReduced2_T_71; 
  assign _notCDom_normDistReduced2_T_73=notCDom_reduced2AbsSigSum[19] ? 6'h23:_notCDom_normDistReduced2_T_72; 
  assign _notCDom_normDistReduced2_T_74=notCDom_reduced2AbsSigSum[20] ? 6'h22:_notCDom_normDistReduced2_T_73; 
  assign _notCDom_normDistReduced2_T_75=notCDom_reduced2AbsSigSum[21] ? 6'h21:_notCDom_normDistReduced2_T_74; 
  assign _notCDom_normDistReduced2_T_76=notCDom_reduced2AbsSigSum[22] ? 6'h20:_notCDom_normDistReduced2_T_75; 
  assign _notCDom_normDistReduced2_T_77=notCDom_reduced2AbsSigSum[23] ? 6'h1f:_notCDom_normDistReduced2_T_76; 
  assign _notCDom_normDistReduced2_T_78=notCDom_reduced2AbsSigSum[24] ? 6'h1e:_notCDom_normDistReduced2_T_77; 
  assign _notCDom_normDistReduced2_T_79=notCDom_reduced2AbsSigSum[25] ? 6'h1d:_notCDom_normDistReduced2_T_78; 
  assign _notCDom_normDistReduced2_T_80=notCDom_reduced2AbsSigSum[26] ? 6'h1c:_notCDom_normDistReduced2_T_79; 
  assign _notCDom_normDistReduced2_T_81=notCDom_reduced2AbsSigSum[27] ? 6'h1b:_notCDom_normDistReduced2_T_80; 
  assign _notCDom_normDistReduced2_T_82=notCDom_reduced2AbsSigSum[28] ? 6'h1a:_notCDom_normDistReduced2_T_81; 
  assign _notCDom_normDistReduced2_T_83=notCDom_reduced2AbsSigSum[29] ? 6'h19:_notCDom_normDistReduced2_T_82; 
  assign _notCDom_normDistReduced2_T_84=notCDom_reduced2AbsSigSum[30] ? 6'h18:_notCDom_normDistReduced2_T_83; 
  assign _notCDom_normDistReduced2_T_85=notCDom_reduced2AbsSigSum[31] ? 6'h17:_notCDom_normDistReduced2_T_84; 
  assign _notCDom_normDistReduced2_T_86=notCDom_reduced2AbsSigSum[32] ? 6'h16:_notCDom_normDistReduced2_T_85; 
  assign _notCDom_normDistReduced2_T_87=notCDom_reduced2AbsSigSum[33] ? 6'h15:_notCDom_normDistReduced2_T_86; 
  assign _notCDom_normDistReduced2_T_88=notCDom_reduced2AbsSigSum[34] ? 6'h14:_notCDom_normDistReduced2_T_87; 
  assign _notCDom_normDistReduced2_T_89=notCDom_reduced2AbsSigSum[35] ? 6'h13:_notCDom_normDistReduced2_T_88; 
  assign _notCDom_normDistReduced2_T_90=notCDom_reduced2AbsSigSum[36] ? 6'h12:_notCDom_normDistReduced2_T_89; 
  assign _notCDom_normDistReduced2_T_91=notCDom_reduced2AbsSigSum[37] ? 6'h11:_notCDom_normDistReduced2_T_90; 
  assign _notCDom_normDistReduced2_T_92=notCDom_reduced2AbsSigSum[38] ? 6'h10:_notCDom_normDistReduced2_T_91; 
  assign _notCDom_normDistReduced2_T_93=notCDom_reduced2AbsSigSum[39] ? 6'hf:_notCDom_normDistReduced2_T_92; 
  assign _notCDom_normDistReduced2_T_94=notCDom_reduced2AbsSigSum[40] ? 6'he:_notCDom_normDistReduced2_T_93; 
  assign _notCDom_normDistReduced2_T_95=notCDom_reduced2AbsSigSum[41] ? 6'hd:_notCDom_normDistReduced2_T_94; 
  assign _notCDom_normDistReduced2_T_96=notCDom_reduced2AbsSigSum[42] ? 6'hc:_notCDom_normDistReduced2_T_95; 
  assign _notCDom_normDistReduced2_T_97=notCDom_reduced2AbsSigSum[43] ? 6'hb:_notCDom_normDistReduced2_T_96; 
  assign _notCDom_normDistReduced2_T_98=notCDom_reduced2AbsSigSum[44] ? 6'ha:_notCDom_normDistReduced2_T_97; 
  assign _notCDom_normDistReduced2_T_99=notCDom_reduced2AbsSigSum[45] ? 6'h9:_notCDom_normDistReduced2_T_98; 
  assign _notCDom_normDistReduced2_T_100=notCDom_reduced2AbsSigSum[46] ? 6'h8:_notCDom_normDistReduced2_T_99; 
  assign _notCDom_normDistReduced2_T_101=notCDom_reduced2AbsSigSum[47] ? 6'h7:_notCDom_normDistReduced2_T_100; 
  assign _notCDom_normDistReduced2_T_102=notCDom_reduced2AbsSigSum[48] ? 6'h6:_notCDom_normDistReduced2_T_101; 
  assign _notCDom_normDistReduced2_T_103=notCDom_reduced2AbsSigSum[49] ? 6'h5:_notCDom_normDistReduced2_T_102; 
  assign _notCDom_normDistReduced2_T_104=notCDom_reduced2AbsSigSum[50] ? 6'h4:_notCDom_normDistReduced2_T_103; 
  assign _notCDom_normDistReduced2_T_105=notCDom_reduced2AbsSigSum[51] ? 6'h3:_notCDom_normDistReduced2_T_104; 
  assign _notCDom_normDistReduced2_T_106=notCDom_reduced2AbsSigSum[52] ? 6'h2:_notCDom_normDistReduced2_T_105; 
  assign _notCDom_normDistReduced2_T_107=notCDom_reduced2AbsSigSum[53] ? 6'h1:_notCDom_normDistReduced2_T_106; 
  assign notCDom_normDistReduced2=notCDom_reduced2AbsSigSum[54] ? 6'h0:_notCDom_normDistReduced2_T_107; 
  assign notCDom_nearNormDist={notCDom_normDistReduced2,1'h0}; 
  assign _notCDom_sExp_T={1'b0,$signed(notCDom_nearNormDist)}; 
  assign _GEN_6={{5{_notCDom_sExp_T[7]}},_notCDom_sExp_T}; 
  assign notCDom_sExp=$signed(io_fromPreMul_sExpSum)-$signed(_GEN_6); 
  assign _GEN_7={127'b0,notCDom_absSigSum}; 
  assign _notCDom_mainSig_T=_GEN_7<<notCDom_nearNormDist; 
  assign notCDom_mainSig=_notCDom_mainSig_T[109:52]; 
  assign notCDom_reduced4SigExtra_reducedVec_0=|notCDom_reduced2AbsSigSum[1:0]; 
  assign notCDom_reduced4SigExtra_reducedVec_1=|notCDom_reduced2AbsSigSum[3:2]; 
  assign notCDom_reduced4SigExtra_reducedVec_2=|notCDom_reduced2AbsSigSum[5:4]; 
  assign notCDom_reduced4SigExtra_reducedVec_3=|notCDom_reduced2AbsSigSum[7:6]; 
  assign notCDom_reduced4SigExtra_reducedVec_4=|notCDom_reduced2AbsSigSum[9:8]; 
  assign notCDom_reduced4SigExtra_reducedVec_5=|notCDom_reduced2AbsSigSum[11:10]; 
  assign notCDom_reduced4SigExtra_reducedVec_6=|notCDom_reduced2AbsSigSum[13:12]; 
  assign notCDom_reduced4SigExtra_reducedVec_7=|notCDom_reduced2AbsSigSum[15:14]; 
  assign notCDom_reduced4SigExtra_reducedVec_8=|notCDom_reduced2AbsSigSum[17:16]; 
  assign notCDom_reduced4SigExtra_reducedVec_9=|notCDom_reduced2AbsSigSum[19:18]; 
  assign notCDom_reduced4SigExtra_reducedVec_10=|notCDom_reduced2AbsSigSum[21:20]; 
  assign notCDom_reduced4SigExtra_reducedVec_11=|notCDom_reduced2AbsSigSum[23:22]; 
  assign notCDom_reduced4SigExtra_reducedVec_12=|notCDom_reduced2AbsSigSum[25:24]; 
  assign notCDom_reduced4SigExtra_reducedVec_13=|notCDom_reduced2AbsSigSum[26]; 
  assign notCDom_reduced4SigExtra_lo={notCDom_reduced4SigExtra_reducedVec_6,notCDom_reduced4SigExtra_reducedVec_5,notCDom_reduced4SigExtra_reducedVec_4,notCDom_reduced4SigExtra_reducedVec_3,notCDom_reduced4SigExtra_reducedVec_2,notCDom_reduced4SigExtra_reducedVec_1,notCDom_reduced4SigExtra_reducedVec_0}; 
  assign _notCDom_reduced4SigExtra_T_2={notCDom_reduced4SigExtra_reducedVec_13,notCDom_reduced4SigExtra_reducedVec_12,notCDom_reduced4SigExtra_reducedVec_11,notCDom_reduced4SigExtra_reducedVec_10,notCDom_reduced4SigExtra_reducedVec_9,notCDom_reduced4SigExtra_reducedVec_8,notCDom_reduced4SigExtra_reducedVec_7,notCDom_reduced4SigExtra_lo}; 
  assign notCDom_reduced4SigExtra_shift=-33'sh100000000>>>~notCDom_normDistReduced2[5:1]; 
  assign _notCDom_reduced4SigExtra_T_10={4'b0,notCDom_reduced4SigExtra_shift[8:5]}; 
  assign _notCDom_reduced4SigExtra_T_12={notCDom_reduced4SigExtra_shift[4:1],4'h0}; 
  assign _notCDom_reduced4SigExtra_T_14=_notCDom_reduced4SigExtra_T_12&8'hf0; 
  assign _notCDom_reduced4SigExtra_T_15=_notCDom_reduced4SigExtra_T_10|_notCDom_reduced4SigExtra_T_14; 
  assign _GEN_8={2'b0,_notCDom_reduced4SigExtra_T_15[7:2]}; 
  assign _notCDom_reduced4SigExtra_T_20=_GEN_8&8'h33; 
  assign _notCDom_reduced4SigExtra_T_22={_notCDom_reduced4SigExtra_T_15[5:0],2'h0}; 
  assign _notCDom_reduced4SigExtra_T_24=_notCDom_reduced4SigExtra_T_22&8'hcc; 
  assign _notCDom_reduced4SigExtra_T_25=_notCDom_reduced4SigExtra_T_20|_notCDom_reduced4SigExtra_T_24; 
  assign _GEN_9={1'b0,_notCDom_reduced4SigExtra_T_25[7:1]}; 
  assign _notCDom_reduced4SigExtra_T_30=_GEN_9&8'h55; 
  assign _notCDom_reduced4SigExtra_T_32={_notCDom_reduced4SigExtra_T_25[6:0],1'h0}; 
  assign _notCDom_reduced4SigExtra_T_34=_notCDom_reduced4SigExtra_T_32&8'haa; 
  assign notCDom_reduced4SigExtra_hi_1=_notCDom_reduced4SigExtra_T_30|_notCDom_reduced4SigExtra_T_34; 
  assign notCDom_reduced4SigExtra_hi_2=notCDom_reduced4SigExtra_shift[9]; 
  assign notCDom_reduced4SigExtra_lo_1=notCDom_reduced4SigExtra_shift[10]; 
  assign notCDom_reduced4SigExtra_hi_4=notCDom_reduced4SigExtra_shift[11]; 
  assign notCDom_reduced4SigExtra_lo_2=notCDom_reduced4SigExtra_shift[12]; 
  assign notCDom_reduced4SigExtra_lo_4=notCDom_reduced4SigExtra_shift[13]; 
  assign _notCDom_reduced4SigExtra_T_39={notCDom_reduced4SigExtra_hi_1,notCDom_reduced4SigExtra_hi_2,notCDom_reduced4SigExtra_lo_1,notCDom_reduced4SigExtra_hi_4,notCDom_reduced4SigExtra_lo_2,notCDom_reduced4SigExtra_lo_4}; 
  assign _GEN_10={1'b0,_notCDom_reduced4SigExtra_T_39}; 
  assign _notCDom_reduced4SigExtra_T_40=_notCDom_reduced4SigExtra_T_2&_GEN_10; 
  assign notCDom_reduced4SigExtra=|_notCDom_reduced4SigExtra_T_40; 
  assign notCDom_sig_hi=notCDom_mainSig[57:3]; 
  assign _notCDom_sig_T_1=|notCDom_mainSig[2:0]; 
  assign notCDom_sig_lo=_notCDom_sig_T_1|notCDom_reduced4SigExtra; 
  assign notCDom_sig={notCDom_sig_hi,notCDom_sig_lo}; 
  assign notCDom_completeCancellation=notCDom_sig[55:54]==2'h0; 
  assign _notCDom_sign_T=io_fromPreMul_signProd^notCDom_signSigSum; 
  assign notCDom_sign=notCDom_completeCancellation ? roundingMode_min:_notCDom_sign_T; 
  assign notNaN_isInfProd=io_fromPreMul_isInfA|io_fromPreMul_isInfB; 
  assign notNaN_isInfOut=notNaN_isInfProd|io_fromPreMul_isInfC; 
  assign _notNaN_addZeros_T=io_fromPreMul_isZeroA|io_fromPreMul_isZeroB; 
  assign notNaN_addZeros=_notNaN_addZeros_T&io_fromPreMul_isZeroC; 
  assign _io_invalidExc_T=io_fromPreMul_isInfA&io_fromPreMul_isZeroB; 
  assign _io_invalidExc_T_1=io_fromPreMul_isSigNaNAny|_io_invalidExc_T; 
  assign _io_invalidExc_T_2=io_fromPreMul_isZeroA&io_fromPreMul_isInfB; 
  assign _io_invalidExc_T_3=_io_invalidExc_T_1|_io_invalidExc_T_2; 
  assign _io_invalidExc_T_6=~io_fromPreMul_isNaNAOrB&notNaN_isInfProd; 
  assign _io_invalidExc_T_7=_io_invalidExc_T_6&io_fromPreMul_isInfC; 
  assign _io_invalidExc_T_8=_io_invalidExc_T_7&io_fromPreMul_doSubMags; 
  assign _io_rawOut_isZero_T_1=~io_fromPreMul_CIsDominant&notCDom_completeCancellation; 
  assign _io_rawOut_sign_T=notNaN_isInfProd&io_fromPreMul_signProd; 
  assign _io_rawOut_sign_T_1=io_fromPreMul_isInfC&CDom_sign; 
  assign _io_rawOut_sign_T_2=_io_rawOut_sign_T|_io_rawOut_sign_T_1; 
  assign _io_rawOut_sign_T_4=notNaN_addZeros&~roundingMode_min; 
  assign _io_rawOut_sign_T_5=_io_rawOut_sign_T_4&io_fromPreMul_signProd; 
  assign _io_rawOut_sign_T_6=_io_rawOut_sign_T_5&CDom_sign; 
  assign _io_rawOut_sign_T_7=_io_rawOut_sign_T_2|_io_rawOut_sign_T_6; 
  assign _io_rawOut_sign_T_8=notNaN_addZeros&roundingMode_min; 
  assign _io_rawOut_sign_T_9=io_fromPreMul_signProd|CDom_sign; 
  assign _io_rawOut_sign_T_10=_io_rawOut_sign_T_8&_io_rawOut_sign_T_9; 
  assign _io_rawOut_sign_T_11=_io_rawOut_sign_T_7|_io_rawOut_sign_T_10; 
  assign _io_rawOut_sign_T_14=~notNaN_isInfOut&~notNaN_addZeros; 
  assign _io_rawOut_sign_T_15=io_fromPreMul_CIsDominant ? CDom_sign:notCDom_sign; 
  assign _io_rawOut_sign_T_16=_io_rawOut_sign_T_14&_io_rawOut_sign_T_15; 
  assign io_invalidExc=_io_invalidExc_T_3|_io_invalidExc_T_8; 
  assign io_rawOut_isNaN=io_fromPreMul_isNaNAOrB|io_fromPreMul_isNaNC; 
  assign io_rawOut_isInf=notNaN_isInfProd|io_fromPreMul_isInfC; 
  assign io_rawOut_isZero=notNaN_addZeros|_io_rawOut_isZero_T_1; 
  assign io_rawOut_sign=_io_rawOut_sign_T_11|_io_rawOut_sign_T_16; 
  assign io_rawOut_sExp=io_fromPreMul_CIsDominant ? $signed(CDom_sExp):$signed(notCDom_sExp); 
  assign io_rawOut_sig=io_fromPreMul_CIsDominant ? CDom_sig:notCDom_sig; 
  assign MulAddRecFNToRaw_postMul_1_covSum=30'h0; 
  assign io_covSum=MulAddRecFNToRaw_postMul_1_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module DivSqrtRawFN_small (
  input clock,
  input reset,
  output io_inReady,
  input io_inValid,
  input io_sqrtOp,
  input io_a_isNaN,
  input io_a_isInf,
  input io_a_isZero,
  input io_a_sign,
  input [9:0] io_a_sExp,
  input [24:0] io_a_sig,
  input io_b_isNaN,
  input io_b_isInf,
  input io_b_isZero,
  input io_b_sign,
  input [9:0] io_b_sExp,
  input [24:0] io_b_sig,
  input [2:0] io_roundingMode,
  output io_rawOutValid_div,
  output io_rawOutValid_sqrt,
  output [2:0] io_roundingModeOut,
  output io_invalidExc,
  output io_infiniteExc,
  output io_rawOut_isNaN,
  output io_rawOut_isInf,
  output io_rawOut_isZero,
  output io_rawOut_sign,
  output [9:0] io_rawOut_sExp,
  output [26:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg [26:0] cycleNum ;  
   reg [31:0] _RAND_0 ;  
   reg sqrtOp_Z ;  
   reg [31:0] _RAND_1 ;  
   reg majorExc_Z ;  
   reg [31:0] _RAND_2 ;  
   reg isNaN_Z ;  
   reg [31:0] _RAND_3 ;  
   reg isInf_Z ;  
   reg [31:0] _RAND_4 ;  
   reg isZero_Z ;  
   reg [31:0] _RAND_5 ;  
   reg sign_Z ;  
   reg [31:0] _RAND_6 ;  
   reg [9:0] sExp_Z ;  
   reg [31:0] _RAND_7 ;  
   reg [22:0] fractB_Z ;  
   reg [31:0] _RAND_8 ;  
   reg [2:0] roundingMode_Z ;  
   reg [31:0] _RAND_9 ;  
   reg [25:0] rem_Z ;  
   reg [31:0] _RAND_10 ;  
   reg notZeroRem_Z ;  
   reg [31:0] _RAND_11 ;  
   reg [25:0] sigX_Z ;  
   reg [31:0] _RAND_12 ;  
   wire _notSigNaNIn_invalidExc_S_div_T ;  
   wire _notSigNaNIn_invalidExc_S_div_T_1 ;  
   wire notSigNaNIn_invalidExc_S_div ;  
   wire _notSigNaNIn_invalidExc_S_sqrt_T_2 ;  
   wire notSigNaNIn_invalidExc_S_sqrt ;  
   wire _majorExc_S_T_2 ;  
   wire _majorExc_S_T_3 ;  
   wire _majorExc_S_T_9 ;  
   wire _majorExc_S_T_10 ;  
   wire _majorExc_S_T_11 ;  
   wire _majorExc_S_T_14 ;  
   wire _majorExc_S_T_15 ;  
   wire _majorExc_S_T_16 ;  
   wire _isNaN_S_T ;  
   wire _isNaN_S_T_1 ;  
   wire _isNaN_S_T_2 ;  
   wire _isInf_S_T ;  
   wire _isZero_S_T ;  
   wire _sign_S_T_1 ;  
   wire sign_S ;  
   wire _specialCaseA_S_T ;  
   wire specialCaseA_S ;  
   wire _specialCaseB_S_T ;  
   wire specialCaseB_S ;  
   wire normalCase_S_div ;  
   wire normalCase_S_sqrt ;  
   wire normalCase_S ;  
   wire sExpQuot_S_div_hi ;  
   wire [7:0] sExpQuot_S_div_lo ;  
   wire [8:0] _sExpQuot_S_div_T_2 ;  
   wire [9:0] _GEN_13 ;  
   wire [10:0] sExpQuot_S_div ;  
   wire _sSatExpQuot_S_div_T ;  
   wire [3:0] sSatExpQuot_S_div_hi ;  
   wire [5:0] sSatExpQuot_S_div_lo ;  
   wire [9:0] sSatExpQuot_S_div ;  
   wire evenSqrt_S ;  
   wire oddSqrt_S ;  
   wire idle ;  
   wire inReady ;  
   wire entering ;  
   wire entering_normalCase ;  
   wire skipCycle2 ;  
   wire _T_1 ;  
   wire _cycleNum_T_1 ;  
   wire [1:0] _cycleNum_T_2 ;  
   wire [25:0] _cycleNum_T_4 ;  
   wire [26:0] _cycleNum_T_5 ;  
   wire [26:0] _cycleNum_T_6 ;  
   wire [26:0] _GEN_14 ;  
   wire [26:0] _cycleNum_T_7 ;  
   wire _cycleNum_T_10 ;  
   wire [25:0] _cycleNum_T_12 ;  
   wire [26:0] _GEN_15 ;  
   wire [26:0] _cycleNum_T_13 ;  
   wire [1:0] _cycleNum_T_14 ;  
   wire [26:0] _GEN_16 ;  
   wire [26:0] _cycleNum_T_15 ;  
   wire [8:0] _sExp_Z_T ;  
   wire [9:0] _sExp_Z_T_1 ;  
   wire _T_3 ;  
   wire _rem_T_1 ;  
   wire [25:0] _rem_T_2 ;  
   wire [25:0] _rem_T_3 ;  
   wire _rem_T_4 ;  
   wire [1:0] rem_hi ;  
   wire [24:0] rem_lo ;  
   wire [26:0] _rem_T_8 ;  
   wire [26:0] _rem_T_9 ;  
   wire [26:0] _GEN_17 ;  
   wire [26:0] _rem_T_10 ;  
   wire [26:0] _rem_T_12 ;  
   wire [26:0] _rem_T_13 ;  
   wire [26:0] rem ;  
   wire [24:0] bitMask ;  
   wire _trialTerm_T_1 ;  
   wire [25:0] _trialTerm_T_2 ;  
   wire [25:0] _trialTerm_T_3 ;  
   wire _trialTerm_T_4 ;  
   wire [24:0] _trialTerm_T_5 ;  
   wire [25:0] _GEN_18 ;  
   wire [25:0] _trialTerm_T_6 ;  
   wire [25:0] _trialTerm_T_8 ;  
   wire [25:0] _trialTerm_T_9 ;  
   wire _trialTerm_T_12 ;  
   wire [23:0] _trialTerm_T_13 ;  
   wire [24:0] _trialTerm_T_14 ;  
   wire [24:0] _trialTerm_T_15 ;  
   wire [25:0] _GEN_19 ;  
   wire [25:0] _trialTerm_T_16 ;  
   wire _trialTerm_T_18 ;  
   wire [26:0] _trialTerm_T_19 ;  
   wire [26:0] _GEN_20 ;  
   wire [26:0] _trialTerm_T_20 ;  
   wire [26:0] _trialTerm_T_21 ;  
   wire [26:0] _GEN_21 ;  
   wire [26:0] trialTerm ;  
   wire [27:0] _trialRem_T ;  
   wire [27:0] _trialRem_T_1 ;  
   wire [27:0] trialRem ;  
   wire newBit ;  
   wire _T_5 ;  
   wire _T_7 ;  
   wire [27:0] _rem_Z_T ;  
   wire [27:0] _rem_Z_T_1 ;  
   wire [27:0] _GEN_10 ;  
   wire _T_9 ;  
   wire _T_10 ;  
   wire _notZeroRem_Z_T ;  
   wire [25:0] _sigX_Z_T_2 ;  
   wire [25:0] _sigX_Z_T_3 ;  
   wire _sigX_Z_T_4 ;  
   wire [24:0] _sigX_Z_T_5 ;  
   wire [25:0] _GEN_22 ;  
   wire [25:0] _sigX_Z_T_6 ;  
   wire [23:0] _sigX_Z_T_8 ;  
   wire [23:0] _sigX_Z_T_9 ;  
   wire [25:0] _GEN_23 ;  
   wire [25:0] _sigX_Z_T_10 ;  
   wire [25:0] _GEN_24 ;  
   wire [25:0] _sigX_Z_T_12 ;  
   wire [25:0] _sigX_Z_T_13 ;  
   wire [25:0] _sigX_Z_T_14 ;  
   wire [26:0] _GEN_25 ;  
   reg [4:0] DivSqrtRawFN_small_state ;  
   reg [31:0] _RAND_13 ;  
   reg DivSqrtRawFN_small_cov[0:31] ;  
   reg [31:0] _RAND_14 ;  
   wire DivSqrtRawFN_small_cov_read_data ;  
   wire [4:0] DivSqrtRawFN_small_cov_read_addr ;  
   wire DivSqrtRawFN_small_cov_write_data ;  
   wire [4:0] DivSqrtRawFN_small_cov_write_addr ;  
   wire DivSqrtRawFN_small_cov_write_mask ;  
   wire DivSqrtRawFN_small_cov_write_en ;  
   reg [29:0] DivSqrtRawFN_small_covSum ;  
   reg [31:0] _RAND_15 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire sqrtOp_Z_shl ;  
   wire [4:0] sqrtOp_Z_pad ;  
   wire [1:0] mux_cond_0_shl ;  
   wire [4:0] mux_cond_0_pad ;  
   wire [2:0] mux_cond_1_shl ;  
   wire [4:0] mux_cond_1_pad ;  
   wire [3:0] mux_cond_2_shl ;  
   wire [4:0] mux_cond_2_pad ;  
   wire [4:0] mux_cond_3_shl ;  
   wire [4:0] mux_cond_3_pad ;  
   wire [4:0] DivSqrtRawFN_small_xor1 ;  
   wire [4:0] DivSqrtRawFN_small_xor6 ;  
   wire [4:0] DivSqrtRawFN_small_xor2 ;  
   wire [4:0] DivSqrtRawFN_small_xor0 ;  
  assign _notSigNaNIn_invalidExc_S_div_T=io_a_isZero&io_b_isZero; 
  assign _notSigNaNIn_invalidExc_S_div_T_1=io_a_isInf&io_b_isInf; 
  assign notSigNaNIn_invalidExc_S_div=_notSigNaNIn_invalidExc_S_div_T|_notSigNaNIn_invalidExc_S_div_T_1; 
  assign _notSigNaNIn_invalidExc_S_sqrt_T_2=~io_a_isNaN&~io_a_isZero; 
  assign notSigNaNIn_invalidExc_S_sqrt=_notSigNaNIn_invalidExc_S_sqrt_T_2&io_a_sign; 
  assign _majorExc_S_T_2=io_a_isNaN&~io_a_sig[22]; 
  assign _majorExc_S_T_3=_majorExc_S_T_2|notSigNaNIn_invalidExc_S_sqrt; 
  assign _majorExc_S_T_9=io_b_isNaN&~io_b_sig[22]; 
  assign _majorExc_S_T_10=_majorExc_S_T_2|_majorExc_S_T_9; 
  assign _majorExc_S_T_11=_majorExc_S_T_10|notSigNaNIn_invalidExc_S_div; 
  assign _majorExc_S_T_14=~io_a_isNaN&~io_a_isInf; 
  assign _majorExc_S_T_15=_majorExc_S_T_14&io_b_isZero; 
  assign _majorExc_S_T_16=_majorExc_S_T_11|_majorExc_S_T_15; 
  assign _isNaN_S_T=io_a_isNaN|notSigNaNIn_invalidExc_S_sqrt; 
  assign _isNaN_S_T_1=io_a_isNaN|io_b_isNaN; 
  assign _isNaN_S_T_2=_isNaN_S_T_1|notSigNaNIn_invalidExc_S_div; 
  assign _isInf_S_T=io_a_isInf|io_b_isZero; 
  assign _isZero_S_T=io_a_isZero|io_b_isInf; 
  assign _sign_S_T_1=~io_sqrtOp&io_b_sign; 
  assign sign_S=io_a_sign^_sign_S_T_1; 
  assign _specialCaseA_S_T=io_a_isNaN|io_a_isInf; 
  assign specialCaseA_S=_specialCaseA_S_T|io_a_isZero; 
  assign _specialCaseB_S_T=io_b_isNaN|io_b_isInf; 
  assign specialCaseB_S=_specialCaseB_S_T|io_b_isZero; 
  assign normalCase_S_div=~specialCaseA_S&~specialCaseB_S; 
  assign normalCase_S_sqrt=~specialCaseA_S&~io_a_sign; 
  assign normalCase_S=io_sqrtOp ? normalCase_S_sqrt:normalCase_S_div; 
  assign sExpQuot_S_div_hi=io_b_sExp[8]; 
  assign sExpQuot_S_div_lo=~io_b_sExp[7:0]; 
  assign _sExpQuot_S_div_T_2={sExpQuot_S_div_hi,sExpQuot_S_div_lo}; 
  assign _GEN_13={{1{_sExpQuot_S_div_T_2[8]}},_sExpQuot_S_div_T_2}; 
  assign sExpQuot_S_div=$signed(io_a_sExp)+$signed(_GEN_13); 
  assign _sSatExpQuot_S_div_T=11'sh1c0<=$signed(sExpQuot_S_div); 
  assign sSatExpQuot_S_div_hi=_sSatExpQuot_S_div_T ? 4'h6:sExpQuot_S_div[9:6]; 
  assign sSatExpQuot_S_div_lo=sExpQuot_S_div[5:0]; 
  assign sSatExpQuot_S_div={sSatExpQuot_S_div_hi,sSatExpQuot_S_div_lo}; 
  assign evenSqrt_S=io_sqrtOp&~io_a_sExp[0]; 
  assign oddSqrt_S=io_sqrtOp&io_a_sExp[0]; 
  assign idle=cycleNum[0]; 
  assign inReady=idle|cycleNum[1]; 
  assign entering=inReady&io_inValid; 
  assign entering_normalCase=entering&normalCase_S; 
  assign skipCycle2=cycleNum[3]&sigX_Z[25]; 
  assign _T_1=~idle|entering; 
  assign _cycleNum_T_1=entering&~normalCase_S; 
  assign _cycleNum_T_2=_cycleNum_T_1 ? 2'h2:2'h0; 
  assign _cycleNum_T_4=io_a_sExp[0] ? 26'h1000000:26'h2000000; 
  assign _cycleNum_T_5=io_sqrtOp ? {1'b0,_cycleNum_T_4}:27'h4000000; 
  assign _cycleNum_T_6=entering_normalCase ? _cycleNum_T_5:27'h0; 
  assign _GEN_14={25'b0,_cycleNum_T_2}; 
  assign _cycleNum_T_7=_GEN_14|_cycleNum_T_6; 
  assign _cycleNum_T_10=~entering&~skipCycle2; 
  assign _cycleNum_T_12=_cycleNum_T_10 ? cycleNum[26:1]:26'h0; 
  assign _GEN_15={1'b0,_cycleNum_T_12}; 
  assign _cycleNum_T_13=_cycleNum_T_7|_GEN_15; 
  assign _cycleNum_T_14=skipCycle2 ? 2'h2:2'h0; 
  assign _GEN_16={25'b0,_cycleNum_T_14}; 
  assign _cycleNum_T_15=_cycleNum_T_13|_GEN_16; 
  assign _sExp_Z_T=io_a_sExp[9:1]; 
  assign _sExp_Z_T_1=$signed(_sExp_Z_T)+9'sh80; 
  assign _T_3=entering_normalCase&~io_sqrtOp; 
  assign _rem_T_1=inReady&~oddSqrt_S; 
  assign _rem_T_2={io_a_sig,1'h0}; 
  assign _rem_T_3=_rem_T_1 ? _rem_T_2:26'h0; 
  assign _rem_T_4=inReady&oddSqrt_S; 
  assign rem_hi=io_a_sig[23:22]-2'h1; 
  assign rem_lo={io_a_sig[21:0],3'h0}; 
  assign _rem_T_8={rem_hi,rem_lo}; 
  assign _rem_T_9=_rem_T_4 ? _rem_T_8:27'h0; 
  assign _GEN_17={1'b0,_rem_T_3}; 
  assign _rem_T_10=_GEN_17|_rem_T_9; 
  assign _rem_T_12={rem_Z,1'h0}; 
  assign _rem_T_13=inReady ? 27'h0:_rem_T_12; 
  assign rem=_rem_T_10|_rem_T_13; 
  assign bitMask=cycleNum[26:2]; 
  assign _trialTerm_T_1=inReady&~io_sqrtOp; 
  assign _trialTerm_T_2={io_b_sig,1'h0}; 
  assign _trialTerm_T_3=_trialTerm_T_1 ? _trialTerm_T_2:26'h0; 
  assign _trialTerm_T_4=inReady&evenSqrt_S; 
  assign _trialTerm_T_5=_trialTerm_T_4 ? 25'h1000000:25'h0; 
  assign _GEN_18={1'b0,_trialTerm_T_5}; 
  assign _trialTerm_T_6=_trialTerm_T_3|_GEN_18; 
  assign _trialTerm_T_8=_rem_T_4 ? 26'h2800000:26'h0; 
  assign _trialTerm_T_9=_trialTerm_T_6|_trialTerm_T_8; 
  assign _trialTerm_T_12=~inReady&~sqrtOp_Z; 
  assign _trialTerm_T_13={1'h1,fractB_Z}; 
  assign _trialTerm_T_14={_trialTerm_T_13,1'h0}; 
  assign _trialTerm_T_15=_trialTerm_T_12 ? _trialTerm_T_14:25'h0; 
  assign _GEN_19={1'b0,_trialTerm_T_15}; 
  assign _trialTerm_T_16=_trialTerm_T_9|_GEN_19; 
  assign _trialTerm_T_18=~inReady&sqrtOp_Z; 
  assign _trialTerm_T_19={sigX_Z,1'h0}; 
  assign _GEN_20={2'b0,bitMask}; 
  assign _trialTerm_T_20=_trialTerm_T_19|_GEN_20; 
  assign _trialTerm_T_21=_trialTerm_T_18 ? _trialTerm_T_20:27'h0; 
  assign _GEN_21={1'b0,_trialTerm_T_16}; 
  assign trialTerm=_GEN_21|_trialTerm_T_21; 
  assign _trialRem_T={1'b0,$signed(rem)}; 
  assign _trialRem_T_1={1'b0,$signed(trialTerm)}; 
  assign trialRem=$signed(_trialRem_T)-$signed(_trialRem_T_1); 
  assign newBit=28'sh0<=$signed(trialRem); 
  assign _T_5=idle|cycleNum[2]; 
  assign _T_7=entering_normalCase|~_T_5; 
  assign _rem_Z_T=$signed(_trialRem_T)-$signed(_trialRem_T_1); 
  assign _rem_Z_T_1=newBit ? _rem_Z_T:{1'b0,rem}; 
  assign _GEN_10=_T_7 ? _rem_Z_T_1:{2'b0,rem_Z}; 
  assign _T_9=~inReady&newBit; 
  assign _T_10=entering_normalCase|_T_9; 
  assign _notZeroRem_Z_T=$signed(trialRem)!=28'sh0; 
  assign _sigX_Z_T_2={newBit,25'h0}; 
  assign _sigX_Z_T_3=_trialTerm_T_1 ? _sigX_Z_T_2:26'h0; 
  assign _sigX_Z_T_4=inReady&io_sqrtOp; 
  assign _sigX_Z_T_5=_sigX_Z_T_4 ? 25'h1000000:25'h0; 
  assign _GEN_22={1'b0,_sigX_Z_T_5}; 
  assign _sigX_Z_T_6=_sigX_Z_T_3|_GEN_22; 
  assign _sigX_Z_T_8={newBit,23'h0}; 
  assign _sigX_Z_T_9=_rem_T_4 ? _sigX_Z_T_8:24'h0; 
  assign _GEN_23={2'b0,_sigX_Z_T_9}; 
  assign _sigX_Z_T_10=_sigX_Z_T_6|_GEN_23; 
  assign _GEN_24={1'b0,bitMask}; 
  assign _sigX_Z_T_12=sigX_Z|_GEN_24; 
  assign _sigX_Z_T_13=inReady ? 26'h0:_sigX_Z_T_12; 
  assign _sigX_Z_T_14=_sigX_Z_T_10|_sigX_Z_T_13; 
  assign _GEN_25={26'b0,notZeroRem_Z}; 
  assign io_inReady=idle|cycleNum[1]; 
  assign io_rawOutValid_div=cycleNum[1]&~sqrtOp_Z; 
  assign io_rawOutValid_sqrt=cycleNum[1]&sqrtOp_Z; 
  assign io_roundingModeOut=roundingMode_Z; 
  assign io_invalidExc=majorExc_Z&isNaN_Z; 
  assign io_infiniteExc=majorExc_Z&~isNaN_Z; 
  assign io_rawOut_isNaN=isNaN_Z; 
  assign io_rawOut_isInf=isInf_Z; 
  assign io_rawOut_isZero=isZero_Z; 
  assign io_rawOut_sign=sign_Z; 
  assign io_rawOut_sExp=sExp_Z; 
  assign io_rawOut_sig=_trialTerm_T_19|_GEN_25; 
  assign DivSqrtRawFN_small_cov_read_addr=DivSqrtRawFN_small_state; 
  assign DivSqrtRawFN_small_cov_read_data=DivSqrtRawFN_small_cov[DivSqrtRawFN_small_cov_read_addr]; 
  assign DivSqrtRawFN_small_cov_write_data=1'h1; 
  assign DivSqrtRawFN_small_cov_write_addr=DivSqrtRawFN_small_state; 
  assign DivSqrtRawFN_small_cov_write_mask=1'h1; 
  assign DivSqrtRawFN_small_cov_write_en=1'h1; 
  assign mux_cond_0=_T_10; 
  assign mux_cond_1=newBit; 
  assign mux_cond_2=skipCycle2; 
  assign mux_cond_3=_cycleNum_T_10; 
  assign sqrtOp_Z_shl=sqrtOp_Z; 
  assign sqrtOp_Z_pad={4'h0,sqrtOp_Z_shl}; 
  assign mux_cond_0_shl={mux_cond_0,1'h0}; 
  assign mux_cond_0_pad={3'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,2'h0}; 
  assign mux_cond_1_pad={2'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl={mux_cond_2,3'h0}; 
  assign mux_cond_2_pad={1'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,4'h0}; 
  assign mux_cond_3_pad=mux_cond_3_shl; 
  assign DivSqrtRawFN_small_xor1=sqrtOp_Z_pad^mux_cond_0_pad; 
  assign DivSqrtRawFN_small_xor6=mux_cond_2_pad^mux_cond_3_pad; 
  assign DivSqrtRawFN_small_xor2=mux_cond_1_pad^DivSqrtRawFN_small_xor6; 
  assign DivSqrtRawFN_small_xor0=DivSqrtRawFN_small_xor1^DivSqrtRawFN_small_xor2; 
  assign io_covSum=DivSqrtRawFN_small_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              cycleNum <=27'h0;
            end 
          else 
            if (reset)
               begin 
                 cycleNum <=27'h1;
               end 
             else 
               if (_T_1)
                  begin 
                    cycleNum <=_cycleNum_T_15;
                  end 
         if (metaReset)
            begin 
              sqrtOp_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 sqrtOp_Z <=io_sqrtOp;
               end 
         if (metaReset)
            begin 
              majorExc_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      majorExc_Z <=_majorExc_S_T_3;
                    end 
                  else 
                    begin 
                      majorExc_Z <=_majorExc_S_T_16;
                    end 
               end 
         if (metaReset)
            begin 
              isNaN_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      isNaN_Z <=_isNaN_S_T;
                    end 
                  else 
                    begin 
                      isNaN_Z <=_isNaN_S_T_2;
                    end 
               end 
         if (metaReset)
            begin 
              isInf_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      isInf_Z <=io_a_isInf;
                    end 
                  else 
                    begin 
                      isInf_Z <=_isInf_S_T;
                    end 
               end 
         if (metaReset)
            begin 
              isZero_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      isZero_Z <=io_a_isZero;
                    end 
                  else 
                    begin 
                      isZero_Z <=_isZero_S_T;
                    end 
               end 
         if (metaReset)
            begin 
              sign_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 sign_Z <=sign_S;
               end 
         if (metaReset)
            begin 
              sExp_Z <=10'h0;
            end 
          else 
            if (entering_normalCase)
               begin 
                 if (io_sqrtOp)
                    begin 
                      sExp_Z <=_sExp_Z_T_1;
                    end 
                  else 
                    begin 
                      sExp_Z <=sSatExpQuot_S_div;
                    end 
               end 
         if (metaReset)
            begin 
              fractB_Z <=23'h0;
            end 
          else 
            if (_T_3)
               begin 
                 fractB_Z <=io_b_sig[22:0];
               end 
         if (metaReset)
            begin 
              roundingMode_Z <=3'h0;
            end 
          else 
            if (entering_normalCase)
               begin 
                 roundingMode_Z <=io_roundingMode;
               end 
         if (metaReset)
            begin 
              rem_Z <=26'h0;
            end 
          else 
            begin 
              rem_Z <=_GEN_10[25:0];
            end 
         if (metaReset)
            begin 
              notZeroRem_Z <=1'h0;
            end 
          else 
            if (_T_10)
               begin 
                 notZeroRem_Z <=_notZeroRem_Z_T;
               end 
         if (metaReset)
            begin 
              sigX_Z <=26'h0;
            end 
          else 
            if (_T_10)
               begin 
                 sigX_Z <=_sigX_Z_T_14;
               end 
         DivSqrtRawFN_small_state <=DivSqrtRawFN_small_xor0;
         if (!(DivSqrtRawFN_small_cov_read_data))
            begin 
              DivSqrtRawFN_small_covSum <=DivSqrtRawFN_small_covSum+1'h1;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (DivSqrtRawFN_small_cov_write_en&DivSqrtRawFN_small_cov_write_mask)
            begin 
              DivSqrtRawFN_small_cov [DivSqrtRawFN_small_cov_write_addr]<=DivSqrtRawFN_small_cov_write_data;
            end 
       end
  
endmodule
 
module RoundAnyRawFNToRecFN_5 (
  input io_invalidExc,
  input io_infiniteExc,
  input io_in_isNaN,
  input io_in_isInf,
  input io_in_isZero,
  input io_in_sign,
  input [9:0] io_in_sExp,
  input [26:0] io_in_sig,
  input [2:0] io_roundingMode,
  input io_detectTininess,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundingMode_near_even ;  
   wire roundingMode_min ;  
   wire roundingMode_max ;  
   wire roundingMode_near_maxMag ;  
   wire roundingMode_odd ;  
   wire _roundMagUp_T ;  
   wire _roundMagUp_T_2 ;  
   wire roundMagUp ;  
   wire doShiftSigDown1 ;  
   wire roundMask_msb ;  
   wire [7:0] roundMask_lsbs ;  
   wire roundMask_msb_1 ;  
   wire [6:0] roundMask_lsbs_1 ;  
   wire roundMask_msb_2 ;  
   wire [5:0] roundMask_lsbs_2 ;  
   wire [64:0] roundMask_shift ;  
   wire [15:0] _roundMask_T_7 ;  
   wire [15:0] _roundMask_T_9 ;  
   wire [15:0] _roundMask_T_11 ;  
   wire [15:0] _roundMask_T_12 ;  
   wire [15:0] _GEN_0 ;  
   wire [15:0] _roundMask_T_17 ;  
   wire [15:0] _roundMask_T_19 ;  
   wire [15:0] _roundMask_T_21 ;  
   wire [15:0] _roundMask_T_22 ;  
   wire [15:0] _GEN_1 ;  
   wire [15:0] _roundMask_T_27 ;  
   wire [15:0] _roundMask_T_29 ;  
   wire [15:0] _roundMask_T_31 ;  
   wire [15:0] _roundMask_T_32 ;  
   wire [15:0] _GEN_2 ;  
   wire [15:0] _roundMask_T_37 ;  
   wire [15:0] _roundMask_T_39 ;  
   wire [15:0] _roundMask_T_41 ;  
   wire [15:0] roundMask_hi ;  
   wire roundMask_hi_1 ;  
   wire roundMask_lo ;  
   wire roundMask_hi_3 ;  
   wire roundMask_lo_1 ;  
   wire roundMask_hi_5 ;  
   wire roundMask_lo_3 ;  
   wire [21:0] _roundMask_T_47 ;  
   wire [21:0] _roundMask_T_49 ;  
   wire [21:0] roundMask_hi_6 ;  
   wire [24:0] _roundMask_T_50 ;  
   wire roundMask_hi_7 ;  
   wire roundMask_lo_6 ;  
   wire roundMask_lo_7 ;  
   wire [2:0] _roundMask_T_53 ;  
   wire [2:0] _roundMask_T_54 ;  
   wire [24:0] _roundMask_T_55 ;  
   wire [24:0] _roundMask_T_56 ;  
   wire [24:0] _GEN_3 ;  
   wire [24:0] roundMask_hi_9 ;  
   wire [26:0] roundMask ;  
   wire [25:0] shiftedRoundMask_lo ;  
   wire [26:0] shiftedRoundMask ;  
   wire [26:0] roundPosMask ;  
   wire [26:0] _roundPosBit_T ;  
   wire roundPosBit ;  
   wire [26:0] _anyRoundExtra_T ;  
   wire anyRoundExtra ;  
   wire anyRound ;  
   wire _roundIncr_T ;  
   wire _roundIncr_T_1 ;  
   wire _roundIncr_T_2 ;  
   wire roundIncr ;  
   wire [26:0] _roundedSig_T ;  
   wire [25:0] _roundedSig_T_2 ;  
   wire _roundedSig_T_3 ;  
   wire _roundedSig_T_5 ;  
   wire [25:0] _roundedSig_T_7 ;  
   wire [25:0] _roundedSig_T_9 ;  
   wire [26:0] _roundedSig_T_11 ;  
   wire _roundedSig_T_13 ;  
   wire [25:0] _roundedSig_T_15 ;  
   wire [25:0] _GEN_4 ;  
   wire [25:0] _roundedSig_T_16 ;  
   wire [25:0] roundedSig ;  
   wire [2:0] _sRoundedExp_T_1 ;  
   wire [9:0] _GEN_5 ;  
   wire [10:0] sRoundedExp ;  
   wire [8:0] common_expOut ;  
   wire [22:0] common_fractOut ;  
   wire [3:0] _common_overflow_T ;  
   wire common_overflow ;  
   wire common_totalUnderflow ;  
   wire unboundedRange_roundPosBit ;  
   wire _unboundedRange_anyRound_T_1 ;  
   wire _unboundedRange_anyRound_T_3 ;  
   wire unboundedRange_anyRound ;  
   wire _unboundedRange_roundIncr_T_1 ;  
   wire _unboundedRange_roundIncr_T_2 ;  
   wire unboundedRange_roundIncr ;  
   wire roundCarry ;  
   wire [1:0] _common_underflow_T ;  
   wire _common_underflow_T_1 ;  
   wire _common_underflow_T_2 ;  
   wire _common_underflow_T_5 ;  
   wire _common_underflow_T_6 ;  
   wire _common_underflow_T_10 ;  
   wire _common_underflow_T_12 ;  
   wire _common_underflow_T_13 ;  
   wire _common_underflow_T_14 ;  
   wire _common_underflow_T_15 ;  
   wire _common_underflow_T_17 ;  
   wire common_underflow ;  
   wire common_inexact ;  
   wire isNaNOut ;  
   wire notNaN_isSpecialInfOut ;  
   wire _commonCase_T_2 ;  
   wire commonCase ;  
   wire overflow ;  
   wire underflow ;  
   wire _inexact_T ;  
   wire inexact ;  
   wire overflow_roundMagUp ;  
   wire _pegMinNonzeroMagOut_T ;  
   wire _pegMinNonzeroMagOut_T_1 ;  
   wire pegMinNonzeroMagOut ;  
   wire pegMaxFiniteMagOut ;  
   wire _notNaN_isInfOut_T ;  
   wire notNaN_isInfOut ;  
   wire signOut ;  
   wire _expOut_T ;  
   wire [8:0] _expOut_T_1 ;  
   wire [8:0] _expOut_T_3 ;  
   wire [8:0] _expOut_T_5 ;  
   wire [8:0] _expOut_T_7 ;  
   wire [8:0] _expOut_T_8 ;  
   wire [8:0] _expOut_T_10 ;  
   wire [8:0] _expOut_T_11 ;  
   wire [8:0] _expOut_T_13 ;  
   wire [8:0] _expOut_T_14 ;  
   wire [8:0] _expOut_T_15 ;  
   wire [8:0] _expOut_T_16 ;  
   wire [8:0] _expOut_T_17 ;  
   wire [8:0] _expOut_T_18 ;  
   wire [8:0] _expOut_T_19 ;  
   wire [8:0] _expOut_T_20 ;  
   wire [8:0] expOut ;  
   wire _fractOut_T ;  
   wire _fractOut_T_1 ;  
   wire [22:0] _fractOut_T_2 ;  
   wire [22:0] _fractOut_T_3 ;  
   wire [22:0] _fractOut_T_5 ;  
   wire [22:0] fractOut ;  
   wire [9:0] io_out_hi ;  
   wire [1:0] io_exceptionFlags_lo ;  
   wire [2:0] io_exceptionFlags_hi ;  
   wire [29:0] RoundAnyRawFNToRecFN_5_covSum ;  
  assign roundingMode_near_even=io_roundingMode==3'h0; 
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign roundingMode_max=io_roundingMode==3'h3; 
  assign roundingMode_near_maxMag=io_roundingMode==3'h4; 
  assign roundingMode_odd=io_roundingMode==3'h6; 
  assign _roundMagUp_T=roundingMode_min&io_in_sign; 
  assign _roundMagUp_T_2=roundingMode_max&~io_in_sign; 
  assign roundMagUp=_roundMagUp_T|_roundMagUp_T_2; 
  assign doShiftSigDown1=io_in_sig[26]; 
  assign roundMask_msb=~io_in_sExp[8]; 
  assign roundMask_lsbs=~io_in_sExp[7:0]; 
  assign roundMask_msb_1=roundMask_lsbs[7]; 
  assign roundMask_lsbs_1=roundMask_lsbs[6:0]; 
  assign roundMask_msb_2=roundMask_lsbs_1[6]; 
  assign roundMask_lsbs_2=roundMask_lsbs_1[5:0]; 
  assign roundMask_shift=-65'sh10000000000000000>>>roundMask_lsbs_2; 
  assign _roundMask_T_7={8'b0,roundMask_shift[57:50]}; 
  assign _roundMask_T_9={roundMask_shift[49:42],8'h0}; 
  assign _roundMask_T_11=_roundMask_T_9&16'hff00; 
  assign _roundMask_T_12=_roundMask_T_7|_roundMask_T_11; 
  assign _GEN_0={4'b0,_roundMask_T_12[15:4]}; 
  assign _roundMask_T_17=_GEN_0&16'hf0f; 
  assign _roundMask_T_19={_roundMask_T_12[11:0],4'h0}; 
  assign _roundMask_T_21=_roundMask_T_19&16'hf0f0; 
  assign _roundMask_T_22=_roundMask_T_17|_roundMask_T_21; 
  assign _GEN_1={2'b0,_roundMask_T_22[15:2]}; 
  assign _roundMask_T_27=_GEN_1&16'h3333; 
  assign _roundMask_T_29={_roundMask_T_22[13:0],2'h0}; 
  assign _roundMask_T_31=_roundMask_T_29&16'hcccc; 
  assign _roundMask_T_32=_roundMask_T_27|_roundMask_T_31; 
  assign _GEN_2={1'b0,_roundMask_T_32[15:1]}; 
  assign _roundMask_T_37=_GEN_2&16'h5555; 
  assign _roundMask_T_39={_roundMask_T_32[14:0],1'h0}; 
  assign _roundMask_T_41=_roundMask_T_39&16'haaaa; 
  assign roundMask_hi=_roundMask_T_37|_roundMask_T_41; 
  assign roundMask_hi_1=roundMask_shift[58]; 
  assign roundMask_lo=roundMask_shift[59]; 
  assign roundMask_hi_3=roundMask_shift[60]; 
  assign roundMask_lo_1=roundMask_shift[61]; 
  assign roundMask_hi_5=roundMask_shift[62]; 
  assign roundMask_lo_3=roundMask_shift[63]; 
  assign _roundMask_T_47={roundMask_hi,roundMask_hi_1,roundMask_lo,roundMask_hi_3,roundMask_lo_1,roundMask_hi_5,roundMask_lo_3}; 
  assign _roundMask_T_49=roundMask_msb_2 ? 22'h0:~_roundMask_T_47; 
  assign roundMask_hi_6=~_roundMask_T_49; 
  assign _roundMask_T_50={roundMask_hi_6,3'h7}; 
  assign roundMask_hi_7=roundMask_shift[0]; 
  assign roundMask_lo_6=roundMask_shift[1]; 
  assign roundMask_lo_7=roundMask_shift[2]; 
  assign _roundMask_T_53={roundMask_hi_7,roundMask_lo_6,roundMask_lo_7}; 
  assign _roundMask_T_54=roundMask_msb_2 ? _roundMask_T_53:3'h0; 
  assign _roundMask_T_55=roundMask_msb_1 ? _roundMask_T_50:{22'b0,_roundMask_T_54}; 
  assign _roundMask_T_56=roundMask_msb ? _roundMask_T_55:25'h0; 
  assign _GEN_3={24'b0,doShiftSigDown1}; 
  assign roundMask_hi_9=_roundMask_T_56|_GEN_3; 
  assign roundMask={roundMask_hi_9,2'h3}; 
  assign shiftedRoundMask_lo=roundMask[26:1]; 
  assign shiftedRoundMask={1'h0,shiftedRoundMask_lo}; 
  assign roundPosMask=~shiftedRoundMask&roundMask; 
  assign _roundPosBit_T=io_in_sig&roundPosMask; 
  assign roundPosBit=|_roundPosBit_T; 
  assign _anyRoundExtra_T=io_in_sig&shiftedRoundMask; 
  assign anyRoundExtra=|_anyRoundExtra_T; 
  assign anyRound=roundPosBit|anyRoundExtra; 
  assign _roundIncr_T=roundingMode_near_even|roundingMode_near_maxMag; 
  assign _roundIncr_T_1=_roundIncr_T&roundPosBit; 
  assign _roundIncr_T_2=roundMagUp&anyRound; 
  assign roundIncr=_roundIncr_T_1|_roundIncr_T_2; 
  assign _roundedSig_T=io_in_sig|roundMask; 
  assign _roundedSig_T_2=_roundedSig_T[26:2]+25'h1; 
  assign _roundedSig_T_3=roundingMode_near_even&roundPosBit; 
  assign _roundedSig_T_5=_roundedSig_T_3&~anyRoundExtra; 
  assign _roundedSig_T_7=_roundedSig_T_5 ? shiftedRoundMask_lo:26'h0; 
  assign _roundedSig_T_9=_roundedSig_T_2&~_roundedSig_T_7; 
  assign _roundedSig_T_11=io_in_sig&~roundMask; 
  assign _roundedSig_T_13=roundingMode_odd&anyRound; 
  assign _roundedSig_T_15=_roundedSig_T_13 ? roundPosMask[26:1]:26'h0; 
  assign _GEN_4={1'b0,_roundedSig_T_11[26:2]}; 
  assign _roundedSig_T_16=_GEN_4|_roundedSig_T_15; 
  assign roundedSig=roundIncr ? _roundedSig_T_9:_roundedSig_T_16; 
  assign _sRoundedExp_T_1={1'b0,$signed(roundedSig[25:24])}; 
  assign _GEN_5={{7{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; 
  assign sRoundedExp=$signed(io_in_sExp)+$signed(_GEN_5); 
  assign common_expOut=sRoundedExp[8:0]; 
  assign common_fractOut=doShiftSigDown1 ? roundedSig[23:1]:roundedSig[22:0]; 
  assign _common_overflow_T=sRoundedExp[10:7]; 
  assign common_overflow=$signed(_common_overflow_T)>=4'sh3; 
  assign common_totalUnderflow=$signed(sRoundedExp)<11'sh6b; 
  assign unboundedRange_roundPosBit=doShiftSigDown1 ? io_in_sig[2]:io_in_sig[1]; 
  assign _unboundedRange_anyRound_T_1=doShiftSigDown1&io_in_sig[2]; 
  assign _unboundedRange_anyRound_T_3=|io_in_sig[1:0]; 
  assign unboundedRange_anyRound=_unboundedRange_anyRound_T_1|_unboundedRange_anyRound_T_3; 
  assign _unboundedRange_roundIncr_T_1=_roundIncr_T&unboundedRange_roundPosBit; 
  assign _unboundedRange_roundIncr_T_2=roundMagUp&unboundedRange_anyRound; 
  assign unboundedRange_roundIncr=_unboundedRange_roundIncr_T_1|_unboundedRange_roundIncr_T_2; 
  assign roundCarry=doShiftSigDown1 ? roundedSig[25]:roundedSig[24]; 
  assign _common_underflow_T=io_in_sExp[9:8]; 
  assign _common_underflow_T_1=$signed(_common_underflow_T)<=2'sh0; 
  assign _common_underflow_T_2=anyRound&_common_underflow_T_1; 
  assign _common_underflow_T_5=doShiftSigDown1 ? roundMask[3]:roundMask[2]; 
  assign _common_underflow_T_6=_common_underflow_T_2&_common_underflow_T_5; 
  assign _common_underflow_T_10=doShiftSigDown1 ? roundMask[4]:roundMask[3]; 
  assign _common_underflow_T_12=io_detectTininess&~_common_underflow_T_10; 
  assign _common_underflow_T_13=_common_underflow_T_12&roundCarry; 
  assign _common_underflow_T_14=_common_underflow_T_13&roundPosBit; 
  assign _common_underflow_T_15=_common_underflow_T_14&unboundedRange_roundIncr; 
  assign _common_underflow_T_17=_common_underflow_T_6&~_common_underflow_T_15; 
  assign common_underflow=common_totalUnderflow|_common_underflow_T_17; 
  assign common_inexact=common_totalUnderflow|anyRound; 
  assign isNaNOut=io_invalidExc|io_in_isNaN; 
  assign notNaN_isSpecialInfOut=io_infiniteExc|io_in_isInf; 
  assign _commonCase_T_2=~isNaNOut&~notNaN_isSpecialInfOut; 
  assign commonCase=_commonCase_T_2&~io_in_isZero; 
  assign overflow=commonCase&common_overflow; 
  assign underflow=commonCase&common_underflow; 
  assign _inexact_T=commonCase&common_inexact; 
  assign inexact=overflow|_inexact_T; 
  assign overflow_roundMagUp=_roundIncr_T|roundMagUp; 
  assign _pegMinNonzeroMagOut_T=commonCase&common_totalUnderflow; 
  assign _pegMinNonzeroMagOut_T_1=roundMagUp|roundingMode_odd; 
  assign pegMinNonzeroMagOut=_pegMinNonzeroMagOut_T&_pegMinNonzeroMagOut_T_1; 
  assign pegMaxFiniteMagOut=overflow&~overflow_roundMagUp; 
  assign _notNaN_isInfOut_T=overflow&overflow_roundMagUp; 
  assign notNaN_isInfOut=notNaN_isSpecialInfOut|_notNaN_isInfOut_T; 
  assign signOut=isNaNOut ? 1'h0:io_in_sign; 
  assign _expOut_T=io_in_isZero|common_totalUnderflow; 
  assign _expOut_T_1=_expOut_T ? 9'h1c0:9'h0; 
  assign _expOut_T_3=common_expOut&~_expOut_T_1; 
  assign _expOut_T_5=pegMinNonzeroMagOut ? 9'h194:9'h0; 
  assign _expOut_T_7=_expOut_T_3&~_expOut_T_5; 
  assign _expOut_T_8=pegMaxFiniteMagOut ? 9'h80:9'h0; 
  assign _expOut_T_10=_expOut_T_7&~_expOut_T_8; 
  assign _expOut_T_11=notNaN_isInfOut ? 9'h40:9'h0; 
  assign _expOut_T_13=_expOut_T_10&~_expOut_T_11; 
  assign _expOut_T_14=pegMinNonzeroMagOut ? 9'h6b:9'h0; 
  assign _expOut_T_15=_expOut_T_13|_expOut_T_14; 
  assign _expOut_T_16=pegMaxFiniteMagOut ? 9'h17f:9'h0; 
  assign _expOut_T_17=_expOut_T_15|_expOut_T_16; 
  assign _expOut_T_18=notNaN_isInfOut ? 9'h180:9'h0; 
  assign _expOut_T_19=_expOut_T_17|_expOut_T_18; 
  assign _expOut_T_20=isNaNOut ? 9'h1c0:9'h0; 
  assign expOut=_expOut_T_19|_expOut_T_20; 
  assign _fractOut_T=isNaNOut|io_in_isZero; 
  assign _fractOut_T_1=_fractOut_T|common_totalUnderflow; 
  assign _fractOut_T_2=isNaNOut ? 23'h400000:23'h0; 
  assign _fractOut_T_3=_fractOut_T_1 ? _fractOut_T_2:common_fractOut; 
  assign _fractOut_T_5=pegMaxFiniteMagOut ? 23'h7fffff:23'h0; 
  assign fractOut=_fractOut_T_3|_fractOut_T_5; 
  assign io_out_hi={signOut,expOut}; 
  assign io_exceptionFlags_lo={underflow,inexact}; 
  assign io_exceptionFlags_hi={io_invalidExc,io_infiniteExc,overflow}; 
  assign io_out={io_out_hi,fractOut}; 
  assign io_exceptionFlags={io_exceptionFlags_hi,io_exceptionFlags_lo}; 
  assign RoundAnyRawFNToRecFN_5_covSum=30'h0; 
  assign io_covSum=RoundAnyRawFNToRecFN_5_covSum; 
  assign metaAssert=1'h0; 
endmodule
 
module DivSqrtRawFN_small_1 (
  input clock,
  input reset,
  output io_inReady,
  input io_inValid,
  input io_sqrtOp,
  input io_a_isNaN,
  input io_a_isInf,
  input io_a_isZero,
  input io_a_sign,
  input [12:0] io_a_sExp,
  input [53:0] io_a_sig,
  input io_b_isNaN,
  input io_b_isInf,
  input io_b_isZero,
  input io_b_sign,
  input [12:0] io_b_sExp,
  input [53:0] io_b_sig,
  input [2:0] io_roundingMode,
  output io_rawOutValid_div,
  output io_rawOutValid_sqrt,
  output [2:0] io_roundingModeOut,
  output io_invalidExc,
  output io_infiniteExc,
  output io_rawOut_isNaN,
  output io_rawOut_isInf,
  output io_rawOut_isZero,
  output io_rawOut_sign,
  output [12:0] io_rawOut_sExp,
  output [55:0] io_rawOut_sig,
  output [29:0] io_covSum,
  output metaAssert,
  input metaReset) ; 
   reg [55:0] cycleNum ;  
   reg [63:0] _RAND_0 ;  
   reg sqrtOp_Z ;  
   reg [31:0] _RAND_1 ;  
   reg majorExc_Z ;  
   reg [31:0] _RAND_2 ;  
   reg isNaN_Z ;  
   reg [31:0] _RAND_3 ;  
   reg isInf_Z ;  
   reg [31:0] _RAND_4 ;  
   reg isZero_Z ;  
   reg [31:0] _RAND_5 ;  
   reg sign_Z ;  
   reg [31:0] _RAND_6 ;  
   reg [12:0] sExp_Z ;  
   reg [31:0] _RAND_7 ;  
   reg [51:0] fractB_Z ;  
   reg [63:0] _RAND_8 ;  
   reg [2:0] roundingMode_Z ;  
   reg [31:0] _RAND_9 ;  
   reg [54:0] rem_Z ;  
   reg [63:0] _RAND_10 ;  
   reg notZeroRem_Z ;  
   reg [31:0] _RAND_11 ;  
   reg [54:0] sigX_Z ;  
   reg [63:0] _RAND_12 ;  
   wire _notSigNaNIn_invalidExc_S_div_T ;  
   wire _notSigNaNIn_invalidExc_S_div_T_1 ;  
   wire notSigNaNIn_invalidExc_S_div ;  
   wire _notSigNaNIn_invalidExc_S_sqrt_T_2 ;  
   wire notSigNaNIn_invalidExc_S_sqrt ;  
   wire _majorExc_S_T_2 ;  
   wire _majorExc_S_T_3 ;  
   wire _majorExc_S_T_9 ;  
   wire _majorExc_S_T_10 ;  
   wire _majorExc_S_T_11 ;  
   wire _majorExc_S_T_14 ;  
   wire _majorExc_S_T_15 ;  
   wire _majorExc_S_T_16 ;  
   wire _isNaN_S_T ;  
   wire _isNaN_S_T_1 ;  
   wire _isNaN_S_T_2 ;  
   wire _isInf_S_T ;  
   wire _isZero_S_T ;  
   wire _sign_S_T_1 ;  
   wire sign_S ;  
   wire _specialCaseA_S_T ;  
   wire specialCaseA_S ;  
   wire _specialCaseB_S_T ;  
   wire specialCaseB_S ;  
   wire normalCase_S_div ;  
   wire normalCase_S_sqrt ;  
   wire normalCase_S ;  
   wire sExpQuot_S_div_hi ;  
   wire [10:0] sExpQuot_S_div_lo ;  
   wire [11:0] _sExpQuot_S_div_T_2 ;  
   wire [12:0] _GEN_13 ;  
   wire [13:0] sExpQuot_S_div ;  
   wire _sSatExpQuot_S_div_T ;  
   wire [3:0] sSatExpQuot_S_div_hi ;  
   wire [8:0] sSatExpQuot_S_div_lo ;  
   wire [12:0] sSatExpQuot_S_div ;  
   wire evenSqrt_S ;  
   wire oddSqrt_S ;  
   wire idle ;  
   wire inReady ;  
   wire entering ;  
   wire entering_normalCase ;  
   wire skipCycle2 ;  
   wire _T_1 ;  
   wire _cycleNum_T_1 ;  
   wire [1:0] _cycleNum_T_2 ;  
   wire [54:0] _cycleNum_T_4 ;  
   wire [55:0] _cycleNum_T_5 ;  
   wire [55:0] _cycleNum_T_6 ;  
   wire [55:0] _GEN_14 ;  
   wire [55:0] _cycleNum_T_7 ;  
   wire _cycleNum_T_10 ;  
   wire [54:0] _cycleNum_T_12 ;  
   wire [55:0] _GEN_15 ;  
   wire [55:0] _cycleNum_T_13 ;  
   wire [1:0] _cycleNum_T_14 ;  
   wire [55:0] _GEN_16 ;  
   wire [55:0] _cycleNum_T_15 ;  
   wire [11:0] _sExp_Z_T ;  
   wire [12:0] _sExp_Z_T_1 ;  
   wire _T_3 ;  
   wire _rem_T_1 ;  
   wire [54:0] _rem_T_2 ;  
   wire [54:0] _rem_T_3 ;  
   wire _rem_T_4 ;  
   wire [1:0] rem_hi ;  
   wire [53:0] rem_lo ;  
   wire [55:0] _rem_T_8 ;  
   wire [55:0] _rem_T_9 ;  
   wire [55:0] _GEN_17 ;  
   wire [55:0] _rem_T_10 ;  
   wire [55:0] _rem_T_12 ;  
   wire [55:0] _rem_T_13 ;  
   wire [55:0] rem ;  
   wire [53:0] bitMask ;  
   wire _trialTerm_T_1 ;  
   wire [54:0] _trialTerm_T_2 ;  
   wire [54:0] _trialTerm_T_3 ;  
   wire _trialTerm_T_4 ;  
   wire [53:0] _trialTerm_T_5 ;  
   wire [54:0] _GEN_18 ;  
   wire [54:0] _trialTerm_T_6 ;  
   wire [54:0] _trialTerm_T_8 ;  
   wire [54:0] _trialTerm_T_9 ;  
   wire _trialTerm_T_12 ;  
   wire [52:0] _trialTerm_T_13 ;  
   wire [53:0] _trialTerm_T_14 ;  
   wire [53:0] _trialTerm_T_15 ;  
   wire [54:0] _GEN_19 ;  
   wire [54:0] _trialTerm_T_16 ;  
   wire _trialTerm_T_18 ;  
   wire [55:0] _trialTerm_T_19 ;  
   wire [55:0] _GEN_20 ;  
   wire [55:0] _trialTerm_T_20 ;  
   wire [55:0] _trialTerm_T_21 ;  
   wire [55:0] _GEN_21 ;  
   wire [55:0] trialTerm ;  
   wire [56:0] _trialRem_T ;  
   wire [56:0] _trialRem_T_1 ;  
   wire [56:0] trialRem ;  
   wire newBit ;  
   wire _T_5 ;  
   wire _T_7 ;  
   wire [56:0] _rem_Z_T ;  
   wire [56:0] _rem_Z_T_1 ;  
   wire [56:0] _GEN_10 ;  
   wire _T_9 ;  
   wire _T_10 ;  
   wire _notZeroRem_Z_T ;  
   wire [54:0] _sigX_Z_T_2 ;  
   wire [54:0] _sigX_Z_T_3 ;  
   wire _sigX_Z_T_4 ;  
   wire [53:0] _sigX_Z_T_5 ;  
   wire [54:0] _GEN_22 ;  
   wire [54:0] _sigX_Z_T_6 ;  
   wire [52:0] _sigX_Z_T_8 ;  
   wire [52:0] _sigX_Z_T_9 ;  
   wire [54:0] _GEN_23 ;  
   wire [54:0] _sigX_Z_T_10 ;  
   wire [54:0] _GEN_24 ;  
   wire [54:0] _sigX_Z_T_12 ;  
   wire [54:0] _sigX_Z_T_13 ;  
   wire [54:0] _sigX_Z_T_14 ;  
   wire [55:0] _GEN_25 ;  
   reg [4:0] DivSqrtRawFN_small_1_state ;  
   reg [31:0] _RAND_13 ;  
   reg DivSqrtRawFN_small_1_cov[0:31] ;  
   reg [31:0] _RAND_14 ;  
   wire DivSqrtRawFN_small_1_cov_read_data ;  
   wire [4:0] DivSqrtRawFN_small_1_cov_read_addr ;  
   wire DivSqrtRawFN_small_1_cov_write_data ;  
   wire [4:0] DivSqrtRawFN_small_1_cov_write_addr ;  
   wire DivSqrtRawFN_small_1_cov_write_mask ;  
   wire DivSqrtRawFN_small_1_cov_write_en ;  
   reg [29:0] DivSqrtRawFN_small_1_covSum ;  
   reg [31:0] _RAND_15 ;  
   wire mux_cond_0 ;  
   wire mux_cond_1 ;  
   wire mux_cond_2 ;  
   wire mux_cond_3 ;  
   wire sqrtOp_Z_shl ;  
   wire [4:0] sqrtOp_Z_pad ;  
   wire [1:0] mux_cond_0_shl ;  
   wire [4:0] mux_cond_0_pad ;  
   wire [2:0] mux_cond_1_shl ;  
   wire [4:0] mux_cond_1_pad ;  
   wire [3:0] mux_cond_2_shl ;  
   wire [4:0] mux_cond_2_pad ;  
   wire [4:0] mux_cond_3_shl ;  
   wire [4:0] mux_cond_3_pad ;  
   wire [4:0] DivSqrtRawFN_small_1_xor1 ;  
   wire [4:0] DivSqrtRawFN_small_1_xor6 ;  
   wire [4:0] DivSqrtRawFN_small_1_xor2 ;  
   wire [4:0] DivSqrtRawFN_small_1_xor0 ;  
  assign _notSigNaNIn_invalidExc_S_div_T=io_a_isZero&io_b_isZero; 
  assign _notSigNaNIn_invalidExc_S_div_T_1=io_a_isInf&io_b_isInf; 
  assign notSigNaNIn_invalidExc_S_div=_notSigNaNIn_invalidExc_S_div_T|_notSigNaNIn_invalidExc_S_div_T_1; 
  assign _notSigNaNIn_invalidExc_S_sqrt_T_2=~io_a_isNaN&~io_a_isZero; 
  assign notSigNaNIn_invalidExc_S_sqrt=_notSigNaNIn_invalidExc_S_sqrt_T_2&io_a_sign; 
  assign _majorExc_S_T_2=io_a_isNaN&~io_a_sig[51]; 
  assign _majorExc_S_T_3=_majorExc_S_T_2|notSigNaNIn_invalidExc_S_sqrt; 
  assign _majorExc_S_T_9=io_b_isNaN&~io_b_sig[51]; 
  assign _majorExc_S_T_10=_majorExc_S_T_2|_majorExc_S_T_9; 
  assign _majorExc_S_T_11=_majorExc_S_T_10|notSigNaNIn_invalidExc_S_div; 
  assign _majorExc_S_T_14=~io_a_isNaN&~io_a_isInf; 
  assign _majorExc_S_T_15=_majorExc_S_T_14&io_b_isZero; 
  assign _majorExc_S_T_16=_majorExc_S_T_11|_majorExc_S_T_15; 
  assign _isNaN_S_T=io_a_isNaN|notSigNaNIn_invalidExc_S_sqrt; 
  assign _isNaN_S_T_1=io_a_isNaN|io_b_isNaN; 
  assign _isNaN_S_T_2=_isNaN_S_T_1|notSigNaNIn_invalidExc_S_div; 
  assign _isInf_S_T=io_a_isInf|io_b_isZero; 
  assign _isZero_S_T=io_a_isZero|io_b_isInf; 
  assign _sign_S_T_1=~io_sqrtOp&io_b_sign; 
  assign sign_S=io_a_sign^_sign_S_T_1; 
  assign _specialCaseA_S_T=io_a_isNaN|io_a_isInf; 
  assign specialCaseA_S=_specialCaseA_S_T|io_a_isZero; 
  assign _specialCaseB_S_T=io_b_isNaN|io_b_isInf; 
  assign specialCaseB_S=_specialCaseB_S_T|io_b_isZero; 
  assign normalCase_S_div=~specialCaseA_S&~specialCaseB_S; 
  assign normalCase_S_sqrt=~specialCaseA_S&~io_a_sign; 
  assign normalCase_S=io_sqrtOp ? normalCase_S_sqrt:normalCase_S_div; 
  assign sExpQuot_S_div_hi=io_b_sExp[11]; 
  assign sExpQuot_S_div_lo=~io_b_sExp[10:0]; 
  assign _sExpQuot_S_div_T_2={sExpQuot_S_div_hi,sExpQuot_S_div_lo}; 
  assign _GEN_13={{1{_sExpQuot_S_div_T_2[11]}},_sExpQuot_S_div_T_2}; 
  assign sExpQuot_S_div=$signed(io_a_sExp)+$signed(_GEN_13); 
  assign _sSatExpQuot_S_div_T=14'she00<=$signed(sExpQuot_S_div); 
  assign sSatExpQuot_S_div_hi=_sSatExpQuot_S_div_T ? 4'h6:sExpQuot_S_div[12:9]; 
  assign sSatExpQuot_S_div_lo=sExpQuot_S_div[8:0]; 
  assign sSatExpQuot_S_div={sSatExpQuot_S_div_hi,sSatExpQuot_S_div_lo}; 
  assign evenSqrt_S=io_sqrtOp&~io_a_sExp[0]; 
  assign oddSqrt_S=io_sqrtOp&io_a_sExp[0]; 
  assign idle=cycleNum[0]; 
  assign inReady=idle|cycleNum[1]; 
  assign entering=inReady&io_inValid; 
  assign entering_normalCase=entering&normalCase_S; 
  assign skipCycle2=cycleNum[3]&sigX_Z[54]; 
  assign _T_1=~idle|entering; 
  assign _cycleNum_T_1=entering&~normalCase_S; 
  assign _cycleNum_T_2=_cycleNum_T_1 ? 2'h2:2'h0; 
  assign _cycleNum_T_4=io_a_sExp[0] ? 55'h20000000000000:55'h40000000000000; 
  assign _cycleNum_T_5=io_sqrtOp ? {1'b0,_cycleNum_T_4}:56'h80000000000000; 
  assign _cycleNum_T_6=entering_normalCase ? _cycleNum_T_5:56'h0; 
  assign _GEN_14={54'b0,_cycleNum_T_2}; 
  assign _cycleNum_T_7=_GEN_14|_cycleNum_T_6; 
  assign _cycleNum_T_10=~entering&~skipCycle2; 
  assign _cycleNum_T_12=_cycleNum_T_10 ? cycleNum[55:1]:55'h0; 
  assign _GEN_15={1'b0,_cycleNum_T_12}; 
  assign _cycleNum_T_13=_cycleNum_T_7|_GEN_15; 
  assign _cycleNum_T_14=skipCycle2 ? 2'h2:2'h0; 
  assign _GEN_16={54'b0,_cycleNum_T_14}; 
  assign _cycleNum_T_15=_cycleNum_T_13|_GEN_16; 
  assign _sExp_Z_T=io_a_sExp[12:1]; 
  assign _sExp_Z_T_1=$signed(_sExp_Z_T)+12'sh400; 
  assign _T_3=entering_normalCase&~io_sqrtOp; 
  assign _rem_T_1=inReady&~oddSqrt_S; 
  assign _rem_T_2={io_a_sig,1'h0}; 
  assign _rem_T_3=_rem_T_1 ? _rem_T_2:55'h0; 
  assign _rem_T_4=inReady&oddSqrt_S; 
  assign rem_hi=io_a_sig[52:51]-2'h1; 
  assign rem_lo={io_a_sig[50:0],3'h0}; 
  assign _rem_T_8={rem_hi,rem_lo}; 
  assign _rem_T_9=_rem_T_4 ? _rem_T_8:56'h0; 
  assign _GEN_17={1'b0,_rem_T_3}; 
  assign _rem_T_10=_GEN_17|_rem_T_9; 
  assign _rem_T_12={rem_Z,1'h0}; 
  assign _rem_T_13=inReady ? 56'h0:_rem_T_12; 
  assign rem=_rem_T_10|_rem_T_13; 
  assign bitMask=cycleNum[55:2]; 
  assign _trialTerm_T_1=inReady&~io_sqrtOp; 
  assign _trialTerm_T_2={io_b_sig,1'h0}; 
  assign _trialTerm_T_3=_trialTerm_T_1 ? _trialTerm_T_2:55'h0; 
  assign _trialTerm_T_4=inReady&evenSqrt_S; 
  assign _trialTerm_T_5=_trialTerm_T_4 ? 54'h20000000000000:54'h0; 
  assign _GEN_18={1'b0,_trialTerm_T_5}; 
  assign _trialTerm_T_6=_trialTerm_T_3|_GEN_18; 
  assign _trialTerm_T_8=_rem_T_4 ? 55'h50000000000000:55'h0; 
  assign _trialTerm_T_9=_trialTerm_T_6|_trialTerm_T_8; 
  assign _trialTerm_T_12=~inReady&~sqrtOp_Z; 
  assign _trialTerm_T_13={1'h1,fractB_Z}; 
  assign _trialTerm_T_14={_trialTerm_T_13,1'h0}; 
  assign _trialTerm_T_15=_trialTerm_T_12 ? _trialTerm_T_14:54'h0; 
  assign _GEN_19={1'b0,_trialTerm_T_15}; 
  assign _trialTerm_T_16=_trialTerm_T_9|_GEN_19; 
  assign _trialTerm_T_18=~inReady&sqrtOp_Z; 
  assign _trialTerm_T_19={sigX_Z,1'h0}; 
  assign _GEN_20={2'b0,bitMask}; 
  assign _trialTerm_T_20=_trialTerm_T_19|_GEN_20; 
  assign _trialTerm_T_21=_trialTerm_T_18 ? _trialTerm_T_20:56'h0; 
  assign _GEN_21={1'b0,_trialTerm_T_16}; 
  assign trialTerm=_GEN_21|_trialTerm_T_21; 
  assign _trialRem_T={1'b0,$signed(rem)}; 
  assign _trialRem_T_1={1'b0,$signed(trialTerm)}; 
  assign trialRem=$signed(_trialRem_T)-$signed(_trialRem_T_1); 
  assign newBit=57'sh0<=$signed(trialRem); 
  assign _T_5=idle|cycleNum[2]; 
  assign _T_7=entering_normalCase|~_T_5; 
  assign _rem_Z_T=$signed(_trialRem_T)-$signed(_trialRem_T_1); 
  assign _rem_Z_T_1=newBit ? _rem_Z_T:{1'b0,rem}; 
  assign _GEN_10=_T_7 ? _rem_Z_T_1:{2'b0,rem_Z}; 
  assign _T_9=~inReady&newBit; 
  assign _T_10=entering_normalCase|_T_9; 
  assign _notZeroRem_Z_T=$signed(trialRem)!=57'sh0; 
  assign _sigX_Z_T_2={newBit,54'h0}; 
  assign _sigX_Z_T_3=_trialTerm_T_1 ? _sigX_Z_T_2:55'h0; 
  assign _sigX_Z_T_4=inReady&io_sqrtOp; 
  assign _sigX_Z_T_5=_sigX_Z_T_4 ? 54'h20000000000000:54'h0; 
  assign _GEN_22={1'b0,_sigX_Z_T_5}; 
  assign _sigX_Z_T_6=_sigX_Z_T_3|_GEN_22; 
  assign _sigX_Z_T_8={newBit,52'h0}; 
  assign _sigX_Z_T_9=_rem_T_4 ? _sigX_Z_T_8:53'h0; 
  assign _GEN_23={2'b0,_sigX_Z_T_9}; 
  assign _sigX_Z_T_10=_sigX_Z_T_6|_GEN_23; 
  assign _GEN_24={1'b0,bitMask}; 
  assign _sigX_Z_T_12=sigX_Z|_GEN_24; 
  assign _sigX_Z_T_13=inReady ? 55'h0:_sigX_Z_T_12; 
  assign _sigX_Z_T_14=_sigX_Z_T_10|_sigX_Z_T_13; 
  assign _GEN_25={55'b0,notZeroRem_Z}; 
  assign io_inReady=idle|cycleNum[1]; 
  assign io_rawOutValid_div=cycleNum[1]&~sqrtOp_Z; 
  assign io_rawOutValid_sqrt=cycleNum[1]&sqrtOp_Z; 
  assign io_roundingModeOut=roundingMode_Z; 
  assign io_invalidExc=majorExc_Z&isNaN_Z; 
  assign io_infiniteExc=majorExc_Z&~isNaN_Z; 
  assign io_rawOut_isNaN=isNaN_Z; 
  assign io_rawOut_isInf=isInf_Z; 
  assign io_rawOut_isZero=isZero_Z; 
  assign io_rawOut_sign=sign_Z; 
  assign io_rawOut_sExp=sExp_Z; 
  assign io_rawOut_sig=_trialTerm_T_19|_GEN_25; 
  assign DivSqrtRawFN_small_1_cov_read_addr=DivSqrtRawFN_small_1_state; 
  assign DivSqrtRawFN_small_1_cov_read_data=DivSqrtRawFN_small_1_cov[DivSqrtRawFN_small_1_cov_read_addr]; 
  assign DivSqrtRawFN_small_1_cov_write_data=1'h1; 
  assign DivSqrtRawFN_small_1_cov_write_addr=DivSqrtRawFN_small_1_state; 
  assign DivSqrtRawFN_small_1_cov_write_mask=1'h1; 
  assign DivSqrtRawFN_small_1_cov_write_en=1'h1; 
  assign mux_cond_0=_T_10; 
  assign mux_cond_1=newBit; 
  assign mux_cond_2=skipCycle2; 
  assign mux_cond_3=_cycleNum_T_10; 
  assign sqrtOp_Z_shl=sqrtOp_Z; 
  assign sqrtOp_Z_pad={4'h0,sqrtOp_Z_shl}; 
  assign mux_cond_0_shl={mux_cond_0,1'h0}; 
  assign mux_cond_0_pad={3'h0,mux_cond_0_shl}; 
  assign mux_cond_1_shl={mux_cond_1,2'h0}; 
  assign mux_cond_1_pad={2'h0,mux_cond_1_shl}; 
  assign mux_cond_2_shl={mux_cond_2,3'h0}; 
  assign mux_cond_2_pad={1'h0,mux_cond_2_shl}; 
  assign mux_cond_3_shl={mux_cond_3,4'h0}; 
  assign mux_cond_3_pad=mux_cond_3_shl; 
  assign DivSqrtRawFN_small_1_xor1=sqrtOp_Z_pad^mux_cond_0_pad; 
  assign DivSqrtRawFN_small_1_xor6=mux_cond_2_pad^mux_cond_3_pad; 
  assign DivSqrtRawFN_small_1_xor2=mux_cond_1_pad^DivSqrtRawFN_small_1_xor6; 
  assign DivSqrtRawFN_small_1_xor0=DivSqrtRawFN_small_1_xor1^DivSqrtRawFN_small_1_xor2; 
  assign io_covSum=DivSqrtRawFN_small_1_covSum; 
  assign metaAssert=1'h0; initial
    begin 
    end  
  always @( posedge clock)
       begin 
         if (metaReset)
            begin 
              cycleNum <=56'h0;
            end 
          else 
            if (reset)
               begin 
                 cycleNum <=56'h1;
               end 
             else 
               if (_T_1)
                  begin 
                    cycleNum <=_cycleNum_T_15;
                  end 
         if (metaReset)
            begin 
              sqrtOp_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 sqrtOp_Z <=io_sqrtOp;
               end 
         if (metaReset)
            begin 
              majorExc_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      majorExc_Z <=_majorExc_S_T_3;
                    end 
                  else 
                    begin 
                      majorExc_Z <=_majorExc_S_T_16;
                    end 
               end 
         if (metaReset)
            begin 
              isNaN_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      isNaN_Z <=_isNaN_S_T;
                    end 
                  else 
                    begin 
                      isNaN_Z <=_isNaN_S_T_2;
                    end 
               end 
         if (metaReset)
            begin 
              isInf_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      isInf_Z <=io_a_isInf;
                    end 
                  else 
                    begin 
                      isInf_Z <=_isInf_S_T;
                    end 
               end 
         if (metaReset)
            begin 
              isZero_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 if (io_sqrtOp)
                    begin 
                      isZero_Z <=io_a_isZero;
                    end 
                  else 
                    begin 
                      isZero_Z <=_isZero_S_T;
                    end 
               end 
         if (metaReset)
            begin 
              sign_Z <=1'h0;
            end 
          else 
            if (entering)
               begin 
                 sign_Z <=sign_S;
               end 
         if (metaReset)
            begin 
              sExp_Z <=13'h0;
            end 
          else 
            if (entering_normalCase)
               begin 
                 if (io_sqrtOp)
                    begin 
                      sExp_Z <=_sExp_Z_T_1;
                    end 
                  else 
                    begin 
                      sExp_Z <=sSatExpQuot_S_div;
                    end 
               end 
         if (metaReset)
            begin 
              fractB_Z <=52'h0;
            end 
          else 
            if (_T_3)
               begin 
                 fractB_Z <=io_b_sig[51:0];
               end 
         if (metaReset)
            begin 
              roundingMode_Z <=3'h0;
            end 
          else 
            if (entering_normalCase)
               begin 
                 roundingMode_Z <=io_roundingMode;
               end 
         if (metaReset)
            begin 
              rem_Z <=55'h0;
            end 
          else 
            begin 
              rem_Z <=_GEN_10[54:0];
            end 
         if (metaReset)
            begin 
              notZeroRem_Z <=1'h0;
            end 
          else 
            if (_T_10)
               begin 
                 notZeroRem_Z <=_notZeroRem_Z_T;
               end 
         if (metaReset)
            begin 
              sigX_Z <=55'h0;
            end 
          else 
            if (_T_10)
               begin 
                 sigX_Z <=_sigX_Z_T_14;
               end 
         DivSqrtRawFN_small_1_state <=DivSqrtRawFN_small_1_xor0;
         if (!(DivSqrtRawFN_small_1_cov_read_data))
            begin 
              DivSqrtRawFN_small_1_covSum <=DivSqrtRawFN_small_1_covSum+1'h1;
            end 
       end
  
  always @( posedge clock)
       begin 
         if (DivSqrtRawFN_small_1_cov_write_en&DivSqrtRawFN_small_1_cov_write_mask)
            begin 
              DivSqrtRawFN_small_1_cov [DivSqrtRawFN_small_1_cov_write_addr]<=DivSqrtRawFN_small_1_cov_write_data;
            end 
       end
  
endmodule
 
module RoundAnyRawFNToRecFN_6 (
  input io_invalidExc,
  input io_infiniteExc,
  input io_in_isNaN,
  input io_in_isInf,
  input io_in_isZero,
  input io_in_sign,
  input [12:0] io_in_sExp,
  input [55:0] io_in_sig,
  input [2:0] io_roundingMode,
  input io_detectTininess,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output [29:0] io_covSum,
  output metaAssert) ; 
   wire roundingMode_near_even ;  
   wire roundingMode_min ;  
   wire roundingMode_max ;  
   wire roundingMode_near_maxMag ;  
   wire roundingMode_odd ;  
   wire _roundMagUp_T ;  
   wire _roundMagUp_T_2 ;  
   wire roundMagUp ;  
   wire doShiftSigDown1 ;  
   wire roundMask_msb ;  
   wire [10:0] roundMask_lsbs ;  
   wire roundMask_msb_1 ;  
   wire [9:0] roundMask_lsbs_1 ;  
   wire roundMask_msb_2 ;  
   wire [8:0] roundMask_lsbs_2 ;  
   wire roundMask_msb_3 ;  
   wire [7:0] roundMask_lsbs_3 ;  
   wire roundMask_msb_4 ;  
   wire [6:0] roundMask_lsbs_4 ;  
   wire roundMask_msb_5 ;  
   wire [5:0] roundMask_lsbs_5 ;  
   wire [64:0] roundMask_shift ;  
   wire [31:0] _roundMask_T_7 ;  
   wire [31:0] _roundMask_T_9 ;  
   wire [31:0] _roundMask_T_11 ;  
   wire [31:0] _roundMask_T_12 ;  
   wire [31:0] _GEN_0 ;  
   wire [31:0] _roundMask_T_17 ;  
   wire [31:0] _roundMask_T_19 ;  
   wire [31:0] _roundMask_T_21 ;  
   wire [31:0] _roundMask_T_22 ;  
   wire [31:0] _GEN_1 ;  
   wire [31:0] _roundMask_T_27 ;  
   wire [31:0] _roundMask_T_29 ;  
   wire [31:0] _roundMask_T_31 ;  
   wire [31:0] _roundMask_T_32 ;  
   wire [31:0] _GEN_2 ;  
   wire [31:0] _roundMask_T_37 ;  
   wire [31:0] _roundMask_T_39 ;  
   wire [31:0] _roundMask_T_41 ;  
   wire [31:0] _roundMask_T_42 ;  
   wire [31:0] _GEN_3 ;  
   wire [31:0] _roundMask_T_47 ;  
   wire [31:0] _roundMask_T_49 ;  
   wire [31:0] _roundMask_T_51 ;  
   wire [31:0] roundMask_hi ;  
   wire [15:0] _roundMask_T_57 ;  
   wire [15:0] _roundMask_T_59 ;  
   wire [15:0] _roundMask_T_61 ;  
   wire [15:0] _roundMask_T_62 ;  
   wire [15:0] _GEN_4 ;  
   wire [15:0] _roundMask_T_67 ;  
   wire [15:0] _roundMask_T_69 ;  
   wire [15:0] _roundMask_T_71 ;  
   wire [15:0] _roundMask_T_72 ;  
   wire [15:0] _GEN_5 ;  
   wire [15:0] _roundMask_T_77 ;  
   wire [15:0] _roundMask_T_79 ;  
   wire [15:0] _roundMask_T_81 ;  
   wire [15:0] _roundMask_T_82 ;  
   wire [15:0] _GEN_6 ;  
   wire [15:0] _roundMask_T_87 ;  
   wire [15:0] _roundMask_T_89 ;  
   wire [15:0] _roundMask_T_91 ;  
   wire [15:0] roundMask_hi_1 ;  
   wire roundMask_hi_2 ;  
   wire roundMask_lo ;  
   wire roundMask_lo_1 ;  
   wire [50:0] _roundMask_T_94 ;  
   wire [50:0] _roundMask_T_96 ;  
   wire [50:0] _roundMask_T_99 ;  
   wire [50:0] _roundMask_T_102 ;  
   wire [50:0] _roundMask_T_105 ;  
   wire [50:0] roundMask_hi_4 ;  
   wire [53:0] _roundMask_T_106 ;  
   wire roundMask_hi_5 ;  
   wire roundMask_lo_4 ;  
   wire roundMask_lo_5 ;  
   wire [2:0] _roundMask_T_109 ;  
   wire [2:0] _roundMask_T_110 ;  
   wire [2:0] _roundMask_T_111 ;  
   wire [2:0] _roundMask_T_112 ;  
   wire [2:0] _roundMask_T_113 ;  
   wire [53:0] _roundMask_T_114 ;  
   wire [53:0] _roundMask_T_115 ;  
   wire [53:0] _GEN_7 ;  
   wire [53:0] roundMask_hi_7 ;  
   wire [55:0] roundMask ;  
   wire [54:0] shiftedRoundMask_lo ;  
   wire [55:0] shiftedRoundMask ;  
   wire [55:0] roundPosMask ;  
   wire [55:0] _roundPosBit_T ;  
   wire roundPosBit ;  
   wire [55:0] _anyRoundExtra_T ;  
   wire anyRoundExtra ;  
   wire anyRound ;  
   wire _roundIncr_T ;  
   wire _roundIncr_T_1 ;  
   wire _roundIncr_T_2 ;  
   wire roundIncr ;  
   wire [55:0] _roundedSig_T ;  
   wire [54:0] _roundedSig_T_2 ;  
   wire _roundedSig_T_3 ;  
   wire _roundedSig_T_5 ;  
   wire [54:0] _roundedSig_T_7 ;  
   wire [54:0] _roundedSig_T_9 ;  
   wire [55:0] _roundedSig_T_11 ;  
   wire _roundedSig_T_13 ;  
   wire [54:0] _roundedSig_T_15 ;  
   wire [54:0] _GEN_8 ;  
   wire [54:0] _roundedSig_T_16 ;  
   wire [54:0] roundedSig ;  
   wire [2:0] _sRoundedExp_T_1 ;  
   wire [12:0] _GEN_9 ;  
   wire [13:0] sRoundedExp ;  
   wire [11:0] common_expOut ;  
   wire [51:0] common_fractOut ;  
   wire [3:0] _common_overflow_T ;  
   wire common_overflow ;  
   wire common_totalUnderflow ;  
   wire unboundedRange_roundPosBit ;  
   wire _unboundedRange_anyRound_T_1 ;  
   wire _unboundedRange_anyRound_T_3 ;  
   wire unboundedRange_anyRound ;  
   wire _unboundedRange_roundIncr_T_1 ;  
   wire _unboundedRange_roundIncr_T_2 ;  
   wire unboundedRange_roundIncr ;  
   wire roundCarry ;  
   wire [1:0] _common_underflow_T ;  
   wire _common_underflow_T_1 ;  
   wire _common_underflow_T_2 ;  
   wire _common_underflow_T_5 ;  
   wire _common_underflow_T_6 ;  
   wire _common_underflow_T_10 ;  
   wire _common_underflow_T_12 ;  
   wire _common_underflow_T_13 ;  
   wire _common_underflow_T_14 ;  
   wire _common_underflow_T_15 ;  
   wire _common_underflow_T_17 ;  
   wire common_underflow ;  
   wire common_inexact ;  
   wire isNaNOut ;  
   wire notNaN_isSpecialInfOut ;  
   wire _commonCase_T_2 ;  
   wire commonCase ;  
   wire overflow ;  
   wire underflow ;  
   wire _inexact_T ;  
   wire inexact ;  
   wire overflow_roundMagUp ;  
   wire _pegMinNonzeroMagOut_T ;  
   wire _pegMinNonzeroMagOut_T_1 ;  
   wire pegMinNonzeroMagOut ;  
   wire pegMaxFiniteMagOut ;  
   wire _notNaN_isInfOut_T ;  
   wire notNaN_isInfOut ;  
   wire signOut ;  
   wire _expOut_T ;  
   wire [11:0] _expOut_T_1 ;  
   wire [11:0] _expOut_T_3 ;  
   wire [11:0] _expOut_T_5 ;  
   wire [11:0] _expOut_T_7 ;  
   wire [11:0] _expOut_T_8 ;  
   wire [11:0] _expOut_T_10 ;  
   wire [11:0] _expOut_T_11 ;  
   wire [11:0] _expOut_T_13 ;  
   wire [11:0] _expOut_T_14 ;  
   wire [11:0] _expOut_T_15 ;  
   wire [11:0] _expOut_T_16 ;  
   wire [11:0] _expOut_T_17 ;  
   wire [11:0] _expOut_T_18 ;  
   wire [11:0] _expOut_T_19 ;  
   wire [11:0] _expOut_T_20 ;  
   wire [11:0] expOut ;  
   wire _fractOut_T ;  
   wire _fractOut_T_1 ;  
   wire [51:0] _fractOut_T_2 ;  
   wire [51:0] _fractOut_T_3 ;  
   wire [51:0] _fractOut_T_5 ;  
   wire [51:0] fractOut ;  
   wire [12:0] io_out_hi ;  
   wire [1:0] io_exceptionFlags_lo ;  
   wire [2:0] io_exceptionFlags_hi ;  
   wire [29:0] RoundAnyRawFNToRecFN_6_covSum ;  
  assign roundingMode_near_even=io_roundingMode==3'h0; 
  assign roundingMode_min=io_roundingMode==3'h2; 
  assign roundingMode_max=io_roundingMode==3'h3; 
  assign roundingMode_near_maxMag=io_roundingMode==3'h4; 
  assign roundingMode_odd=io_roundingMode==3'h6; 
  assign _roundMagUp_T=roundingMode_min&io_in_sign; 
  assign _roundMagUp_T_2=roundingMode_max&~io_in_sign; 
  assign roundMagUp=_roundMagUp_T|_roundMagUp_T_2; 
  assign doShiftSigDown1=io_in_sig[55]; 
  assign roundMask_msb=~io_in_sExp[11]; 
  assign roundMask_lsbs=~io_in_sExp[10:0]; 
  assign roundMask_msb_1=roundMask_lsbs[10]; 
  assign roundMask_lsbs_1=roundMask_lsbs[9:0]; 
  assign roundMask_msb_2=roundMask_lsbs_1[9]; 
  assign roundMask_lsbs_2=roundMask_lsbs_1[8:0]; 
  assign roundMask_msb_3=roundMask_lsbs_2[8]; 
  assign roundMask_lsbs_3=roundMask_lsbs_2[7:0]; 
  assign roundMask_msb_4=roundMask_lsbs_3[7]; 
  assign roundMask_lsbs_4=roundMask_lsbs_3[6:0]; 
  assign roundMask_msb_5=roundMask_lsbs_4[6]; 
  assign roundMask_lsbs_5=roundMask_lsbs_4[5:0]; 
  assign roundMask_shift=-65'sh10000000000000000>>>roundMask_lsbs_5; 
  assign _roundMask_T_7={16'b0,roundMask_shift[44:29]}; 
  assign _roundMask_T_9={roundMask_shift[28:13],16'h0}; 
  assign _roundMask_T_11=_roundMask_T_9&32'hffff0000; 
  assign _roundMask_T_12=_roundMask_T_7|_roundMask_T_11; 
  assign _GEN_0={8'b0,_roundMask_T_12[31:8]}; 
  assign _roundMask_T_17=_GEN_0&32'hff00ff; 
  assign _roundMask_T_19={_roundMask_T_12[23:0],8'h0}; 
  assign _roundMask_T_21=_roundMask_T_19&32'hff00ff00; 
  assign _roundMask_T_22=_roundMask_T_17|_roundMask_T_21; 
  assign _GEN_1={4'b0,_roundMask_T_22[31:4]}; 
  assign _roundMask_T_27=_GEN_1&32'hf0f0f0f; 
  assign _roundMask_T_29={_roundMask_T_22[27:0],4'h0}; 
  assign _roundMask_T_31=_roundMask_T_29&32'hf0f0f0f0; 
  assign _roundMask_T_32=_roundMask_T_27|_roundMask_T_31; 
  assign _GEN_2={2'b0,_roundMask_T_32[31:2]}; 
  assign _roundMask_T_37=_GEN_2&32'h33333333; 
  assign _roundMask_T_39={_roundMask_T_32[29:0],2'h0}; 
  assign _roundMask_T_41=_roundMask_T_39&32'hcccccccc; 
  assign _roundMask_T_42=_roundMask_T_37|_roundMask_T_41; 
  assign _GEN_3={1'b0,_roundMask_T_42[31:1]}; 
  assign _roundMask_T_47=_GEN_3&32'h55555555; 
  assign _roundMask_T_49={_roundMask_T_42[30:0],1'h0}; 
  assign _roundMask_T_51=_roundMask_T_49&32'haaaaaaaa; 
  assign roundMask_hi=_roundMask_T_47|_roundMask_T_51; 
  assign _roundMask_T_57={8'b0,roundMask_shift[60:53]}; 
  assign _roundMask_T_59={roundMask_shift[52:45],8'h0}; 
  assign _roundMask_T_61=_roundMask_T_59&16'hff00; 
  assign _roundMask_T_62=_roundMask_T_57|_roundMask_T_61; 
  assign _GEN_4={4'b0,_roundMask_T_62[15:4]}; 
  assign _roundMask_T_67=_GEN_4&16'hf0f; 
  assign _roundMask_T_69={_roundMask_T_62[11:0],4'h0}; 
  assign _roundMask_T_71=_roundMask_T_69&16'hf0f0; 
  assign _roundMask_T_72=_roundMask_T_67|_roundMask_T_71; 
  assign _GEN_5={2'b0,_roundMask_T_72[15:2]}; 
  assign _roundMask_T_77=_GEN_5&16'h3333; 
  assign _roundMask_T_79={_roundMask_T_72[13:0],2'h0}; 
  assign _roundMask_T_81=_roundMask_T_79&16'hcccc; 
  assign _roundMask_T_82=_roundMask_T_77|_roundMask_T_81; 
  assign _GEN_6={1'b0,_roundMask_T_82[15:1]}; 
  assign _roundMask_T_87=_GEN_6&16'h5555; 
  assign _roundMask_T_89={_roundMask_T_82[14:0],1'h0}; 
  assign _roundMask_T_91=_roundMask_T_89&16'haaaa; 
  assign roundMask_hi_1=_roundMask_T_87|_roundMask_T_91; 
  assign roundMask_hi_2=roundMask_shift[61]; 
  assign roundMask_lo=roundMask_shift[62]; 
  assign roundMask_lo_1=roundMask_shift[63]; 
  assign _roundMask_T_94={roundMask_hi,roundMask_hi_1,roundMask_hi_2,roundMask_lo,roundMask_lo_1}; 
  assign _roundMask_T_96=roundMask_msb_5 ? 51'h0:~_roundMask_T_94; 
  assign _roundMask_T_99=roundMask_msb_4 ? 51'h0:_roundMask_T_96[50:0]; 
  assign _roundMask_T_102=roundMask_msb_3 ? 51'h0:_roundMask_T_99[50:0]; 
  assign _roundMask_T_105=roundMask_msb_2 ? 51'h0:_roundMask_T_102[50:0]; 
  assign roundMask_hi_4=~_roundMask_T_105; 
  assign _roundMask_T_106={roundMask_hi_4,3'h7}; 
  assign roundMask_hi_5=roundMask_shift[0]; 
  assign roundMask_lo_4=roundMask_shift[1]; 
  assign roundMask_lo_5=roundMask_shift[2]; 
  assign _roundMask_T_109={roundMask_hi_5,roundMask_lo_4,roundMask_lo_5}; 
  assign _roundMask_T_110=roundMask_msb_5 ? _roundMask_T_109:3'h0; 
  assign _roundMask_T_111=roundMask_msb_4 ? _roundMask_T_110:3'h0; 
  assign _roundMask_T_112=roundMask_msb_3 ? _roundMask_T_111:3'h0; 
  assign _roundMask_T_113=roundMask_msb_2 ? _roundMask_T_112:3'h0; 
  assign _roundMask_T_114=roundMask_msb_1 ? _roundMask_T_106:{51'b0,_roundMask_T_113}; 
  assign _roundMask_T_115=roundMask_msb ? _roundMask_T_114:54'h0; 
  assign _GEN_7={53'b0,doShiftSigDown1}; 
  assign roundMask_hi_7=_roundMask_T_115|_GEN_7; 
  assign roundMask={roundMask_hi_7,2'h3}; 
  assign shiftedRoundMask_lo=roundMask[55:1]; 
  assign shiftedRoundMask={1'h0,shiftedRoundMask_lo}; 
  assign roundPosMask=~shiftedRoundMask&roundMask; 
  assign _roundPosBit_T=io_in_sig&roundPosMask; 
  assign roundPosBit=|_roundPosBit_T; 
  assign _anyRoundExtra_T=io_in_sig&shiftedRoundMask; 
  assign anyRoundExtra=|_anyRoundExtra_T; 
  assign anyRound=roundPosBit|anyRoundExtra; 
  assign _roundIncr_T=roundingMode_near_even|roundingMode_near_maxMag; 
  assign _roundIncr_T_1=_roundIncr_T&roundPosBit; 
  assign _roundIncr_T_2=roundMagUp&anyRound; 
  assign roundIncr=_roundIncr_T_1|_roundIncr_T_2; 
  assign _roundedSig_T=io_in_sig|roundMask; 
  assign _roundedSig_T_2=_roundedSig_T[55:2]+54'h1; 
  assign _roundedSig_T_3=roundingMode_near_even&roundPosBit; 
  assign _roundedSig_T_5=_roundedSig_T_3&~anyRoundExtra; 
  assign _roundedSig_T_7=_roundedSig_T_5 ? shiftedRoundMask_lo:55'h0; 
  assign _roundedSig_T_9=_roundedSig_T_2&~_roundedSig_T_7; 
  assign _roundedSig_T_11=io_in_sig&~roundMask; 
  assign _roundedSig_T_13=roundingMode_odd&anyRound; 
  assign _roundedSig_T_15=_roundedSig_T_13 ? roundPosMask[55:1]:55'h0; 
  assign _GEN_8={1'b0,_roundedSig_T_11[55:2]}; 
  assign _roundedSig_T_16=_GEN_8|_roundedSig_T_15; 
  assign roundedSig=roundIncr ? _roundedSig_T_9:_roundedSig_T_16; 
  assign _sRoundedExp_T_1={1'b0,$signed(roundedSig[54:53])}; 
  assign _GEN_9={{10{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; 
  assign sRoundedExp=$signed(io_in_sExp)+$signed(_GEN_9); 
  assign common_expOut=sRoundedExp[11:0]; 
  assign common_fractOut=doShiftSigDown1 ? roundedSig[52:1]:roundedSig[51:0]; 
  assign _common_overflow_T=sRoundedExp[13:10]; 
  assign common_overflow=$signed(_common_overflow_T)>=4'sh3; 
  assign common_totalUnderflow=$signed(sRoundedExp)<14'sh3ce; 
  assign unboundedRange_roundPosBit=doShiftSigDown1 ? io_in_sig[2]:io_in_sig[1]; 
  assign _unboundedRange_anyRound_T_1=doShiftSigDown1&io_in_sig[2]; 
  assign _unboundedRange_anyRound_T_3=|io_in_sig[1:0]; 
  assign unboundedRange_anyRound=_unboundedRange_anyRound_T_1|_unboundedRange_anyRound_T_3; 
  assign _unboundedRange_roundIncr_T_1=_roundIncr_T&unboundedRange_roundPosBit; 
  assign _unboundedRange_roundIncr_T_2=roundMagUp&unboundedRange_anyRound; 
  assign unboundedRange_roundIncr=_unboundedRange_roundIncr_T_1|_unboundedRange_roundIncr_T_2; 
  assign roundCarry=doShiftSigDown1 ? roundedSig[54]:roundedSig[53]; 
  assign _common_underflow_T=io_in_sExp[12:11]; 
  assign _common_underflow_T_1=$signed(_common_underflow_T)<=2'sh0; 
  assign _common_underflow_T_2=anyRound&_common_underflow_T_1; 
  assign _common_underflow_T_5=doShiftSigDown1 ? roundMask[3]:roundMask[2]; 
  assign _common_underflow_T_6=_common_underflow_T_2&_common_underflow_T_5; 
  assign _common_underflow_T_10=doShiftSigDown1 ? roundMask[4]:roundMask[3]; 
  assign _common_underflow_T_12=io_detectTininess&~_common_underflow_T_10; 
  assign _common_underflow_T_13=_common_underflow_T_12&roundCarry; 
  assign _common_underflow_T_14=_common_underflow_T_13&roundPosBit; 
  assign _common_underflow_T_15=_common_underflow_T_14&unboundedRange_roundIncr; 
  assign _common_underflow_T_17=_common_underflow_T_6&~_common_underflow_T_15; 
  assign common_underflow=common_totalUnderflow|_common_underflow_T_17; 
  assign common_inexact=common_totalUnderflow|anyRound; 
  assign isNaNOut=io_invalidExc|io_in_isNaN; 
  assign notNaN_isSpecialInfOut=io_infiniteExc|io_in_isInf; 
  assign _commonCase_T_2=~isNaNOut&~notNaN_isSpecialInfOut; 
  assign commonCase=_commonCase_T_2&~io_in_isZero; 
  assign overflow=commonCase&common_overflow; 
  assign underflow=commonCase&common_underflow; 
  assign _inexact_T=commonCase&common_inexact; 
  assign inexact=overflow|_inexact_T; 
  assign overflow_roundMagUp=_roundIncr_T|roundMagUp; 
  assign _pegMinNonzeroMagOut_T=commonCase&common_totalUnderflow; 
  assign _pegMinNonzeroMagOut_T_1=roundMagUp|roundingMode_odd; 
  assign pegMinNonzeroMagOut=_pegMinNonzeroMagOut_T&_pegMinNonzeroMagOut_T_1; 
  assign pegMaxFiniteMagOut=overflow&~overflow_roundMagUp; 
  assign _notNaN_isInfOut_T=overflow&overflow_roundMagUp; 
  assign notNaN_isInfOut=notNaN_isSpecialInfOut|_notNaN_isInfOut_T; 
  assign signOut=isNaNOut ? 1'h0:io_in_sign; 
  assign _expOut_T=io_in_isZero|common_totalUnderflow; 
  assign _expOut_T_1=_expOut_T ? 12'he00:12'h0; 
  assign _expOut_T_3=common_expOut&~_expOut_T_1; 
  assign _expOut_T_5=pegMinNonzeroMagOut ? 12'hc31:12'h0; 
  assign _expOut_T_7=_expOut_T_3&~_expOut_T_5; 
  assign _expOut_T_8=pegMaxFiniteMagOut ? 12'h400:12'h0; 
  assign _expOut_T_10=_expOut_T_7&~_expOut_T_8; 
  assign _expOut_T_11=notNaN_isInfOut ? 12'h200:12'h0; 
  assign _expOut_T_13=_expOut_T_10&~_expOut_T_11; 
  assign _expOut_T_14=pegMinNonzeroMagOut ? 12'h3ce:12'h0; 
  assign _expOut_T_15=_expOut_T_13|_expOut_T_14; 
  assign _expOut_T_16=pegMaxFiniteMagOut ? 12'hbff:12'h0; 
  assign _expOut_T_17=_expOut_T_15|_expOut_T_16; 
  assign _expOut_T_18=notNaN_isInfOut ? 12'hc00:12'h0; 
  assign _expOut_T_19=_expOut_T_17|_expOut_T_18; 
  assign _expOut_T_20=isNaNOut ? 12'he00:12'h0; 
  assign expOut=_expOut_T_19|_expOut_T_20; 
  assign _fractOut_T=isNaNOut|io_in_isZero; 
  assign _fractOut_T_1=_fractOut_T|common_totalUnderflow; 
  assign _fractOut_T_2=isNaNOut ? 52'h8000000000000:52'h0; 
  assign _fractOut_T_3=_fractOut_T_1 ? _fractOut_T_2:common_fractOut; 
  assign _fractOut_T_5=pegMaxFiniteMagOut ? 52'hfffffffffffff:52'h0; 
  assign fractOut=_fractOut_T_3|_fractOut_T_5; 
  assign io_out_hi={signOut,expOut}; 
  assign io_exceptionFlags_lo={underflow,inexact}; 
  assign io_exceptionFlags_hi={io_invalidExc,io_infiniteExc,overflow}; 
  assign io_out={io_out_hi,fractOut}; 
  assign io_exceptionFlags={io_exceptionFlags_hi,io_exceptionFlags_lo}; 
  assign RoundAnyRawFNToRecFN_6_covSum=30'h0; 
  assign io_covSum=RoundAnyRawFNToRecFN_6_covSum; 
  assign metaAssert=1'h0; 
endmodule
 




