module IntXbar (
  input auto_int_in_0,
  input auto_int_in_1,
  output auto_int_out_0,
  output auto_int_out_1) ; 
  assign auto_int_out_0=auto_int_in_0; 
  assign auto_int_out_1=auto_int_in_1; 
endmodule
 
module NonSyncResetSynchronizerPrimitiveShiftReg_d3 (
  input clock,
  input io_d,
  output io_q) ; 
   reg sync_0 ;  
   reg sync_1 ;  
   reg sync_2 ;  
  always @( posedge clock)
       begin 
         sync_0 <=sync_1;
         sync_1 <=sync_2;
         sync_2 <=io_d;
       end
  
  assign io_q=sync_0; 
endmodule
 
module SynchronizerShiftReg_w2_d3 (
  input clock,
  input [1:0] io_d,
  output [1:0] io_q) ; 
   wire _output_chain_1_io_q ;  
   wire _output_chain_io_q ;  
  NonSyncResetSynchronizerPrimitiveShiftReg_d3 output_chain(.clock(clock),.io_d(io_d[0]),.io_q(_output_chain_io_q)); 
  NonSyncResetSynchronizerPrimitiveShiftReg_d3 output_chain_1(.clock(clock),.io_d(io_d[1]),.io_q(_output_chain_1_io_q)); 
  assign io_q={_output_chain_1_io_q,_output_chain_io_q}; 
endmodule
 
module IntSyncAsyncCrossingSink (
  input clock,
  input auto_in_sync_0,
  input auto_in_sync_1,
  output auto_out_0,
  output auto_out_1) ; 
   wire [1:0] _chain_io_q ;  
  SynchronizerShiftReg_w2_d3 chain(.clock(clock),.io_d({auto_in_sync_1,auto_in_sync_0}),.io_q(_chain_io_q)); 
  assign auto_out_0=_chain_io_q[0]; 
  assign auto_out_1=_chain_io_q[1]; 
endmodule
 
module SimpleClockGroupSource (
  input clock,
  input reset,
  output auto_out_member_subsystem_sbus_5_clock,
  output auto_out_member_subsystem_sbus_5_reset,
  output auto_out_member_subsystem_sbus_4_clock,
  output auto_out_member_subsystem_sbus_4_reset,
  output auto_out_member_subsystem_sbus_3_clock,
  output auto_out_member_subsystem_sbus_3_reset,
  output auto_out_member_subsystem_sbus_2_clock,
  output auto_out_member_subsystem_sbus_2_reset,
  output auto_out_member_subsystem_sbus_1_clock,
  output auto_out_member_subsystem_sbus_1_reset,
  output auto_out_member_subsystem_sbus_0_clock,
  output auto_out_member_subsystem_sbus_0_reset) ; 
  assign auto_out_member_subsystem_sbus_5_clock=clock; 
  assign auto_out_member_subsystem_sbus_5_reset=reset; 
  assign auto_out_member_subsystem_sbus_4_clock=clock; 
  assign auto_out_member_subsystem_sbus_4_reset=reset; 
  assign auto_out_member_subsystem_sbus_3_clock=clock; 
  assign auto_out_member_subsystem_sbus_3_reset=reset; 
  assign auto_out_member_subsystem_sbus_2_clock=clock; 
  assign auto_out_member_subsystem_sbus_2_reset=reset; 
  assign auto_out_member_subsystem_sbus_1_clock=clock; 
  assign auto_out_member_subsystem_sbus_1_reset=reset; 
  assign auto_out_member_subsystem_sbus_0_clock=clock; 
  assign auto_out_member_subsystem_sbus_0_reset=reset; 
endmodule
 
module FixedClockBroadcast (
  input auto_in_clock,
  input auto_in_reset,
  output auto_out_2_clock,
  output auto_out_2_reset,
  output auto_out_1_clock,
  output auto_out_0_clock,
  output auto_out_0_reset) ; 
  assign auto_out_2_clock=auto_in_clock; 
  assign auto_out_2_reset=auto_in_reset; 
  assign auto_out_1_clock=auto_in_clock; 
  assign auto_out_0_clock=auto_in_clock; 
  assign auto_out_0_reset=auto_in_reset; 
endmodule
 
module TLMonitor (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [3:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [3:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [3:0] source ;  
   reg [31:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [3:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [15:0] inflight ;  
   reg [63:0] inflight_opcodes ;  
   reg [127:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [63:0] _a_opcode_lookup_T_1=inflight_opcodes>>{58'h0,io_in_d_bits_source,2'h0} ;  
   wire [15:0] _GEN_0={12'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [15:0] _GEN_2={12'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [15:0] inflight_1 ;  
   reg [127:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_bits_size<4'h7 ;  
   wire _GEN_6=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_7=_GEN_4&_GEN_5&_GEN_6 ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_9=io_in_a_bits_param>3'h2 ;  
   wire _GEN_10=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_11=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_13={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_14=_GEN_4&_GEN_13 ;  
   wire _GEN_15=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_16={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_17={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_18={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_19=io_in_a_bits_mask!=mask ;  
   wire _GEN_20=_GEN_4&(_GEN_14|_GEN_5&(_GEN_15|_GEN_16|_GEN_17|_GEN_6)|io_in_a_bits_size<4'h9&_GEN_18) ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_22=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_23=_GEN_4&io_in_a_bits_size<4'h4&(_GEN_15|_GEN_13|_GEN_16|_GEN_17) ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_26=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_27=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_28=io_in_d_bits_size<4'h3 ;  
   wire _GEN_29=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_30=io_in_d_bits_param==2'h2 ;  
   wire _GEN_31=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_32=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_33=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_35=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_36=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_37=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [127:0] _GEN_38={121'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [15:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 16'h1<<_GEN_0:16'h0 ;  
   wire _GEN_39=io_in_d_valid&d_first_1 ;  
   wire _GEN_40=_GEN_39&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_41=_GEN_40&same_cycle_resp&~reset ;  
   wire _GEN_42=_GEN_40&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_43={4'h0,io_in_d_bits_size} ;  
   wire _GEN_44=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [15:0] _GEN_45=inflight>>_GEN_0 ;  
   wire [15:0] _GEN_46=inflight>>_GEN_2 ;  
   wire [127:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_38 ;  
   wire [15:0] _GEN_47=inflight_1>>_GEN_2 ;  
   wire [127:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_38 ;  
  always @( posedge clock)
       begin 
         if (_GEN_8&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~(_GEN_14|_GEN_5&(_GEN_15|{io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0|_GEN_16|_GEN_17|_GEN_18|_GEN_6)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(_GEN_4&_GEN_14))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_45[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~reset&~(_GEN_46[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_43!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_40 ? 16'h1<<_GEN_2:16'h0)|a_set_wo_ready==16'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==16'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~(_GEN_47[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&_GEN_43!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==16'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_48={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_48 ;  
   wire [142:0] _GEN_49={136'h0,io_in_d_bits_source,3'h0} ;  
   wire [142:0] _d_opcodes_clr_T_5=143'hF<<{137'h0,io_in_d_bits_source,2'h0} ;  
   wire [130:0] _a_opcodes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{125'h0,io_in_a_bits_source,2'h0} ;  
   wire [142:0] _d_sizes_clr_T_5=143'hFF<<_GEN_49 ;  
   wire [131:0] _a_sizes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{125'h0,io_in_a_bits_source,3'h0} ;  
   wire [142:0] _d_sizes_clr_T_11=143'hFF<<_GEN_49 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_50=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_51=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=16'h0;
              inflight_opcodes <=64'h0;
              inflight_sizes <=128'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=16'h0;
              inflight_sizes_1 <=128'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? 16'h1<<_GEN_0:16'h0))&~(_GEN_50 ? 16'h1<<_GEN_2:16'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[63:0]:64'h0))&~(_GEN_50 ? _d_opcodes_clr_T_5[63:0]:64'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[127:0]:128'h0))&~(_GEN_50 ? _d_sizes_clr_T_5[127:0]:128'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_51 ? 16'h1<<_GEN_2:16'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_51 ? _d_sizes_clr_T_11[127:0]:128'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLMonitor_1 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [1:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_b_ready,
  input io_in_b_valid,
  input [1:0] io_in_b_bits_param,
  input [31:0] io_in_b_bits_address,
  input io_in_c_ready,
  input io_in_c_valid,
  input [2:0] io_in_c_bits_opcode,
  input [2:0] io_in_c_bits_param,
  input [3:0] io_in_c_bits_size,
  input [1:0] io_in_c_bits_source,
  input [31:0] io_in_c_bits_address,
  input io_in_c_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [1:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt,
  input io_in_e_valid,
  input [1:0] io_in_e_bits_sink) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire [26:0] _GEN_0={23'h0,io_in_c_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [1:0] source ;  
   reg [31:0] address ;  
   wire _d_first_T_3=io_in_d_ready&io_in_d_valid ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [1:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [8:0] b_first_counter ;  
   reg [1:0] param_2 ;  
   reg [31:0] address_1 ;  
   wire _c_first_T_1=io_in_c_ready&io_in_c_valid ;  
   reg [8:0] c_first_counter ;  
   reg [2:0] opcode_3 ;  
   reg [2:0] param_3 ;  
   reg [3:0] size_3 ;  
   reg [1:0] source_3 ;  
   reg [31:0] address_2 ;  
   reg [2:0] inflight ;  
   reg [11:0] inflight_opcodes ;  
   reg [23:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [11:0] _a_opcode_lookup_T_1=inflight_opcodes>>{8'h0,io_in_d_bits_source,2'h0} ;  
   wire [3:0] _GEN_1={2'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [3:0] _GEN_3={2'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [2:0] inflight_1 ;  
   reg [23:0] inflight_sizes_1 ;  
   reg [8:0] c_first_counter_1 ;  
   wire c_first_1=c_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   wire _GEN_4=io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1] ;  
   wire [3:0] _GEN_5={2'h0,io_in_c_bits_source} ;  
   wire _GEN_6=_c_first_T_1&c_first_1&_GEN_4 ;  
   reg [31:0] watchdog_1 ;  
   reg [3:0] inflight_2 ;  
   reg [8:0] d_first_counter_3 ;  
   wire d_first_3=d_first_counter_3==9'h0 ;  
   wire _GEN_7=_d_first_T_3&d_first_3&io_in_d_bits_opcode[2]&~(io_in_d_bits_opcode[1]) ;  
   wire [3:0] _GEN_8={2'h0,io_in_d_bits_sink} ;  
   wire [3:0] d_set=_GEN_7 ? 4'h1<<_GEN_8:4'h0 ;  
   wire [3:0] _GEN_9={2'h0,io_in_e_bits_sink} ;  
   wire _source_ok_T=io_in_a_bits_source==2'h0 ;  
   wire _source_ok_T_1=io_in_a_bits_source==2'h1 ;  
   wire _source_ok_T_2=io_in_a_bits_source==2'h2 ;  
   wire source_ok=_source_ok_T|_source_ok_T_1|_source_ok_T_2 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_10=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_11=io_in_a_bits_size<4'hD ;  
   wire _GEN_12=_GEN_11&(_source_ok_T|_source_ok_T_1|_source_ok_T_2) ;  
   wire _GEN_13=io_in_a_bits_size<4'h7 ;  
   wire _GEN_14=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_15=_GEN_12&_GEN_13&_GEN_14 ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_17=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_18={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_19={io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0 ;  
   wire _GEN_20={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_21={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_22={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_23=_GEN_17|_GEN_18 ;  
   wire _GEN_24=_source_ok_T&io_in_a_bits_size==4'h6&_GEN_11&(_GEN_23|_GEN_19|_GEN_20|_GEN_21|_GEN_22|_GEN_14) ;  
   wire _GEN_25=io_in_a_bits_param>3'h2 ;  
   wire _GEN_26=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_27=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_28=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_29=_GEN_11&_GEN_18 ;  
   wire _GEN_30=io_in_a_bits_mask!=mask ;  
   wire _GEN_31=_GEN_12&(_GEN_29|_GEN_13&(_GEN_17|_GEN_20|_GEN_21|_GEN_14)|io_in_a_bits_size<4'h9&_GEN_22) ;  
   wire _GEN_32=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_33=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_34=_GEN_12&io_in_a_bits_size<4'h4&(_GEN_23|_GEN_20|_GEN_21) ;  
   wire _GEN_35=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_36=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_37=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source==2'h0|io_in_d_bits_source==2'h1|io_in_d_bits_source==2'h2 ;  
   wire _GEN_38=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_39=io_in_d_bits_size<4'h3 ;  
   wire _GEN_40=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_41=io_in_d_bits_param==2'h2 ;  
   wire _GEN_42=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_43=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_44=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_45=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_46=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire [19:0] _GEN_47={io_in_b_bits_address[31:14],~(io_in_b_bits_address[13:12])} ;  
   wire [5:0] _GEN_48={io_in_b_bits_address[31:28],~(io_in_b_bits_address[27:26])} ;  
   wire [15:0] _GEN_49={io_in_b_bits_address[31:26],io_in_b_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_50={io_in_b_bits_address[31:17],~(io_in_b_bits_address[16])} ;  
   wire _GEN_51=io_in_b_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_52={io_in_b_bits_address[31],~(io_in_b_bits_address[30:29])} ;  
   wire _GEN_53=io_in_b_valid&~reset ;  
   wire _source_ok_T_8=io_in_c_bits_source==2'h0 ;  
   wire _source_ok_T_9=io_in_c_bits_source==2'h1 ;  
   wire _source_ok_T_10=io_in_c_bits_source==2'h2 ;  
   wire source_ok_2=_source_ok_T_8|_source_ok_T_9|_source_ok_T_10 ;  
   wire [26:0] _is_aligned_mask_T_7=27'hFFF<<_GEN_0 ;  
   wire [11:0] _GEN_54=io_in_c_bits_address[11:0]&~(_is_aligned_mask_T_7[11:0]) ;  
   wire [19:0] _GEN_55={io_in_c_bits_address[31:14],~(io_in_c_bits_address[13:12])} ;  
   wire [5:0] _GEN_56={io_in_c_bits_address[31:28],~(io_in_c_bits_address[27:26])} ;  
   wire [15:0] _GEN_57={io_in_c_bits_address[31:26],io_in_c_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_58={io_in_c_bits_address[31:17],~(io_in_c_bits_address[16])} ;  
   wire _GEN_59=io_in_c_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_60={io_in_c_bits_address[31],~(io_in_c_bits_address[30:29])} ;  
   wire address_ok_1=~(|_GEN_55)|~(|_GEN_56)|~(|_GEN_57)|~(|(io_in_c_bits_address[31:12]))|~(|_GEN_58)|~_GEN_59|~(|_GEN_60) ;  
   wire _GEN_61=io_in_c_valid&io_in_c_bits_opcode==3'h4&~reset ;  
   wire _GEN_62=io_in_c_bits_size<4'h3 ;  
   wire _GEN_63=io_in_c_valid&io_in_c_bits_opcode==3'h5&~reset ;  
   wire _GEN_64=io_in_c_bits_size<4'hD ;  
   wire _GEN_65=_GEN_64&(_source_ok_T_8|_source_ok_T_9|_source_ok_T_10)&io_in_c_bits_size<4'h7&~_GEN_59 ;  
   wire _GEN_66=io_in_c_valid&io_in_c_bits_opcode==3'h6&~reset ;  
   wire _GEN_67=_source_ok_T_8&io_in_c_bits_size==4'h6&_GEN_64&(~(|(io_in_c_bits_address[31:12]))|~(|_GEN_55)|~(|_GEN_58)|~(|_GEN_57)|~(|_GEN_56)|~(|_GEN_60)|~_GEN_59) ;  
   wire _GEN_68=io_in_c_valid&(&io_in_c_bits_opcode)&~reset ;  
   wire _GEN_69=io_in_c_valid&io_in_c_bits_opcode==3'h0&~reset ;  
   wire _GEN_70=io_in_c_valid&io_in_c_bits_opcode==3'h1&~reset ;  
   wire _GEN_71=io_in_c_valid&io_in_c_bits_opcode==3'h2&~reset ;  
   wire _GEN_72=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_73=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_74=io_in_b_valid&(|b_first_counter)&~reset ;  
   wire _GEN_75=io_in_c_valid&(|c_first_counter)&~reset ;  
   wire [23:0] _GEN_76={19'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [3:0] _a_set_wo_ready_T=4'h1<<_GEN_1 ;  
   wire [2:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[2:0]:3'h0 ;  
   wire _GEN_77=io_in_d_valid&d_first_1 ;  
   wire _GEN_78=_GEN_77&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [2:0] _GEN_79={1'h0,io_in_d_bits_source} ;  
   wire _GEN_80=_GEN_78&same_cycle_resp&~reset ;  
   wire _GEN_81=_GEN_78&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_82={4'h0,io_in_d_bits_size} ;  
   wire _same_cycle_resp_T_3=io_in_c_valid&c_first_1 ;  
   wire [3:0] _c_set_wo_ready_T=4'h1<<_GEN_5 ;  
   wire [2:0] c_set_wo_ready=_same_cycle_resp_T_3&_GEN_4 ? _c_set_wo_ready_T[2:0]:3'h0 ;  
   wire _GEN_83=io_in_d_valid&d_first_2 ;  
   wire _GEN_84=_GEN_83&d_release_ack ;  
   wire same_cycle_resp_1=_same_cycle_resp_T_3&io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1]&io_in_c_bits_source==io_in_d_bits_source ;  
   wire [2:0] _GEN_85=inflight>>io_in_a_bits_source ;  
   wire [2:0] _GEN_86=inflight>>_GEN_79 ;  
   wire [23:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_76 ;  
   wire [3:0] _d_clr_wo_ready_T=4'h1<<_GEN_3 ;  
   wire [2:0] _GEN_87=inflight_1>>io_in_c_bits_source ;  
   wire [2:0] _GEN_88=inflight_1>>_GEN_79 ;  
   wire [23:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_76 ;  
   wire [3:0] _d_clr_wo_ready_T_1=4'h1<<_GEN_3 ;  
   wire [3:0] _GEN_89=inflight_2>>_GEN_8 ;  
   wire [3:0] _GEN_90=(d_set|inflight_2)>>_GEN_9 ;  
  always @( posedge clock)
       begin 
         if (_GEN_16&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(_GEN_29|_GEN_13&(_GEN_17|_GEN_19|_GEN_20|_GEN_21|_GEN_22|_GEN_14)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~_GEN_34)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~_GEN_34)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~(_GEN_12&_GEN_29))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&~(~(|(io_in_b_bits_address[31:12]))|~(|_GEN_47)|~(|_GEN_50)|~(|_GEN_49)|~(|_GEN_48)|~(|_GEN_52)|~_GEN_51))
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&~(~(|_GEN_47)|~(|_GEN_48)|~(|_GEN_49)|~(|(io_in_b_bits_address[31:12]))|~(|_GEN_50)|~_GEN_51|~(|_GEN_52)))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&(|(io_in_b_bits_address[5:0])))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&(&io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&~_GEN_65)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&~_GEN_67)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&~_GEN_65)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&~_GEN_67)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&io_in_b_bits_param!=param_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&io_in_b_bits_address!=address_1)
            begin 
              if (1)$display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_opcode!=opcode_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_param!=param_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_size!=size_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_source!=source_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_address!=address_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel address changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_85[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&~reset&~(_GEN_86[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&_GEN_82!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_77&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_78 ? _d_clr_wo_ready_T[2:0]:3'h0)|a_set_wo_ready==3'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==3'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~reset&_GEN_87[0])
            begin 
              if (1)$display("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&~reset&~(_GEN_88[0]|same_cycle_resp_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&same_cycle_resp_1&~reset&io_in_d_bits_size!=io_in_c_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&~same_cycle_resp_1&~reset&_GEN_82!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&c_first_1&io_in_c_valid&io_in_c_bits_source==io_in_d_bits_source&d_release_ack&~(io_in_c_bits_opcode==3'h4|io_in_c_bits_opcode==3'h5)&~reset&~(~io_in_d_ready|io_in_c_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if ((|c_set_wo_ready)&~reset&c_set_wo_ready==(_GEN_84 ? _d_clr_wo_ready_T_1[2:0]:3'h0))
            begin 
              if (1)$display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==3'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~reset&_GEN_89[0])
            begin 
              if (1)$display("Assertion failed: 'D' channel re-used a sink ID (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_e_valid&~reset&~(_GEN_90[0]))
            begin 
              if (1)$display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:55)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_91={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_91 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_91 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_91 ;  
   wire [26:0] _d_first_beats1_decode_T_13=27'hFFF<<_GEN_91 ;  
   wire [26:0] _c_first_beats1_decode_T_1=27'hFFF<<_GEN_0 ;  
   wire [26:0] _c_first_beats1_decode_T_5=27'hFFF<<_GEN_0 ;  
   wire _GEN_92=_d_first_T_3&d_first_1&~d_release_ack ;  
   wire [46:0] _GEN_93={42'h0,io_in_d_bits_source,3'h0} ;  
   wire _GEN_94=_d_first_T_3&d_first_2&d_release_ack ;  
   wire [3:0] _d_clr_T=4'h1<<_GEN_3 ;  
   wire [3:0] _a_set_T=4'h1<<_GEN_1 ;  
   wire [46:0] _d_opcodes_clr_T_5=47'hF<<{43'h0,io_in_d_bits_source,2'h0} ;  
   wire [34:0] _a_opcodes_set_T_1={31'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{31'h0,io_in_a_bits_source,2'h0} ;  
   wire [46:0] _d_sizes_clr_T_5=47'hFF<<_GEN_93 ;  
   wire [35:0] _a_sizes_set_T_1={31'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:5'h0}<<{31'h0,io_in_a_bits_source,3'h0} ;  
   wire [3:0] _d_clr_T_1=4'h1<<_GEN_3 ;  
   wire [3:0] _c_set_T=4'h1<<_GEN_5 ;  
   wire [46:0] _d_sizes_clr_T_11=47'hFF<<_GEN_93 ;  
   wire [35:0] _c_sizes_set_T_1={31'h0,_GEN_6 ? {io_in_c_bits_size,1'h1}:5'h0}<<{31'h0,io_in_c_bits_source,3'h0} ;  
   wire b_first_done=io_in_b_ready&io_in_b_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              b_first_counter <=9'h0;
              c_first_counter <=9'h0;
              inflight <=3'h0;
              inflight_opcodes <=12'h0;
              inflight_sizes <=24'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=3'h0;
              inflight_sizes_1 <=24'h0;
              c_first_counter_1 <=9'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
              inflight_2 <=4'h0;
              d_first_counter_3 <=9'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_3)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   if (d_first_3)
                      d_first_counter_3 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_13[11:3]):9'h0;
                    else 
                      d_first_counter_3 <=d_first_counter_3-9'h1;
                 end 
              if (b_first_done)
                 begin 
                   if (|b_first_counter)
                      b_first_counter <=b_first_counter-9'h1;
                    else 
                      b_first_counter <=9'h0;
                 end 
              if (_c_first_T_1)
                 begin 
                   if (|c_first_counter)
                      c_first_counter <=c_first_counter-9'h1;
                    else 
                      c_first_counter <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_1[11:3]):9'h0;
                   if (c_first_1)
                      c_first_counter_1 <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      c_first_counter_1 <=c_first_counter_1-9'h1;
                 end 
              inflight <=(inflight|(_GEN_2 ? _a_set_T[2:0]:3'h0))&~(_GEN_92 ? _d_clr_T[2:0]:3'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[11:0]:12'h0))&~(_GEN_92 ? _d_opcodes_clr_T_5[11:0]:12'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[23:0]:24'h0))&~(_GEN_92 ? _d_sizes_clr_T_5[23:0]:24'h0);
              if (_a_first_T_1|_d_first_T_3)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=(inflight_1|(_GEN_6 ? _c_set_T[2:0]:3'h0))&~(_GEN_94 ? _d_clr_T_1[2:0]:3'h0);
              inflight_sizes_1 <=(inflight_sizes_1|(_GEN_6 ? _c_sizes_set_T_1[23:0]:24'h0))&~(_GEN_94 ? _d_sizes_clr_T_11[23:0]:24'h0);
              if (_c_first_T_1|_d_first_T_3)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight_2 <=(inflight_2|d_set)&~(io_in_e_valid ? 4'h1<<_GEN_9:4'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_3&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
         if (b_first_done&~(|b_first_counter))
            begin 
              param_2 <=io_in_b_bits_param;
              address_1 <=io_in_b_bits_address;
            end 
         if (_c_first_T_1&~(|c_first_counter))
            begin 
              opcode_3 <=io_in_c_bits_opcode;
              param_3 <=io_in_c_bits_param;
              size_3 <=io_in_c_bits_size;
              source_3 <=io_in_c_bits_source;
              address_2 <=io_in_c_bits_address;
            end 
       end
  
endmodule
 
module TLXbar (
  input clock,
  input reset,
  output auto_in_1_a_ready,
  input auto_in_1_a_valid,
  input [2:0] auto_in_1_a_bits_opcode,
  input [2:0] auto_in_1_a_bits_param,
  input [3:0] auto_in_1_a_bits_size,
  input [1:0] auto_in_1_a_bits_source,
  input [31:0] auto_in_1_a_bits_address,
  input [7:0] auto_in_1_a_bits_mask,
  input [63:0] auto_in_1_a_bits_data,
  input auto_in_1_a_bits_corrupt,
  input auto_in_1_b_ready,
  output auto_in_1_b_valid,
  output [1:0] auto_in_1_b_bits_param,
  output [31:0] auto_in_1_b_bits_address,
  output auto_in_1_c_ready,
  input auto_in_1_c_valid,
  input [2:0] auto_in_1_c_bits_opcode,
  input [2:0] auto_in_1_c_bits_param,
  input [3:0] auto_in_1_c_bits_size,
  input [1:0] auto_in_1_c_bits_source,
  input [31:0] auto_in_1_c_bits_address,
  input [63:0] auto_in_1_c_bits_data,
  input auto_in_1_c_bits_corrupt,
  input auto_in_1_d_ready,
  output auto_in_1_d_valid,
  output [2:0] auto_in_1_d_bits_opcode,
  output [1:0] auto_in_1_d_bits_param,
  output [3:0] auto_in_1_d_bits_size,
  output [1:0] auto_in_1_d_bits_source,
  output [1:0] auto_in_1_d_bits_sink,
  output auto_in_1_d_bits_denied,
  output [63:0] auto_in_1_d_bits_data,
  output auto_in_1_d_bits_corrupt,
  input auto_in_1_e_valid,
  input [1:0] auto_in_1_e_bits_sink,
  output auto_in_0_a_ready,
  input auto_in_0_a_valid,
  input [2:0] auto_in_0_a_bits_opcode,
  input [2:0] auto_in_0_a_bits_param,
  input [3:0] auto_in_0_a_bits_size,
  input [3:0] auto_in_0_a_bits_source,
  input [31:0] auto_in_0_a_bits_address,
  input [7:0] auto_in_0_a_bits_mask,
  input [63:0] auto_in_0_a_bits_data,
  input auto_in_0_a_bits_corrupt,
  input auto_in_0_d_ready,
  output auto_in_0_d_valid,
  output [2:0] auto_in_0_d_bits_opcode,
  output [1:0] auto_in_0_d_bits_param,
  output [3:0] auto_in_0_d_bits_size,
  output [3:0] auto_in_0_d_bits_source,
  output [1:0] auto_in_0_d_bits_sink,
  output auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output auto_in_0_d_bits_corrupt,
  input auto_out_2_a_ready,
  output auto_out_2_a_valid,
  output [2:0] auto_out_2_a_bits_opcode,
  output [2:0] auto_out_2_a_bits_param,
  output [3:0] auto_out_2_a_bits_size,
  output [4:0] auto_out_2_a_bits_source,
  output [30:0] auto_out_2_a_bits_address,
  output [7:0] auto_out_2_a_bits_mask,
  output [63:0] auto_out_2_a_bits_data,
  output auto_out_2_a_bits_corrupt,
  output auto_out_2_d_ready,
  input auto_out_2_d_valid,
  input [2:0] auto_out_2_d_bits_opcode,
  input [3:0] auto_out_2_d_bits_size,
  input [4:0] auto_out_2_d_bits_source,
  input auto_out_2_d_bits_denied,
  input [63:0] auto_out_2_d_bits_data,
  input auto_out_2_d_bits_corrupt,
  input auto_out_1_a_ready,
  output auto_out_1_a_valid,
  output [2:0] auto_out_1_a_bits_opcode,
  output [2:0] auto_out_1_a_bits_param,
  output [2:0] auto_out_1_a_bits_size,
  output [4:0] auto_out_1_a_bits_source,
  output [31:0] auto_out_1_a_bits_address,
  output [7:0] auto_out_1_a_bits_mask,
  output [63:0] auto_out_1_a_bits_data,
  output auto_out_1_a_bits_corrupt,
  output auto_out_1_b_ready,
  input auto_out_1_b_valid,
  input [1:0] auto_out_1_b_bits_param,
  input [31:0] auto_out_1_b_bits_address,
  input auto_out_1_c_ready,
  output auto_out_1_c_valid,
  output [2:0] auto_out_1_c_bits_opcode,
  output [2:0] auto_out_1_c_bits_param,
  output [2:0] auto_out_1_c_bits_size,
  output [4:0] auto_out_1_c_bits_source,
  output [31:0] auto_out_1_c_bits_address,
  output [63:0] auto_out_1_c_bits_data,
  output auto_out_1_c_bits_corrupt,
  output auto_out_1_d_ready,
  input auto_out_1_d_valid,
  input [2:0] auto_out_1_d_bits_opcode,
  input [1:0] auto_out_1_d_bits_param,
  input [2:0] auto_out_1_d_bits_size,
  input [4:0] auto_out_1_d_bits_source,
  input [1:0] auto_out_1_d_bits_sink,
  input auto_out_1_d_bits_denied,
  input [63:0] auto_out_1_d_bits_data,
  input auto_out_1_d_bits_corrupt,
  output auto_out_1_e_valid,
  output [1:0] auto_out_1_e_bits_sink,
  input auto_out_0_a_ready,
  output auto_out_0_a_valid,
  output [2:0] auto_out_0_a_bits_opcode,
  output [2:0] auto_out_0_a_bits_param,
  output [3:0] auto_out_0_a_bits_size,
  output [4:0] auto_out_0_a_bits_source,
  output [27:0] auto_out_0_a_bits_address,
  output [7:0] auto_out_0_a_bits_mask,
  output [63:0] auto_out_0_a_bits_data,
  output auto_out_0_a_bits_corrupt,
  output auto_out_0_d_ready,
  input auto_out_0_d_valid,
  input [2:0] auto_out_0_d_bits_opcode,
  input [1:0] auto_out_0_d_bits_param,
  input [3:0] auto_out_0_d_bits_size,
  input [4:0] auto_out_0_d_bits_source,
  input auto_out_0_d_bits_sink,
  input auto_out_0_d_bits_denied,
  input [63:0] auto_out_0_d_bits_data,
  input auto_out_0_d_bits_corrupt) ; 
   wire allowed_4_2 ;  
   wire allowed_4_1 ;  
   wire allowed_4_0 ;  
   wire allowed_3_2 ;  
   wire allowed_3_1 ;  
   wire allowed_3_0 ;  
   wire allowed_2_1 ;  
   wire allowed_2_0 ;  
   wire allowed_1_1 ;  
   wire allowed_1_0 ;  
   wire allowed_1 ;  
   wire allowed_0 ;  
   wire [4:0] in_0_a_bits_source={1'h0,auto_in_0_a_bits_source} ;  
   wire [4:0] in_1_a_bits_source={3'h4,auto_in_1_a_bits_source} ;  
   wire [1:0] out_0_d_bits_sink={1'h0,auto_out_0_d_bits_sink} ;  
   wire [3:0] out_1_d_bits_size={1'h0,auto_out_1_d_bits_size} ;  
   wire requestAIO_0_0=auto_in_0_a_bits_address[31:30]==2'h0 ;  
   wire requestAIO_0_1=auto_in_0_a_bits_address[31:30]==2'h2 ;  
   wire requestAIO_0_2={auto_in_0_a_bits_address[31],~(auto_in_0_a_bits_address[30])}==2'h0 ;  
   wire requestAIO_1_0=auto_in_1_a_bits_address[31:30]==2'h0 ;  
   wire requestAIO_1_1=auto_in_1_a_bits_address[31:30]==2'h2 ;  
   wire requestAIO_1_2={auto_in_1_a_bits_address[31],~(auto_in_1_a_bits_address[30])}==2'h0 ;  
   wire requestDOI_0_1=auto_out_0_d_bits_source[4:2]==3'h4 ;  
   wire requestDOI_1_1=auto_out_1_d_bits_source[4:2]==3'h4 ;  
   wire requestDOI_2_1=auto_out_2_d_bits_source[4:2]==3'h4 ;  
   wire portsAOI_filtered_0_valid=auto_in_0_a_valid&requestAIO_0_0 ;  
   wire portsAOI_filtered_1_valid=auto_in_0_a_valid&requestAIO_0_1 ;  
   wire portsAOI_filtered_2_valid=auto_in_0_a_valid&requestAIO_0_2 ;  
   wire _portsAOI_in_0_a_ready_T_4=requestAIO_0_0&auto_out_0_a_ready&allowed_0|requestAIO_0_1&auto_out_1_a_ready&allowed_1_0|requestAIO_0_2&auto_out_2_a_ready&allowed_2_0 ;  
   wire portsAOI_filtered_1_0_valid=auto_in_1_a_valid&requestAIO_1_0 ;  
   wire portsAOI_filtered_1_1_valid=auto_in_1_a_valid&requestAIO_1_1 ;  
   wire portsAOI_filtered_1_2_valid=auto_in_1_a_valid&requestAIO_1_2 ;  
   wire _portsAOI_in_1_a_ready_T_4=requestAIO_1_0&auto_out_0_a_ready&allowed_1|requestAIO_1_1&auto_out_1_a_ready&allowed_1_1|requestAIO_1_2&auto_out_2_a_ready&allowed_2_1 ;  
   wire portsDIO_filtered_0_valid=auto_out_0_d_valid&~(auto_out_0_d_bits_source[4]) ;  
   wire portsDIO_filtered_1_valid=auto_out_0_d_valid&requestDOI_0_1 ;  
   wire portsDIO_filtered_1_0_valid=auto_out_1_d_valid&~(auto_out_1_d_bits_source[4]) ;  
   wire portsDIO_filtered_1_1_valid=auto_out_1_d_valid&requestDOI_1_1 ;  
   wire portsDIO_filtered_2_0_valid=auto_out_2_d_valid&~(auto_out_2_d_bits_source[4]) ;  
   wire portsDIO_filtered_2_1_valid=auto_out_2_d_valid&requestDOI_2_1 ;  
   reg [8:0] beatsLeft ;  
   wire idle=beatsLeft==9'h0 ;  
   wire [1:0] readys_valid={portsAOI_filtered_1_0_valid,portsAOI_filtered_0_valid} ;  
   reg [1:0] readys_mask ;  
   wire [1:0] _readys_filter_T_1=readys_valid&~readys_mask ;  
   wire [1:0] readys_readys=~({readys_mask[1],_readys_filter_T_1[1]|readys_mask[0]}&({_readys_filter_T_1[0],portsAOI_filtered_1_0_valid}|_readys_filter_T_1)) ;  
   wire winner_0=readys_readys[0]&portsAOI_filtered_0_valid ;  
   wire winner_1=readys_readys[1]&portsAOI_filtered_1_0_valid ;  
   wire _out_0_a_valid_T=portsAOI_filtered_0_valid|portsAOI_filtered_1_0_valid ;  
   reg state_0 ;  
   reg state_1 ;  
   wire muxState_0=idle ? winner_0:state_0 ;  
   wire muxState_1=idle ? winner_1:state_1 ;  
  assign allowed_0=idle ? readys_readys[0]:state_0; 
  assign allowed_1=idle ? readys_readys[1]:state_1; 
   wire out_0_a_valid=idle ? _out_0_a_valid_T:state_0&portsAOI_filtered_0_valid|state_1&portsAOI_filtered_1_0_valid ;  
   reg [8:0] beatsLeft_1 ;  
   wire idle_1=beatsLeft_1==9'h0 ;  
   wire [1:0] readys_valid_1={portsAOI_filtered_1_1_valid,portsAOI_filtered_1_valid} ;  
   reg [1:0] readys_mask_1 ;  
   wire [1:0] _readys_filter_T_3=readys_valid_1&~readys_mask_1 ;  
   wire [1:0] readys_readys_1=~({readys_mask_1[1],_readys_filter_T_3[1]|readys_mask_1[0]}&({_readys_filter_T_3[0],portsAOI_filtered_1_1_valid}|_readys_filter_T_3)) ;  
   wire winner_1_0=readys_readys_1[0]&portsAOI_filtered_1_valid ;  
   wire winner_1_1=readys_readys_1[1]&portsAOI_filtered_1_1_valid ;  
   wire _out_1_a_valid_T=portsAOI_filtered_1_valid|portsAOI_filtered_1_1_valid ;  
   reg state_1_0 ;  
   reg state_1_1 ;  
   wire muxState_1_0=idle_1 ? winner_1_0:state_1_0 ;  
   wire muxState_1_1=idle_1 ? winner_1_1:state_1_1 ;  
  assign allowed_1_0=idle_1 ? readys_readys_1[0]:state_1_0; 
  assign allowed_1_1=idle_1 ? readys_readys_1[1]:state_1_1; 
   wire out_1_a_valid=idle_1 ? _out_1_a_valid_T:state_1_0&portsAOI_filtered_1_valid|state_1_1&portsAOI_filtered_1_1_valid ;  
   reg [8:0] beatsLeft_2 ;  
   wire idle_2=beatsLeft_2==9'h0 ;  
   wire [1:0] readys_valid_2={portsAOI_filtered_1_2_valid,portsAOI_filtered_2_valid} ;  
   reg [1:0] readys_mask_2 ;  
   wire [1:0] _readys_filter_T_5=readys_valid_2&~readys_mask_2 ;  
   wire [1:0] readys_readys_2=~({readys_mask_2[1],_readys_filter_T_5[1]|readys_mask_2[0]}&({_readys_filter_T_5[0],portsAOI_filtered_1_2_valid}|_readys_filter_T_5)) ;  
   wire winner_2_0=readys_readys_2[0]&portsAOI_filtered_2_valid ;  
   wire winner_2_1=readys_readys_2[1]&portsAOI_filtered_1_2_valid ;  
   wire _out_2_a_valid_T=portsAOI_filtered_2_valid|portsAOI_filtered_1_2_valid ;  
   reg state_2_0 ;  
   reg state_2_1 ;  
   wire muxState_2_0=idle_2 ? winner_2_0:state_2_0 ;  
   wire muxState_2_1=idle_2 ? winner_2_1:state_2_1 ;  
  assign allowed_2_0=idle_2 ? readys_readys_2[0]:state_2_0; 
  assign allowed_2_1=idle_2 ? readys_readys_2[1]:state_2_1; 
   wire out_2_a_valid=idle_2 ? _out_2_a_valid_T:state_2_0&portsAOI_filtered_2_valid|state_2_1&portsAOI_filtered_1_2_valid ;  
   reg [8:0] beatsLeft_3 ;  
   wire idle_3=beatsLeft_3==9'h0 ;  
   wire [2:0] readys_valid_3={portsDIO_filtered_2_0_valid,portsDIO_filtered_1_0_valid,portsDIO_filtered_0_valid} ;  
   reg [2:0] readys_mask_3 ;  
   wire [2:0] _readys_filter_T_7=readys_valid_3&~readys_mask_3 ;  
   wire [3:0] _GEN={_readys_filter_T_7[1:0],portsDIO_filtered_2_0_valid,portsDIO_filtered_1_0_valid}|{_readys_filter_T_7,portsDIO_filtered_2_0_valid} ;  
   wire [2:0] readys_readys_3=~({readys_mask_3[2],_readys_filter_T_7[2]|readys_mask_3[1],_GEN[3]|readys_mask_3[0]}&(_GEN[2:0]|{_readys_filter_T_7[2],_GEN[3:2]})) ;  
   wire winner_3_0=readys_readys_3[0]&portsDIO_filtered_0_valid ;  
   wire winner_3_1=readys_readys_3[1]&portsDIO_filtered_1_0_valid ;  
   wire winner_3_2=readys_readys_3[2]&portsDIO_filtered_2_0_valid ;  
   wire _in_0_d_valid_T=portsDIO_filtered_0_valid|portsDIO_filtered_1_0_valid ;  
   reg state_3_0 ;  
   reg state_3_1 ;  
   reg state_3_2 ;  
   wire muxState_3_0=idle_3 ? winner_3_0:state_3_0 ;  
   wire muxState_3_1=idle_3 ? winner_3_1:state_3_1 ;  
   wire muxState_3_2=idle_3 ? winner_3_2:state_3_2 ;  
  assign allowed_3_0=idle_3 ? readys_readys_3[0]:state_3_0; 
  assign allowed_3_1=idle_3 ? readys_readys_3[1]:state_3_1; 
  assign allowed_3_2=idle_3 ? readys_readys_3[2]:state_3_2; 
   wire in_0_d_valid=idle_3 ? _in_0_d_valid_T|portsDIO_filtered_2_0_valid:state_3_0&portsDIO_filtered_0_valid|state_3_1&portsDIO_filtered_1_0_valid|state_3_2&portsDIO_filtered_2_0_valid ;  
   wire _in_0_d_bits_T_4=muxState_3_0&auto_out_0_d_bits_corrupt|muxState_3_1&auto_out_1_d_bits_corrupt|muxState_3_2&auto_out_2_d_bits_corrupt ;  
   wire _in_0_d_bits_T_14=muxState_3_0&auto_out_0_d_bits_denied|muxState_3_1&auto_out_1_d_bits_denied|muxState_3_2&auto_out_2_d_bits_denied ;  
   wire [1:0] _in_0_d_bits_T_18=(muxState_3_0 ? out_0_d_bits_sink:2'h0)|(muxState_3_1 ? auto_out_1_d_bits_sink:2'h0) ;  
   wire [3:0] _in_0_d_bits_T_24=(muxState_3_0 ? auto_out_0_d_bits_source[3:0]:4'h0)|(muxState_3_1 ? auto_out_1_d_bits_source[3:0]:4'h0)|(muxState_3_2 ? auto_out_2_d_bits_source[3:0]:4'h0) ;  
   wire [3:0] _in_0_d_bits_T_29=(muxState_3_0 ? auto_out_0_d_bits_size:4'h0)|(muxState_3_1 ? out_1_d_bits_size:4'h0)|(muxState_3_2 ? auto_out_2_d_bits_size:4'h0) ;  
   wire [1:0] _in_0_d_bits_T_33=(muxState_3_0 ? auto_out_0_d_bits_param:2'h0)|(muxState_3_1 ? auto_out_1_d_bits_param:2'h0) ;  
   wire [2:0] _in_0_d_bits_T_39=(muxState_3_0 ? auto_out_0_d_bits_opcode:3'h0)|(muxState_3_1 ? auto_out_1_d_bits_opcode:3'h0)|(muxState_3_2 ? auto_out_2_d_bits_opcode:3'h0) ;  
   reg [8:0] beatsLeft_4 ;  
   wire idle_4=beatsLeft_4==9'h0 ;  
   wire [2:0] readys_valid_4={portsDIO_filtered_2_1_valid,portsDIO_filtered_1_1_valid,portsDIO_filtered_1_valid} ;  
   reg [2:0] readys_mask_4 ;  
   wire [2:0] _readys_filter_T_9=readys_valid_4&~readys_mask_4 ;  
   wire [3:0] _GEN_0={_readys_filter_T_9[1:0],portsDIO_filtered_2_1_valid,portsDIO_filtered_1_1_valid}|{_readys_filter_T_9,portsDIO_filtered_2_1_valid} ;  
   wire [2:0] readys_readys_4=~({readys_mask_4[2],_readys_filter_T_9[2]|readys_mask_4[1],_GEN_0[3]|readys_mask_4[0]}&(_GEN_0[2:0]|{_readys_filter_T_9[2],_GEN_0[3:2]})) ;  
   wire winner_4_0=readys_readys_4[0]&portsDIO_filtered_1_valid ;  
   wire winner_4_1=readys_readys_4[1]&portsDIO_filtered_1_1_valid ;  
   wire winner_4_2=readys_readys_4[2]&portsDIO_filtered_2_1_valid ;  
   wire _in_1_d_valid_T=portsDIO_filtered_1_valid|portsDIO_filtered_1_1_valid ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~winner_0|~winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_out_0_a_valid_T|winner_0|winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
         if (~reset&~(~winner_1_0|~winner_1_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_out_1_a_valid_T|winner_1_0|winner_1_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
         if (~reset&~(~winner_2_0|~winner_2_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_out_2_a_valid_T|winner_2_0|winner_2_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
         if (~reset&~((~winner_3_0|~winner_3_1)&(~(winner_3_0|winner_3_1)|~winner_3_2)))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~(_in_0_d_valid_T|portsDIO_filtered_2_0_valid)|winner_3_0|winner_3_1|winner_3_2))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
         if (~reset&~((~winner_4_0|~winner_4_1)&(~(winner_4_0|winner_4_1)|~winner_4_2)))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~(_in_1_d_valid_T|portsDIO_filtered_2_1_valid)|winner_4_0|winner_4_1|winner_4_2))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg state_4_0 ;  
   reg state_4_1 ;  
   reg state_4_2 ;  
   wire muxState_4_0=idle_4 ? winner_4_0:state_4_0 ;  
   wire muxState_4_1=idle_4 ? winner_4_1:state_4_1 ;  
   wire muxState_4_2=idle_4 ? winner_4_2:state_4_2 ;  
  assign allowed_4_0=idle_4 ? readys_readys_4[0]:state_4_0; 
  assign allowed_4_1=idle_4 ? readys_readys_4[1]:state_4_1; 
  assign allowed_4_2=idle_4 ? readys_readys_4[2]:state_4_2; 
   wire in_1_d_valid=idle_4 ? _in_1_d_valid_T|portsDIO_filtered_2_1_valid:state_4_0&portsDIO_filtered_1_valid|state_4_1&portsDIO_filtered_1_1_valid|state_4_2&portsDIO_filtered_2_1_valid ;  
   wire _in_1_d_bits_T_4=muxState_4_0&auto_out_0_d_bits_corrupt|muxState_4_1&auto_out_1_d_bits_corrupt|muxState_4_2&auto_out_2_d_bits_corrupt ;  
   wire _in_1_d_bits_T_14=muxState_4_0&auto_out_0_d_bits_denied|muxState_4_1&auto_out_1_d_bits_denied|muxState_4_2&auto_out_2_d_bits_denied ;  
   wire [1:0] _in_1_d_bits_T_18=(muxState_4_0 ? out_0_d_bits_sink:2'h0)|(muxState_4_1 ? auto_out_1_d_bits_sink:2'h0) ;  
   wire [1:0] _in_1_d_bits_T_24=(muxState_4_0 ? auto_out_0_d_bits_source[1:0]:2'h0)|(muxState_4_1 ? auto_out_1_d_bits_source[1:0]:2'h0)|(muxState_4_2 ? auto_out_2_d_bits_source[1:0]:2'h0) ;  
   wire [3:0] _in_1_d_bits_T_29=(muxState_4_0 ? auto_out_0_d_bits_size:4'h0)|(muxState_4_1 ? out_1_d_bits_size:4'h0)|(muxState_4_2 ? auto_out_2_d_bits_size:4'h0) ;  
   wire [1:0] _in_1_d_bits_T_33=(muxState_4_0 ? auto_out_0_d_bits_param:2'h0)|(muxState_4_1 ? auto_out_1_d_bits_param:2'h0) ;  
   wire [2:0] _in_1_d_bits_T_39=(muxState_4_0 ? auto_out_0_d_bits_opcode:3'h0)|(muxState_4_1 ? auto_out_1_d_bits_opcode:3'h0)|(muxState_4_2 ? auto_out_2_d_bits_opcode:3'h0) ;  
   wire [1:0] _readys_mask_T=readys_readys&readys_valid ;  
   wire [1:0] _readys_mask_T_5=readys_readys_1&readys_valid_1 ;  
   wire [1:0] _readys_mask_T_10=readys_readys_2&readys_valid_2 ;  
   wire [2:0] _readys_mask_T_15=readys_readys_3&readys_valid_3 ;  
   wire [2:0] _readys_mask_T_18=_readys_mask_T_15|{_readys_mask_T_15[1:0],1'h0} ;  
   wire [2:0] _readys_mask_T_23=readys_readys_4&readys_valid_4 ;  
   wire [2:0] _readys_mask_T_26=_readys_mask_T_23|{_readys_mask_T_23[1:0],1'h0} ;  
   wire [26:0] _beatsAI_decode_T_1=27'hFFF<<auto_in_0_a_bits_size ;  
   wire [26:0] _beatsAI_decode_T_5=27'hFFF<<auto_in_1_a_bits_size ;  
   wire [26:0] _beatsDO_decode_T_1=27'hFFF<<auto_out_0_d_bits_size ;  
   wire [20:0] _beatsDO_decode_T_5=21'h3F<<auto_out_1_d_bits_size ;  
   wire [22:0] _beatsDO_decode_T_9=23'hFF<<auto_out_2_d_bits_size ;  
   wire latch=idle&auto_out_0_a_ready ;  
   wire latch_1=idle_1&auto_out_1_a_ready ;  
   wire latch_2=idle_2&auto_out_2_a_ready ;  
   wire latch_3=idle_3&auto_in_0_d_ready ;  
   wire latch_4=idle_4&auto_in_1_d_ready ;  
   wire [8:0] maskedBeats_0_3=winner_3_0&auto_out_0_d_bits_opcode[0] ? ~(_beatsDO_decode_T_1[11:3]):9'h0 ;  
   wire [8:0] maskedBeats_0_4=winner_4_0&auto_out_0_d_bits_opcode[0] ? ~(_beatsDO_decode_T_1[11:3]):9'h0 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              beatsLeft <=9'h0;
              readys_mask <=2'h3;
              state_0 <=1'h0;
              state_1 <=1'h0;
              beatsLeft_1 <=9'h0;
              readys_mask_1 <=2'h3;
              state_1_0 <=1'h0;
              state_1_1 <=1'h0;
              beatsLeft_2 <=9'h0;
              readys_mask_2 <=2'h3;
              state_2_0 <=1'h0;
              state_2_1 <=1'h0;
              beatsLeft_3 <=9'h0;
              readys_mask_3 <=3'h7;
              state_3_0 <=1'h0;
              state_3_1 <=1'h0;
              state_3_2 <=1'h0;
              beatsLeft_4 <=9'h0;
              readys_mask_4 <=3'h7;
              state_4_0 <=1'h0;
              state_4_1 <=1'h0;
              state_4_2 <=1'h0;
            end 
          else 
            begin 
              if (latch)
                 beatsLeft <=(winner_0&~(auto_in_0_a_bits_opcode[2]) ? ~(_beatsAI_decode_T_1[11:3]):9'h0)|(winner_1&~(auto_in_1_a_bits_opcode[2]) ? ~(_beatsAI_decode_T_5[11:3]):9'h0);
               else 
                 beatsLeft <=beatsLeft-{8'h0,auto_out_0_a_ready&out_0_a_valid};
              if (latch&(|readys_valid))
                 readys_mask <=_readys_mask_T|{_readys_mask_T[0],1'h0};
              if (idle)
                 begin 
                   state_0 <=winner_0;
                   state_1 <=winner_1;
                 end 
              if (latch_1)
                 beatsLeft_1 <=(winner_1_0&~(auto_in_0_a_bits_opcode[2]) ? ~(_beatsAI_decode_T_1[11:3]):9'h0)|(winner_1_1&~(auto_in_1_a_bits_opcode[2]) ? ~(_beatsAI_decode_T_5[11:3]):9'h0);
               else 
                 beatsLeft_1 <=beatsLeft_1-{8'h0,auto_out_1_a_ready&out_1_a_valid};
              if (latch_1&(|readys_valid_1))
                 readys_mask_1 <=_readys_mask_T_5|{_readys_mask_T_5[0],1'h0};
              if (idle_1)
                 begin 
                   state_1_0 <=winner_1_0;
                   state_1_1 <=winner_1_1;
                 end 
              if (latch_2)
                 beatsLeft_2 <=(winner_2_0&~(auto_in_0_a_bits_opcode[2]) ? ~(_beatsAI_decode_T_1[11:3]):9'h0)|(winner_2_1&~(auto_in_1_a_bits_opcode[2]) ? ~(_beatsAI_decode_T_5[11:3]):9'h0);
               else 
                 beatsLeft_2 <=beatsLeft_2-{8'h0,auto_out_2_a_ready&out_2_a_valid};
              if (latch_2&(|readys_valid_2))
                 readys_mask_2 <=_readys_mask_T_10|{_readys_mask_T_10[0],1'h0};
              if (idle_2)
                 begin 
                   state_2_0 <=winner_2_0;
                   state_2_1 <=winner_2_1;
                 end 
              if (latch_3)
                 beatsLeft_3 <={maskedBeats_0_3[8:5],{maskedBeats_0_3[4:3],maskedBeats_0_3[2:0]|(winner_3_1&auto_out_1_d_bits_opcode[0] ? ~(_beatsDO_decode_T_5[5:3]):3'h0)}|(winner_3_2&auto_out_2_d_bits_opcode[0] ? ~(_beatsDO_decode_T_9[7:3]):5'h0)};
               else 
                 beatsLeft_3 <=beatsLeft_3-{8'h0,auto_in_0_d_ready&in_0_d_valid};
              if (latch_3&(|readys_valid_3))
                 readys_mask_3 <=_readys_mask_T_18|{_readys_mask_T_18[0],2'h0};
              if (idle_3)
                 begin 
                   state_3_0 <=winner_3_0;
                   state_3_1 <=winner_3_1;
                   state_3_2 <=winner_3_2;
                 end 
              if (latch_4)
                 beatsLeft_4 <={maskedBeats_0_4[8:5],{maskedBeats_0_4[4:3],maskedBeats_0_4[2:0]|(winner_4_1&auto_out_1_d_bits_opcode[0] ? ~(_beatsDO_decode_T_5[5:3]):3'h0)}|(winner_4_2&auto_out_2_d_bits_opcode[0] ? ~(_beatsDO_decode_T_9[7:3]):5'h0)};
               else 
                 beatsLeft_4 <=beatsLeft_4-{8'h0,auto_in_1_d_ready&in_1_d_valid};
              if (latch_4&(|readys_valid_4))
                 readys_mask_4 <=_readys_mask_T_26|{_readys_mask_T_26[0],2'h0};
              if (idle_4)
                 begin 
                   state_4_0 <=winner_4_0;
                   state_4_1 <=winner_4_1;
                   state_4_2 <=winner_4_2;
                 end 
            end 
       end
  
  TLMonitor monitor(.clock(clock),.reset(reset),.io_in_a_ready(_portsAOI_in_0_a_ready_T_4),.io_in_a_valid(auto_in_0_a_valid),.io_in_a_bits_opcode(auto_in_0_a_bits_opcode),.io_in_a_bits_param(auto_in_0_a_bits_param),.io_in_a_bits_size(auto_in_0_a_bits_size),.io_in_a_bits_source(auto_in_0_a_bits_source),.io_in_a_bits_address(auto_in_0_a_bits_address),.io_in_a_bits_mask(auto_in_0_a_bits_mask),.io_in_a_bits_corrupt(auto_in_0_a_bits_corrupt),.io_in_d_ready(auto_in_0_d_ready),.io_in_d_valid(in_0_d_valid),.io_in_d_bits_opcode(_in_0_d_bits_T_39),.io_in_d_bits_param(_in_0_d_bits_T_33),.io_in_d_bits_size(_in_0_d_bits_T_29),.io_in_d_bits_source(_in_0_d_bits_T_24),.io_in_d_bits_sink(_in_0_d_bits_T_18),.io_in_d_bits_denied(_in_0_d_bits_T_14),.io_in_d_bits_corrupt(_in_0_d_bits_T_4)); 
  TLMonitor_1 monitor_1(.clock(clock),.reset(reset),.io_in_a_ready(_portsAOI_in_1_a_ready_T_4),.io_in_a_valid(auto_in_1_a_valid),.io_in_a_bits_opcode(auto_in_1_a_bits_opcode),.io_in_a_bits_param(auto_in_1_a_bits_param),.io_in_a_bits_size(auto_in_1_a_bits_size),.io_in_a_bits_source(auto_in_1_a_bits_source),.io_in_a_bits_address(auto_in_1_a_bits_address),.io_in_a_bits_mask(auto_in_1_a_bits_mask),.io_in_a_bits_corrupt(auto_in_1_a_bits_corrupt),.io_in_b_ready(auto_in_1_b_ready),.io_in_b_valid(auto_out_1_b_valid),.io_in_b_bits_param(auto_out_1_b_bits_param),.io_in_b_bits_address(auto_out_1_b_bits_address),.io_in_c_ready(auto_out_1_c_ready),.io_in_c_valid(auto_in_1_c_valid),.io_in_c_bits_opcode(auto_in_1_c_bits_opcode),.io_in_c_bits_param(auto_in_1_c_bits_param),.io_in_c_bits_size(auto_in_1_c_bits_size),.io_in_c_bits_source(auto_in_1_c_bits_source),.io_in_c_bits_address(auto_in_1_c_bits_address),.io_in_c_bits_corrupt(auto_in_1_c_bits_corrupt),.io_in_d_ready(auto_in_1_d_ready),.io_in_d_valid(in_1_d_valid),.io_in_d_bits_opcode(_in_1_d_bits_T_39),.io_in_d_bits_param(_in_1_d_bits_T_33),.io_in_d_bits_size(_in_1_d_bits_T_29),.io_in_d_bits_source(_in_1_d_bits_T_24),.io_in_d_bits_sink(_in_1_d_bits_T_18),.io_in_d_bits_denied(_in_1_d_bits_T_14),.io_in_d_bits_corrupt(_in_1_d_bits_T_4),.io_in_e_valid(auto_in_1_e_valid),.io_in_e_bits_sink(auto_in_1_e_bits_sink)); 
  assign auto_in_1_a_ready=_portsAOI_in_1_a_ready_T_4; 
  assign auto_in_1_b_valid=auto_out_1_b_valid; 
  assign auto_in_1_b_bits_param=auto_out_1_b_bits_param; 
  assign auto_in_1_b_bits_address=auto_out_1_b_bits_address; 
  assign auto_in_1_c_ready=auto_out_1_c_ready; 
  assign auto_in_1_d_valid=in_1_d_valid; 
  assign auto_in_1_d_bits_opcode=_in_1_d_bits_T_39; 
  assign auto_in_1_d_bits_param=_in_1_d_bits_T_33; 
  assign auto_in_1_d_bits_size=_in_1_d_bits_T_29; 
  assign auto_in_1_d_bits_source=_in_1_d_bits_T_24; 
  assign auto_in_1_d_bits_sink=_in_1_d_bits_T_18; 
  assign auto_in_1_d_bits_denied=_in_1_d_bits_T_14; 
  assign auto_in_1_d_bits_data=(muxState_4_0 ? auto_out_0_d_bits_data:64'h0)|(muxState_4_1 ? auto_out_1_d_bits_data:64'h0)|(muxState_4_2 ? auto_out_2_d_bits_data:64'h0); 
  assign auto_in_1_d_bits_corrupt=_in_1_d_bits_T_4; 
  assign auto_in_0_a_ready=_portsAOI_in_0_a_ready_T_4; 
  assign auto_in_0_d_valid=in_0_d_valid; 
  assign auto_in_0_d_bits_opcode=_in_0_d_bits_T_39; 
  assign auto_in_0_d_bits_param=_in_0_d_bits_T_33; 
  assign auto_in_0_d_bits_size=_in_0_d_bits_T_29; 
  assign auto_in_0_d_bits_source=_in_0_d_bits_T_24; 
  assign auto_in_0_d_bits_sink=_in_0_d_bits_T_18; 
  assign auto_in_0_d_bits_denied=_in_0_d_bits_T_14; 
  assign auto_in_0_d_bits_data=(muxState_3_0 ? auto_out_0_d_bits_data:64'h0)|(muxState_3_1 ? auto_out_1_d_bits_data:64'h0)|(muxState_3_2 ? auto_out_2_d_bits_data:64'h0); 
  assign auto_in_0_d_bits_corrupt=_in_0_d_bits_T_4; 
  assign auto_out_2_a_valid=out_2_a_valid; 
  assign auto_out_2_a_bits_opcode=(muxState_2_0 ? auto_in_0_a_bits_opcode:3'h0)|(muxState_2_1 ? auto_in_1_a_bits_opcode:3'h0); 
  assign auto_out_2_a_bits_param=(muxState_2_0 ? auto_in_0_a_bits_param:3'h0)|(muxState_2_1 ? auto_in_1_a_bits_param:3'h0); 
  assign auto_out_2_a_bits_size=(muxState_2_0 ? auto_in_0_a_bits_size:4'h0)|(muxState_2_1 ? auto_in_1_a_bits_size:4'h0); 
  assign auto_out_2_a_bits_source=(muxState_2_0 ? in_0_a_bits_source:5'h0)|(muxState_2_1 ? in_1_a_bits_source:5'h0); 
  assign auto_out_2_a_bits_address=(muxState_2_0 ? auto_in_0_a_bits_address[30:0]:31'h0)|(muxState_2_1 ? auto_in_1_a_bits_address[30:0]:31'h0); 
  assign auto_out_2_a_bits_mask=(muxState_2_0 ? auto_in_0_a_bits_mask:8'h0)|(muxState_2_1 ? auto_in_1_a_bits_mask:8'h0); 
  assign auto_out_2_a_bits_data=(muxState_2_0 ? auto_in_0_a_bits_data:64'h0)|(muxState_2_1 ? auto_in_1_a_bits_data:64'h0); 
  assign auto_out_2_a_bits_corrupt=muxState_2_0&auto_in_0_a_bits_corrupt|muxState_2_1&auto_in_1_a_bits_corrupt; 
  assign auto_out_2_d_ready=~(auto_out_2_d_bits_source[4])&auto_in_0_d_ready&allowed_3_2|requestDOI_2_1&auto_in_1_d_ready&allowed_4_2; 
  assign auto_out_1_a_valid=out_1_a_valid; 
  assign auto_out_1_a_bits_opcode=(muxState_1_0 ? auto_in_0_a_bits_opcode:3'h0)|(muxState_1_1 ? auto_in_1_a_bits_opcode:3'h0); 
  assign auto_out_1_a_bits_param=(muxState_1_0 ? auto_in_0_a_bits_param:3'h0)|(muxState_1_1 ? auto_in_1_a_bits_param:3'h0); 
  assign auto_out_1_a_bits_size=(muxState_1_0 ? auto_in_0_a_bits_size[2:0]:3'h0)|(muxState_1_1 ? auto_in_1_a_bits_size[2:0]:3'h0); 
  assign auto_out_1_a_bits_source=(muxState_1_0 ? in_0_a_bits_source:5'h0)|(muxState_1_1 ? in_1_a_bits_source:5'h0); 
  assign auto_out_1_a_bits_address=(muxState_1_0 ? auto_in_0_a_bits_address:32'h0)|(muxState_1_1 ? auto_in_1_a_bits_address:32'h0); 
  assign auto_out_1_a_bits_mask=(muxState_1_0 ? auto_in_0_a_bits_mask:8'h0)|(muxState_1_1 ? auto_in_1_a_bits_mask:8'h0); 
  assign auto_out_1_a_bits_data=(muxState_1_0 ? auto_in_0_a_bits_data:64'h0)|(muxState_1_1 ? auto_in_1_a_bits_data:64'h0); 
  assign auto_out_1_a_bits_corrupt=muxState_1_0&auto_in_0_a_bits_corrupt|muxState_1_1&auto_in_1_a_bits_corrupt; 
  assign auto_out_1_b_ready=auto_in_1_b_ready; 
  assign auto_out_1_c_valid=auto_in_1_c_valid; 
  assign auto_out_1_c_bits_opcode=auto_in_1_c_bits_opcode; 
  assign auto_out_1_c_bits_param=auto_in_1_c_bits_param; 
  assign auto_out_1_c_bits_size=auto_in_1_c_bits_size[2:0]; 
  assign auto_out_1_c_bits_source={3'h4,auto_in_1_c_bits_source}; 
  assign auto_out_1_c_bits_address=auto_in_1_c_bits_address; 
  assign auto_out_1_c_bits_data=auto_in_1_c_bits_data; 
  assign auto_out_1_c_bits_corrupt=auto_in_1_c_bits_corrupt; 
  assign auto_out_1_d_ready=~(auto_out_1_d_bits_source[4])&auto_in_0_d_ready&allowed_3_1|requestDOI_1_1&auto_in_1_d_ready&allowed_4_1; 
  assign auto_out_1_e_valid=auto_in_1_e_valid; 
  assign auto_out_1_e_bits_sink=auto_in_1_e_bits_sink; 
  assign auto_out_0_a_valid=out_0_a_valid; 
  assign auto_out_0_a_bits_opcode=(muxState_0 ? auto_in_0_a_bits_opcode:3'h0)|(muxState_1 ? auto_in_1_a_bits_opcode:3'h0); 
  assign auto_out_0_a_bits_param=(muxState_0 ? auto_in_0_a_bits_param:3'h0)|(muxState_1 ? auto_in_1_a_bits_param:3'h0); 
  assign auto_out_0_a_bits_size=(muxState_0 ? auto_in_0_a_bits_size:4'h0)|(muxState_1 ? auto_in_1_a_bits_size:4'h0); 
  assign auto_out_0_a_bits_source=(muxState_0 ? in_0_a_bits_source:5'h0)|(muxState_1 ? in_1_a_bits_source:5'h0); 
  assign auto_out_0_a_bits_address=(muxState_0 ? auto_in_0_a_bits_address[27:0]:28'h0)|(muxState_1 ? auto_in_1_a_bits_address[27:0]:28'h0); 
  assign auto_out_0_a_bits_mask=(muxState_0 ? auto_in_0_a_bits_mask:8'h0)|(muxState_1 ? auto_in_1_a_bits_mask:8'h0); 
  assign auto_out_0_a_bits_data=(muxState_0 ? auto_in_0_a_bits_data:64'h0)|(muxState_1 ? auto_in_1_a_bits_data:64'h0); 
  assign auto_out_0_a_bits_corrupt=muxState_0&auto_in_0_a_bits_corrupt|muxState_1&auto_in_1_a_bits_corrupt; 
  assign auto_out_0_d_ready=~(auto_out_0_d_bits_source[4])&auto_in_0_d_ready&allowed_3_0|requestDOI_0_1&auto_in_1_d_ready&allowed_4_0; 
endmodule
 
module TLMonitor_2 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [3:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [3:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [3:0] source ;  
   reg [31:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [3:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [15:0] inflight ;  
   reg [63:0] inflight_opcodes ;  
   reg [127:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [63:0] _a_opcode_lookup_T_1=inflight_opcodes>>{58'h0,io_in_d_bits_source,2'h0} ;  
   wire [15:0] _GEN_0={12'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [15:0] _GEN_2={12'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [15:0] inflight_1 ;  
   reg [127:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_bits_size<4'h7 ;  
   wire _GEN_6=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_7=_GEN_4&_GEN_5&_GEN_6 ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_9=io_in_a_bits_param>3'h2 ;  
   wire _GEN_10=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_11=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_13={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_14=_GEN_4&_GEN_13 ;  
   wire _GEN_15=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_16={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_17={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_18={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_19=io_in_a_bits_mask!=mask ;  
   wire _GEN_20=_GEN_4&(_GEN_14|_GEN_5&(_GEN_15|_GEN_16|_GEN_17|_GEN_6)|io_in_a_bits_size<4'h9&_GEN_18) ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_22=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_23=_GEN_4&io_in_a_bits_size<4'h4&(_GEN_15|_GEN_13|_GEN_16|_GEN_17) ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_26=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_27=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_28=io_in_d_bits_size<4'h3 ;  
   wire _GEN_29=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_30=io_in_d_bits_param==2'h2 ;  
   wire _GEN_31=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_32=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_33=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_35=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_36=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_37=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [127:0] _GEN_38={121'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [15:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 16'h1<<_GEN_0:16'h0 ;  
   wire _GEN_39=io_in_d_valid&d_first_1 ;  
   wire _GEN_40=_GEN_39&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_41=_GEN_40&same_cycle_resp&~reset ;  
   wire _GEN_42=_GEN_40&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_43={4'h0,io_in_d_bits_size} ;  
   wire _GEN_44=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [15:0] _GEN_45=inflight>>_GEN_0 ;  
   wire [15:0] _GEN_46=inflight>>_GEN_2 ;  
   wire [127:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_38 ;  
   wire [15:0] _GEN_47=inflight_1>>_GEN_2 ;  
   wire [127:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_38 ;  
  always @( posedge clock)
       begin 
         if (_GEN_8&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~(_GEN_14|_GEN_5&(_GEN_15|{io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0|_GEN_16|_GEN_17|_GEN_18|_GEN_6)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(_GEN_4&_GEN_14))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_45[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~reset&~(_GEN_46[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_43!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_40 ? 16'h1<<_GEN_2:16'h0)|a_set_wo_ready==16'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==16'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~(_GEN_47[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&_GEN_43!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==16'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_48={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_48 ;  
   wire [142:0] _GEN_49={136'h0,io_in_d_bits_source,3'h0} ;  
   wire [142:0] _d_opcodes_clr_T_5=143'hF<<{137'h0,io_in_d_bits_source,2'h0} ;  
   wire [130:0] _a_opcodes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{125'h0,io_in_a_bits_source,2'h0} ;  
   wire [142:0] _d_sizes_clr_T_5=143'hFF<<_GEN_49 ;  
   wire [131:0] _a_sizes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{125'h0,io_in_a_bits_source,3'h0} ;  
   wire [142:0] _d_sizes_clr_T_11=143'hFF<<_GEN_49 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_50=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_51=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=16'h0;
              inflight_opcodes <=64'h0;
              inflight_sizes <=128'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=16'h0;
              inflight_sizes_1 <=128'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? 16'h1<<_GEN_0:16'h0))&~(_GEN_50 ? 16'h1<<_GEN_2:16'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[63:0]:64'h0))&~(_GEN_50 ? _d_opcodes_clr_T_5[63:0]:64'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[127:0]:128'h0))&~(_GEN_50 ? _d_sizes_clr_T_5[127:0]:128'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_51 ? 16'h1<<_GEN_2:16'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_51 ? _d_sizes_clr_T_11[127:0]:128'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLMonitor_3 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [1:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_b_ready,
  input io_in_b_valid,
  input [1:0] io_in_b_bits_param,
  input [31:0] io_in_b_bits_address,
  input io_in_c_ready,
  input io_in_c_valid,
  input [2:0] io_in_c_bits_opcode,
  input [2:0] io_in_c_bits_param,
  input [3:0] io_in_c_bits_size,
  input [1:0] io_in_c_bits_source,
  input [31:0] io_in_c_bits_address,
  input io_in_c_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [1:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt,
  input io_in_e_valid,
  input [1:0] io_in_e_bits_sink) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire [26:0] _GEN_0={23'h0,io_in_c_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [1:0] source ;  
   reg [31:0] address ;  
   wire _d_first_T_3=io_in_d_ready&io_in_d_valid ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [1:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [8:0] b_first_counter ;  
   reg [1:0] param_2 ;  
   reg [31:0] address_1 ;  
   wire _c_first_T_1=io_in_c_ready&io_in_c_valid ;  
   reg [8:0] c_first_counter ;  
   reg [2:0] opcode_3 ;  
   reg [2:0] param_3 ;  
   reg [3:0] size_3 ;  
   reg [1:0] source_3 ;  
   reg [31:0] address_2 ;  
   reg [2:0] inflight ;  
   reg [11:0] inflight_opcodes ;  
   reg [23:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [11:0] _a_opcode_lookup_T_1=inflight_opcodes>>{8'h0,io_in_d_bits_source,2'h0} ;  
   wire [3:0] _GEN_1={2'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [3:0] _GEN_3={2'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [2:0] inflight_1 ;  
   reg [23:0] inflight_sizes_1 ;  
   reg [8:0] c_first_counter_1 ;  
   wire c_first_1=c_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   wire _GEN_4=io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1] ;  
   wire [3:0] _GEN_5={2'h0,io_in_c_bits_source} ;  
   wire _GEN_6=_c_first_T_1&c_first_1&_GEN_4 ;  
   reg [31:0] watchdog_1 ;  
   reg [3:0] inflight_2 ;  
   reg [8:0] d_first_counter_3 ;  
   wire d_first_3=d_first_counter_3==9'h0 ;  
   wire _GEN_7=_d_first_T_3&d_first_3&io_in_d_bits_opcode[2]&~(io_in_d_bits_opcode[1]) ;  
   wire [3:0] _GEN_8={2'h0,io_in_d_bits_sink} ;  
   wire [3:0] d_set=_GEN_7 ? 4'h1<<_GEN_8:4'h0 ;  
   wire [3:0] _GEN_9={2'h0,io_in_e_bits_sink} ;  
   wire _source_ok_T=io_in_a_bits_source==2'h0 ;  
   wire _source_ok_T_1=io_in_a_bits_source==2'h1 ;  
   wire _source_ok_T_2=io_in_a_bits_source==2'h2 ;  
   wire source_ok=_source_ok_T|_source_ok_T_1|_source_ok_T_2 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_10=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_11=io_in_a_bits_size<4'hD ;  
   wire _GEN_12=_GEN_11&(_source_ok_T|_source_ok_T_1|_source_ok_T_2) ;  
   wire _GEN_13=io_in_a_bits_size<4'h7 ;  
   wire _GEN_14=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_15=_GEN_12&_GEN_13&_GEN_14 ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_17=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_18={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_19={io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0 ;  
   wire _GEN_20={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_21={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_22={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_23=_GEN_17|_GEN_18 ;  
   wire _GEN_24=_source_ok_T&io_in_a_bits_size==4'h6&_GEN_11&(_GEN_23|_GEN_19|_GEN_20|_GEN_21|_GEN_22|_GEN_14) ;  
   wire _GEN_25=io_in_a_bits_param>3'h2 ;  
   wire _GEN_26=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_27=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_28=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_29=_GEN_11&_GEN_18 ;  
   wire _GEN_30=io_in_a_bits_mask!=mask ;  
   wire _GEN_31=_GEN_12&(_GEN_29|_GEN_13&(_GEN_17|_GEN_20|_GEN_21|_GEN_14)|io_in_a_bits_size<4'h9&_GEN_22) ;  
   wire _GEN_32=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_33=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_34=_GEN_12&io_in_a_bits_size<4'h4&(_GEN_23|_GEN_20|_GEN_21) ;  
   wire _GEN_35=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_36=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_37=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source==2'h0|io_in_d_bits_source==2'h1|io_in_d_bits_source==2'h2 ;  
   wire _GEN_38=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_39=io_in_d_bits_size<4'h3 ;  
   wire _GEN_40=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_41=io_in_d_bits_param==2'h2 ;  
   wire _GEN_42=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_43=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_44=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_45=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_46=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire [19:0] _GEN_47={io_in_b_bits_address[31:14],~(io_in_b_bits_address[13:12])} ;  
   wire [5:0] _GEN_48={io_in_b_bits_address[31:28],~(io_in_b_bits_address[27:26])} ;  
   wire [15:0] _GEN_49={io_in_b_bits_address[31:26],io_in_b_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_50={io_in_b_bits_address[31:17],~(io_in_b_bits_address[16])} ;  
   wire _GEN_51=io_in_b_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_52={io_in_b_bits_address[31],~(io_in_b_bits_address[30:29])} ;  
   wire _GEN_53=io_in_b_valid&~reset ;  
   wire _source_ok_T_8=io_in_c_bits_source==2'h0 ;  
   wire _source_ok_T_9=io_in_c_bits_source==2'h1 ;  
   wire _source_ok_T_10=io_in_c_bits_source==2'h2 ;  
   wire source_ok_2=_source_ok_T_8|_source_ok_T_9|_source_ok_T_10 ;  
   wire [26:0] _is_aligned_mask_T_7=27'hFFF<<_GEN_0 ;  
   wire [11:0] _GEN_54=io_in_c_bits_address[11:0]&~(_is_aligned_mask_T_7[11:0]) ;  
   wire [19:0] _GEN_55={io_in_c_bits_address[31:14],~(io_in_c_bits_address[13:12])} ;  
   wire [5:0] _GEN_56={io_in_c_bits_address[31:28],~(io_in_c_bits_address[27:26])} ;  
   wire [15:0] _GEN_57={io_in_c_bits_address[31:26],io_in_c_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_58={io_in_c_bits_address[31:17],~(io_in_c_bits_address[16])} ;  
   wire _GEN_59=io_in_c_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_60={io_in_c_bits_address[31],~(io_in_c_bits_address[30:29])} ;  
   wire address_ok_1=~(|_GEN_55)|~(|_GEN_56)|~(|_GEN_57)|~(|(io_in_c_bits_address[31:12]))|~(|_GEN_58)|~_GEN_59|~(|_GEN_60) ;  
   wire _GEN_61=io_in_c_valid&io_in_c_bits_opcode==3'h4&~reset ;  
   wire _GEN_62=io_in_c_bits_size<4'h3 ;  
   wire _GEN_63=io_in_c_valid&io_in_c_bits_opcode==3'h5&~reset ;  
   wire _GEN_64=io_in_c_bits_size<4'hD ;  
   wire _GEN_65=_GEN_64&(_source_ok_T_8|_source_ok_T_9|_source_ok_T_10)&io_in_c_bits_size<4'h7&~_GEN_59 ;  
   wire _GEN_66=io_in_c_valid&io_in_c_bits_opcode==3'h6&~reset ;  
   wire _GEN_67=_source_ok_T_8&io_in_c_bits_size==4'h6&_GEN_64&(~(|(io_in_c_bits_address[31:12]))|~(|_GEN_55)|~(|_GEN_58)|~(|_GEN_57)|~(|_GEN_56)|~(|_GEN_60)|~_GEN_59) ;  
   wire _GEN_68=io_in_c_valid&(&io_in_c_bits_opcode)&~reset ;  
   wire _GEN_69=io_in_c_valid&io_in_c_bits_opcode==3'h0&~reset ;  
   wire _GEN_70=io_in_c_valid&io_in_c_bits_opcode==3'h1&~reset ;  
   wire _GEN_71=io_in_c_valid&io_in_c_bits_opcode==3'h2&~reset ;  
   wire _GEN_72=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_73=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_74=io_in_b_valid&(|b_first_counter)&~reset ;  
   wire _GEN_75=io_in_c_valid&(|c_first_counter)&~reset ;  
   wire [23:0] _GEN_76={19'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [3:0] _a_set_wo_ready_T=4'h1<<_GEN_1 ;  
   wire [2:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[2:0]:3'h0 ;  
   wire _GEN_77=io_in_d_valid&d_first_1 ;  
   wire _GEN_78=_GEN_77&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [2:0] _GEN_79={1'h0,io_in_d_bits_source} ;  
   wire _GEN_80=_GEN_78&same_cycle_resp&~reset ;  
   wire _GEN_81=_GEN_78&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_82={4'h0,io_in_d_bits_size} ;  
   wire _same_cycle_resp_T_3=io_in_c_valid&c_first_1 ;  
   wire [3:0] _c_set_wo_ready_T=4'h1<<_GEN_5 ;  
   wire [2:0] c_set_wo_ready=_same_cycle_resp_T_3&_GEN_4 ? _c_set_wo_ready_T[2:0]:3'h0 ;  
   wire _GEN_83=io_in_d_valid&d_first_2 ;  
   wire _GEN_84=_GEN_83&d_release_ack ;  
   wire same_cycle_resp_1=_same_cycle_resp_T_3&io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1]&io_in_c_bits_source==io_in_d_bits_source ;  
   wire [2:0] _GEN_85=inflight>>io_in_a_bits_source ;  
   wire [2:0] _GEN_86=inflight>>_GEN_79 ;  
   wire [23:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_76 ;  
   wire [3:0] _d_clr_wo_ready_T=4'h1<<_GEN_3 ;  
   wire [2:0] _GEN_87=inflight_1>>io_in_c_bits_source ;  
   wire [2:0] _GEN_88=inflight_1>>_GEN_79 ;  
   wire [23:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_76 ;  
   wire [3:0] _d_clr_wo_ready_T_1=4'h1<<_GEN_3 ;  
   wire [3:0] _GEN_89=inflight_2>>_GEN_8 ;  
   wire [3:0] _GEN_90=(d_set|inflight_2)>>_GEN_9 ;  
  always @( posedge clock)
       begin 
         if (_GEN_16&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(_GEN_29|_GEN_13&(_GEN_17|_GEN_19|_GEN_20|_GEN_21|_GEN_22|_GEN_14)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~_GEN_34)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~_GEN_34)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~(_GEN_12&_GEN_29))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|_GEN_10))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&~(~(|(io_in_b_bits_address[31:12]))|~(|_GEN_47)|~(|_GEN_50)|~(|_GEN_49)|~(|_GEN_48)|~(|_GEN_52)|~_GEN_51))
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&~(~(|_GEN_47)|~(|_GEN_48)|~(|_GEN_49)|~(|(io_in_b_bits_address[31:12]))|~(|_GEN_50)|~_GEN_51|~(|_GEN_52)))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&(|(io_in_b_bits_address[5:0])))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&(&io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&~_GEN_65)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&~_GEN_67)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_66&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&~_GEN_65)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&~_GEN_67)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_68&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_70&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid param (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck is corrupt (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_72&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&io_in_b_bits_param!=param_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&io_in_b_bits_address!=address_1)
            begin 
              if (1)$display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_opcode!=opcode_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_param!=param_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel param changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_size!=size_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel size changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_source!=source_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel source changed within multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_75&io_in_c_bits_address!=address_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel address changed with multibeat operation (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_85[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&~reset&~(_GEN_86[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&_GEN_82!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_77&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_78 ? _d_clr_wo_ready_T[2:0]:3'h0)|a_set_wo_ready==3'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==3'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~reset&_GEN_87[0])
            begin 
              if (1)$display("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&~reset&~(_GEN_88[0]|same_cycle_resp_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&same_cycle_resp_1&~reset&io_in_d_bits_size!=io_in_c_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&~same_cycle_resp_1&~reset&_GEN_82!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&c_first_1&io_in_c_valid&io_in_c_bits_source==io_in_d_bits_source&d_release_ack&~(io_in_c_bits_opcode==3'h4|io_in_c_bits_opcode==3'h5)&~reset&~(~io_in_d_ready|io_in_c_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if ((|c_set_wo_ready)&~reset&c_set_wo_ready==(_GEN_84 ? _d_clr_wo_ready_T_1[2:0]:3'h0))
            begin 
              if (1)$display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==3'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~reset&_GEN_89[0])
            begin 
              if (1)$display("Assertion failed: 'D' channel re-used a sink ID (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_e_valid&~reset&~(_GEN_90[0]))
            begin 
              if (1)$display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/SystemBus.scala:41:96)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_91={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_91 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_91 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_91 ;  
   wire [26:0] _d_first_beats1_decode_T_13=27'hFFF<<_GEN_91 ;  
   wire [26:0] _c_first_beats1_decode_T_1=27'hFFF<<_GEN_0 ;  
   wire [26:0] _c_first_beats1_decode_T_5=27'hFFF<<_GEN_0 ;  
   wire _GEN_92=_d_first_T_3&d_first_1&~d_release_ack ;  
   wire [46:0] _GEN_93={42'h0,io_in_d_bits_source,3'h0} ;  
   wire _GEN_94=_d_first_T_3&d_first_2&d_release_ack ;  
   wire [3:0] _d_clr_T=4'h1<<_GEN_3 ;  
   wire [3:0] _a_set_T=4'h1<<_GEN_1 ;  
   wire [46:0] _d_opcodes_clr_T_5=47'hF<<{43'h0,io_in_d_bits_source,2'h0} ;  
   wire [34:0] _a_opcodes_set_T_1={31'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{31'h0,io_in_a_bits_source,2'h0} ;  
   wire [46:0] _d_sizes_clr_T_5=47'hFF<<_GEN_93 ;  
   wire [35:0] _a_sizes_set_T_1={31'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:5'h0}<<{31'h0,io_in_a_bits_source,3'h0} ;  
   wire [3:0] _d_clr_T_1=4'h1<<_GEN_3 ;  
   wire [3:0] _c_set_T=4'h1<<_GEN_5 ;  
   wire [46:0] _d_sizes_clr_T_11=47'hFF<<_GEN_93 ;  
   wire [35:0] _c_sizes_set_T_1={31'h0,_GEN_6 ? {io_in_c_bits_size,1'h1}:5'h0}<<{31'h0,io_in_c_bits_source,3'h0} ;  
   wire b_first_done=io_in_b_ready&io_in_b_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              b_first_counter <=9'h0;
              c_first_counter <=9'h0;
              inflight <=3'h0;
              inflight_opcodes <=12'h0;
              inflight_sizes <=24'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=3'h0;
              inflight_sizes_1 <=24'h0;
              c_first_counter_1 <=9'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
              inflight_2 <=4'h0;
              d_first_counter_3 <=9'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_3)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   if (d_first_3)
                      d_first_counter_3 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_13[11:3]):9'h0;
                    else 
                      d_first_counter_3 <=d_first_counter_3-9'h1;
                 end 
              if (b_first_done)
                 begin 
                   if (|b_first_counter)
                      b_first_counter <=b_first_counter-9'h1;
                    else 
                      b_first_counter <=9'h0;
                 end 
              if (_c_first_T_1)
                 begin 
                   if (|c_first_counter)
                      c_first_counter <=c_first_counter-9'h1;
                    else 
                      c_first_counter <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_1[11:3]):9'h0;
                   if (c_first_1)
                      c_first_counter_1 <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      c_first_counter_1 <=c_first_counter_1-9'h1;
                 end 
              inflight <=(inflight|(_GEN_2 ? _a_set_T[2:0]:3'h0))&~(_GEN_92 ? _d_clr_T[2:0]:3'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[11:0]:12'h0))&~(_GEN_92 ? _d_opcodes_clr_T_5[11:0]:12'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[23:0]:24'h0))&~(_GEN_92 ? _d_sizes_clr_T_5[23:0]:24'h0);
              if (_a_first_T_1|_d_first_T_3)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=(inflight_1|(_GEN_6 ? _c_set_T[2:0]:3'h0))&~(_GEN_94 ? _d_clr_T_1[2:0]:3'h0);
              inflight_sizes_1 <=(inflight_sizes_1|(_GEN_6 ? _c_sizes_set_T_1[23:0]:24'h0))&~(_GEN_94 ? _d_sizes_clr_T_11[23:0]:24'h0);
              if (_c_first_T_1|_d_first_T_3)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight_2 <=(inflight_2|d_set)&~(io_in_e_valid ? 4'h1<<_GEN_9:4'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_3&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
         if (b_first_done&~(|b_first_counter))
            begin 
              param_2 <=io_in_b_bits_param;
              address_1 <=io_in_b_bits_address;
            end 
         if (_c_first_T_1&~(|c_first_counter))
            begin 
              opcode_3 <=io_in_c_bits_opcode;
              param_3 <=io_in_c_bits_param;
              size_3 <=io_in_c_bits_size;
              source_3 <=io_in_c_bits_source;
              address_2 <=io_in_c_bits_address;
            end 
       end
  
endmodule
 
module TLFIFOFixer (
  input clock,
  input reset,
  output auto_in_1_a_ready,
  input auto_in_1_a_valid,
  input [2:0] auto_in_1_a_bits_opcode,
  input [2:0] auto_in_1_a_bits_param,
  input [3:0] auto_in_1_a_bits_size,
  input [1:0] auto_in_1_a_bits_source,
  input [31:0] auto_in_1_a_bits_address,
  input [7:0] auto_in_1_a_bits_mask,
  input [63:0] auto_in_1_a_bits_data,
  input auto_in_1_a_bits_corrupt,
  input auto_in_1_b_ready,
  output auto_in_1_b_valid,
  output [1:0] auto_in_1_b_bits_param,
  output [31:0] auto_in_1_b_bits_address,
  output auto_in_1_c_ready,
  input auto_in_1_c_valid,
  input [2:0] auto_in_1_c_bits_opcode,
  input [2:0] auto_in_1_c_bits_param,
  input [3:0] auto_in_1_c_bits_size,
  input [1:0] auto_in_1_c_bits_source,
  input [31:0] auto_in_1_c_bits_address,
  input [63:0] auto_in_1_c_bits_data,
  input auto_in_1_c_bits_corrupt,
  input auto_in_1_d_ready,
  output auto_in_1_d_valid,
  output [2:0] auto_in_1_d_bits_opcode,
  output [1:0] auto_in_1_d_bits_param,
  output [3:0] auto_in_1_d_bits_size,
  output [1:0] auto_in_1_d_bits_source,
  output [1:0] auto_in_1_d_bits_sink,
  output auto_in_1_d_bits_denied,
  output [63:0] auto_in_1_d_bits_data,
  output auto_in_1_d_bits_corrupt,
  input auto_in_1_e_valid,
  input [1:0] auto_in_1_e_bits_sink,
  output auto_in_0_a_ready,
  input auto_in_0_a_valid,
  input [2:0] auto_in_0_a_bits_opcode,
  input [2:0] auto_in_0_a_bits_param,
  input [3:0] auto_in_0_a_bits_size,
  input [3:0] auto_in_0_a_bits_source,
  input [31:0] auto_in_0_a_bits_address,
  input [7:0] auto_in_0_a_bits_mask,
  input [63:0] auto_in_0_a_bits_data,
  input auto_in_0_a_bits_corrupt,
  input auto_in_0_d_ready,
  output auto_in_0_d_valid,
  output [2:0] auto_in_0_d_bits_opcode,
  output [1:0] auto_in_0_d_bits_param,
  output [3:0] auto_in_0_d_bits_size,
  output [3:0] auto_in_0_d_bits_source,
  output [1:0] auto_in_0_d_bits_sink,
  output auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output auto_in_0_d_bits_corrupt,
  input auto_out_1_a_ready,
  output auto_out_1_a_valid,
  output [2:0] auto_out_1_a_bits_opcode,
  output [2:0] auto_out_1_a_bits_param,
  output [3:0] auto_out_1_a_bits_size,
  output [1:0] auto_out_1_a_bits_source,
  output [31:0] auto_out_1_a_bits_address,
  output [7:0] auto_out_1_a_bits_mask,
  output [63:0] auto_out_1_a_bits_data,
  output auto_out_1_a_bits_corrupt,
  output auto_out_1_b_ready,
  input auto_out_1_b_valid,
  input [1:0] auto_out_1_b_bits_param,
  input [31:0] auto_out_1_b_bits_address,
  input auto_out_1_c_ready,
  output auto_out_1_c_valid,
  output [2:0] auto_out_1_c_bits_opcode,
  output [2:0] auto_out_1_c_bits_param,
  output [3:0] auto_out_1_c_bits_size,
  output [1:0] auto_out_1_c_bits_source,
  output [31:0] auto_out_1_c_bits_address,
  output [63:0] auto_out_1_c_bits_data,
  output auto_out_1_c_bits_corrupt,
  output auto_out_1_d_ready,
  input auto_out_1_d_valid,
  input [2:0] auto_out_1_d_bits_opcode,
  input [1:0] auto_out_1_d_bits_param,
  input [3:0] auto_out_1_d_bits_size,
  input [1:0] auto_out_1_d_bits_source,
  input [1:0] auto_out_1_d_bits_sink,
  input auto_out_1_d_bits_denied,
  input [63:0] auto_out_1_d_bits_data,
  input auto_out_1_d_bits_corrupt,
  output auto_out_1_e_valid,
  output [1:0] auto_out_1_e_bits_sink,
  input auto_out_0_a_ready,
  output auto_out_0_a_valid,
  output [2:0] auto_out_0_a_bits_opcode,
  output [2:0] auto_out_0_a_bits_param,
  output [3:0] auto_out_0_a_bits_size,
  output [3:0] auto_out_0_a_bits_source,
  output [31:0] auto_out_0_a_bits_address,
  output [7:0] auto_out_0_a_bits_mask,
  output [63:0] auto_out_0_a_bits_data,
  output auto_out_0_a_bits_corrupt,
  output auto_out_0_d_ready,
  input auto_out_0_d_valid,
  input [2:0] auto_out_0_d_bits_opcode,
  input [1:0] auto_out_0_d_bits_param,
  input [3:0] auto_out_0_d_bits_size,
  input [3:0] auto_out_0_d_bits_source,
  input [1:0] auto_out_0_d_bits_sink,
  input auto_out_0_d_bits_denied,
  input [63:0] auto_out_0_d_bits_data,
  input auto_out_0_d_bits_corrupt) ; 
   wire [1:0] a_id={auto_in_0_a_bits_address[30],~(auto_in_0_a_bits_address[30])} ;  
   wire a_noDomain=a_id==2'h0 ;  
   reg [8:0] a_first_counter ;  
   wire a_first=a_first_counter==9'h0 ;  
   reg [8:0] d_first_counter ;  
   reg flight_0 ;  
   reg flight_1 ;  
   reg flight_2 ;  
   reg flight_3 ;  
   reg flight_4 ;  
   reg flight_5 ;  
   reg flight_6 ;  
   reg flight_7 ;  
   reg flight_8 ;  
   reg flight_9 ;  
   reg flight_10 ;  
   reg flight_11 ;  
   reg flight_12 ;  
   reg flight_13 ;  
   reg flight_14 ;  
   reg flight_15 ;  
   reg [1:0] stalls_id ;  
   reg [1:0] stalls_id_1 ;  
   wire stall=~(auto_in_0_a_bits_source[3])&a_first&(flight_0|flight_1|flight_2|flight_3|flight_4|flight_5|flight_6|flight_7)&(a_noDomain|stalls_id!=a_id)|auto_in_0_a_bits_source[3]&a_first&(flight_8|flight_9|flight_10|flight_11|flight_12|flight_13|flight_14|flight_15)&(a_noDomain|stalls_id_1!=a_id) ;  
   wire nodeIn_a_ready=auto_out_0_a_ready&(auto_in_0_a_bits_address[31]|~stall) ;  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<auto_in_0_a_bits_size ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<auto_out_0_d_bits_size ;  
   wire d_first_first=d_first_counter==9'h0 ;  
   wire _GEN=d_first_first&auto_out_0_d_bits_opcode!=3'h6&auto_in_0_d_ready&auto_out_0_d_valid ;  
   wire _stalls_id_T_4=nodeIn_a_ready&auto_in_0_a_valid ;  
   wire _GEN_0=a_first&_stalls_id_T_4 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              flight_0 <=1'h0;
              flight_1 <=1'h0;
              flight_2 <=1'h0;
              flight_3 <=1'h0;
              flight_4 <=1'h0;
              flight_5 <=1'h0;
              flight_6 <=1'h0;
              flight_7 <=1'h0;
              flight_8 <=1'h0;
              flight_9 <=1'h0;
              flight_10 <=1'h0;
              flight_11 <=1'h0;
              flight_12 <=1'h0;
              flight_13 <=1'h0;
              flight_14 <=1'h0;
              flight_15 <=1'h0;
            end 
          else 
            begin 
              if (_stalls_id_T_4)
                 begin 
                   if (a_first)
                      a_first_counter <=auto_in_0_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                    else 
                      a_first_counter <=a_first_counter-9'h1;
                 end 
              if (auto_in_0_d_ready&auto_out_0_d_valid)
                 begin 
                   if (d_first_first)
                      d_first_counter <=auto_out_0_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                    else 
                      d_first_counter <=d_first_counter-9'h1;
                 end 
              flight_0 <=~(_GEN&auto_out_0_d_bits_source==4'h0)&(_GEN_0&auto_in_0_a_bits_source==4'h0 ? ~(auto_in_0_a_bits_address[31]):flight_0);
              flight_1 <=~(_GEN&auto_out_0_d_bits_source==4'h1)&(_GEN_0&auto_in_0_a_bits_source==4'h1 ? ~(auto_in_0_a_bits_address[31]):flight_1);
              flight_2 <=~(_GEN&auto_out_0_d_bits_source==4'h2)&(_GEN_0&auto_in_0_a_bits_source==4'h2 ? ~(auto_in_0_a_bits_address[31]):flight_2);
              flight_3 <=~(_GEN&auto_out_0_d_bits_source==4'h3)&(_GEN_0&auto_in_0_a_bits_source==4'h3 ? ~(auto_in_0_a_bits_address[31]):flight_3);
              flight_4 <=~(_GEN&auto_out_0_d_bits_source==4'h4)&(_GEN_0&auto_in_0_a_bits_source==4'h4 ? ~(auto_in_0_a_bits_address[31]):flight_4);
              flight_5 <=~(_GEN&auto_out_0_d_bits_source==4'h5)&(_GEN_0&auto_in_0_a_bits_source==4'h5 ? ~(auto_in_0_a_bits_address[31]):flight_5);
              flight_6 <=~(_GEN&auto_out_0_d_bits_source==4'h6)&(_GEN_0&auto_in_0_a_bits_source==4'h6 ? ~(auto_in_0_a_bits_address[31]):flight_6);
              flight_7 <=~(_GEN&auto_out_0_d_bits_source==4'h7)&(_GEN_0&auto_in_0_a_bits_source==4'h7 ? ~(auto_in_0_a_bits_address[31]):flight_7);
              flight_8 <=~(_GEN&auto_out_0_d_bits_source==4'h8)&(_GEN_0&auto_in_0_a_bits_source==4'h8 ? ~(auto_in_0_a_bits_address[31]):flight_8);
              flight_9 <=~(_GEN&auto_out_0_d_bits_source==4'h9)&(_GEN_0&auto_in_0_a_bits_source==4'h9 ? ~(auto_in_0_a_bits_address[31]):flight_9);
              flight_10 <=~(_GEN&auto_out_0_d_bits_source==4'hA)&(_GEN_0&auto_in_0_a_bits_source==4'hA ? ~(auto_in_0_a_bits_address[31]):flight_10);
              flight_11 <=~(_GEN&auto_out_0_d_bits_source==4'hB)&(_GEN_0&auto_in_0_a_bits_source==4'hB ? ~(auto_in_0_a_bits_address[31]):flight_11);
              flight_12 <=~(_GEN&auto_out_0_d_bits_source==4'hC)&(_GEN_0&auto_in_0_a_bits_source==4'hC ? ~(auto_in_0_a_bits_address[31]):flight_12);
              flight_13 <=~(_GEN&auto_out_0_d_bits_source==4'hD)&(_GEN_0&auto_in_0_a_bits_source==4'hD ? ~(auto_in_0_a_bits_address[31]):flight_13);
              flight_14 <=~(_GEN&auto_out_0_d_bits_source==4'hE)&(_GEN_0&auto_in_0_a_bits_source==4'hE ? ~(auto_in_0_a_bits_address[31]):flight_14);
              flight_15 <=~(_GEN&(&auto_out_0_d_bits_source))&(_GEN_0&(&auto_in_0_a_bits_source) ? ~(auto_in_0_a_bits_address[31]):flight_15);
            end 
         if (_stalls_id_T_4&~(auto_in_0_a_bits_source[3])&~(auto_in_0_a_bits_address[31]))
            stalls_id <=a_id;
         if (_stalls_id_T_4&auto_in_0_a_bits_source[3]&~(auto_in_0_a_bits_address[31]))
            stalls_id_1 <=a_id;
       end
  
  TLMonitor_2 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_0_a_valid),.io_in_a_bits_opcode(auto_in_0_a_bits_opcode),.io_in_a_bits_param(auto_in_0_a_bits_param),.io_in_a_bits_size(auto_in_0_a_bits_size),.io_in_a_bits_source(auto_in_0_a_bits_source),.io_in_a_bits_address(auto_in_0_a_bits_address),.io_in_a_bits_mask(auto_in_0_a_bits_mask),.io_in_a_bits_corrupt(auto_in_0_a_bits_corrupt),.io_in_d_ready(auto_in_0_d_ready),.io_in_d_valid(auto_out_0_d_valid),.io_in_d_bits_opcode(auto_out_0_d_bits_opcode),.io_in_d_bits_param(auto_out_0_d_bits_param),.io_in_d_bits_size(auto_out_0_d_bits_size),.io_in_d_bits_source(auto_out_0_d_bits_source),.io_in_d_bits_sink(auto_out_0_d_bits_sink),.io_in_d_bits_denied(auto_out_0_d_bits_denied),.io_in_d_bits_corrupt(auto_out_0_d_bits_corrupt)); 
  TLMonitor_3 monitor_1(.clock(clock),.reset(reset),.io_in_a_ready(auto_out_1_a_ready),.io_in_a_valid(auto_in_1_a_valid),.io_in_a_bits_opcode(auto_in_1_a_bits_opcode),.io_in_a_bits_param(auto_in_1_a_bits_param),.io_in_a_bits_size(auto_in_1_a_bits_size),.io_in_a_bits_source(auto_in_1_a_bits_source),.io_in_a_bits_address(auto_in_1_a_bits_address),.io_in_a_bits_mask(auto_in_1_a_bits_mask),.io_in_a_bits_corrupt(auto_in_1_a_bits_corrupt),.io_in_b_ready(auto_in_1_b_ready),.io_in_b_valid(auto_out_1_b_valid),.io_in_b_bits_param(auto_out_1_b_bits_param),.io_in_b_bits_address(auto_out_1_b_bits_address),.io_in_c_ready(auto_out_1_c_ready),.io_in_c_valid(auto_in_1_c_valid),.io_in_c_bits_opcode(auto_in_1_c_bits_opcode),.io_in_c_bits_param(auto_in_1_c_bits_param),.io_in_c_bits_size(auto_in_1_c_bits_size),.io_in_c_bits_source(auto_in_1_c_bits_source),.io_in_c_bits_address(auto_in_1_c_bits_address),.io_in_c_bits_corrupt(auto_in_1_c_bits_corrupt),.io_in_d_ready(auto_in_1_d_ready),.io_in_d_valid(auto_out_1_d_valid),.io_in_d_bits_opcode(auto_out_1_d_bits_opcode),.io_in_d_bits_param(auto_out_1_d_bits_param),.io_in_d_bits_size(auto_out_1_d_bits_size),.io_in_d_bits_source(auto_out_1_d_bits_source),.io_in_d_bits_sink(auto_out_1_d_bits_sink),.io_in_d_bits_denied(auto_out_1_d_bits_denied),.io_in_d_bits_corrupt(auto_out_1_d_bits_corrupt),.io_in_e_valid(auto_in_1_e_valid),.io_in_e_bits_sink(auto_in_1_e_bits_sink)); 
  assign auto_in_1_a_ready=auto_out_1_a_ready; 
  assign auto_in_1_b_valid=auto_out_1_b_valid; 
  assign auto_in_1_b_bits_param=auto_out_1_b_bits_param; 
  assign auto_in_1_b_bits_address=auto_out_1_b_bits_address; 
  assign auto_in_1_c_ready=auto_out_1_c_ready; 
  assign auto_in_1_d_valid=auto_out_1_d_valid; 
  assign auto_in_1_d_bits_opcode=auto_out_1_d_bits_opcode; 
  assign auto_in_1_d_bits_param=auto_out_1_d_bits_param; 
  assign auto_in_1_d_bits_size=auto_out_1_d_bits_size; 
  assign auto_in_1_d_bits_source=auto_out_1_d_bits_source; 
  assign auto_in_1_d_bits_sink=auto_out_1_d_bits_sink; 
  assign auto_in_1_d_bits_denied=auto_out_1_d_bits_denied; 
  assign auto_in_1_d_bits_data=auto_out_1_d_bits_data; 
  assign auto_in_1_d_bits_corrupt=auto_out_1_d_bits_corrupt; 
  assign auto_in_0_a_ready=nodeIn_a_ready; 
  assign auto_in_0_d_valid=auto_out_0_d_valid; 
  assign auto_in_0_d_bits_opcode=auto_out_0_d_bits_opcode; 
  assign auto_in_0_d_bits_param=auto_out_0_d_bits_param; 
  assign auto_in_0_d_bits_size=auto_out_0_d_bits_size; 
  assign auto_in_0_d_bits_source=auto_out_0_d_bits_source; 
  assign auto_in_0_d_bits_sink=auto_out_0_d_bits_sink; 
  assign auto_in_0_d_bits_denied=auto_out_0_d_bits_denied; 
  assign auto_in_0_d_bits_data=auto_out_0_d_bits_data; 
  assign auto_in_0_d_bits_corrupt=auto_out_0_d_bits_corrupt; 
  assign auto_out_1_a_valid=auto_in_1_a_valid; 
  assign auto_out_1_a_bits_opcode=auto_in_1_a_bits_opcode; 
  assign auto_out_1_a_bits_param=auto_in_1_a_bits_param; 
  assign auto_out_1_a_bits_size=auto_in_1_a_bits_size; 
  assign auto_out_1_a_bits_source=auto_in_1_a_bits_source; 
  assign auto_out_1_a_bits_address=auto_in_1_a_bits_address; 
  assign auto_out_1_a_bits_mask=auto_in_1_a_bits_mask; 
  assign auto_out_1_a_bits_data=auto_in_1_a_bits_data; 
  assign auto_out_1_a_bits_corrupt=auto_in_1_a_bits_corrupt; 
  assign auto_out_1_b_ready=auto_in_1_b_ready; 
  assign auto_out_1_c_valid=auto_in_1_c_valid; 
  assign auto_out_1_c_bits_opcode=auto_in_1_c_bits_opcode; 
  assign auto_out_1_c_bits_param=auto_in_1_c_bits_param; 
  assign auto_out_1_c_bits_size=auto_in_1_c_bits_size; 
  assign auto_out_1_c_bits_source=auto_in_1_c_bits_source; 
  assign auto_out_1_c_bits_address=auto_in_1_c_bits_address; 
  assign auto_out_1_c_bits_data=auto_in_1_c_bits_data; 
  assign auto_out_1_c_bits_corrupt=auto_in_1_c_bits_corrupt; 
  assign auto_out_1_d_ready=auto_in_1_d_ready; 
  assign auto_out_1_e_valid=auto_in_1_e_valid; 
  assign auto_out_1_e_bits_sink=auto_in_1_e_bits_sink; 
  assign auto_out_0_a_valid=auto_in_0_a_valid&(auto_in_0_a_bits_address[31]|~stall); 
  assign auto_out_0_a_bits_opcode=auto_in_0_a_bits_opcode; 
  assign auto_out_0_a_bits_param=auto_in_0_a_bits_param; 
  assign auto_out_0_a_bits_size=auto_in_0_a_bits_size; 
  assign auto_out_0_a_bits_source=auto_in_0_a_bits_source; 
  assign auto_out_0_a_bits_address=auto_in_0_a_bits_address; 
  assign auto_out_0_a_bits_mask=auto_in_0_a_bits_mask; 
  assign auto_out_0_a_bits_data=auto_in_0_a_bits_data; 
  assign auto_out_0_a_bits_corrupt=auto_in_0_a_bits_corrupt; 
  assign auto_out_0_d_ready=auto_in_0_d_ready; 
endmodule
 
module ram_2x4 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [3:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [3:0] W0_data) ; 
   reg [3:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:4'bx; 
endmodule
 
module ram_addr_2x31 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [30:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [30:0] W0_data) ; 
   reg [30:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:31'bx; 
endmodule
 
module ram_2x8 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [7:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [7:0] W0_data) ; 
   reg [7:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:8'bx; 
endmodule
 
module ram_2x3 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [2:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [2:0] W0_data) ; 
   reg [2:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:3'bx; 
endmodule
 
module ram_2x2 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [1:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [1:0] W0_data) ; 
   reg [1:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:2'bx; 
endmodule
 
module ram_2x1 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input W0_data) ; 
   reg Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:1'bx; 
endmodule
 
module Queue (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [30:0] io_enq_bits_addr,
  input [7:0] io_enq_bits_len,
  input [2:0] io_enq_bits_size,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst,
  output io_deq_bits_lock,
  output [3:0] io_deq_bits_cache,
  output [2:0] io_deq_bits_prot,
  output [3:0] io_deq_bits_qos) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x4 ram_id_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_addr_2x31 ram_addr_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_addr),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_addr)); 
  ram_2x8 ram_len_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_len),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_len)); 
  ram_2x3 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_2x2 ram_burst_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_burst),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(2'h1)); 
  ram_2x1 ram_lock_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_lock),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(1'h0)); 
  ram_2x4 ram_cache_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_cache),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(4'h0)); 
  ram_2x3 ram_prot_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_prot),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(3'h2)); 
  ram_2x4 ram_qos_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_qos),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(4'h0)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module ram_data_2x64 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [63:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [63:0] W0_data) ; 
   reg [63:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:64'bx; 
endmodule
 
module Queue_1 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [63:0] io_enq_bits_data,
  input [7:0] io_enq_bits_strb,
  input io_enq_bits_last,
  input io_deq_ready,
  output io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0] io_deq_bits_strb,
  output io_deq_bits_last) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x8 ram_strb_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_strb),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_strb)); 
  ram_2x1 ram_last_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_last),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_last)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_2 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [1:0] io_enq_bits_resp,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x4 ram_id_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_2x2 ram_resp_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_resp),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_resp)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_4 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [63:0] io_enq_bits_data,
  input [1:0] io_enq_bits_resp,
  input io_enq_bits_last,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0] io_deq_bits_resp,
  output io_deq_bits_last) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x4 ram_id_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x2 ram_resp_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_resp),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_resp)); 
  ram_2x1 ram_last_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_last),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_last)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module AXI4Buffer (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [1:0] auto_out_aw_bits_burst,
  output auto_out_aw_bits_lock,
  output [3:0] auto_out_aw_bits_cache,
  output [2:0] auto_out_aw_bits_prot,
  output [3:0] auto_out_aw_bits_qos,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [1:0] auto_out_ar_bits_burst,
  output auto_out_ar_bits_lock,
  output [3:0] auto_out_ar_bits_cache,
  output [2:0] auto_out_ar_bits_prot,
  output [3:0] auto_out_ar_bits_qos,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_last) ; 
  Queue nodeOut_aw_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_aw_ready),.io_enq_valid(auto_in_aw_valid),.io_enq_bits_id(auto_in_aw_bits_id),.io_enq_bits_addr(auto_in_aw_bits_addr),.io_enq_bits_len(auto_in_aw_bits_len),.io_enq_bits_size(auto_in_aw_bits_size),.io_deq_ready(auto_out_aw_ready),.io_deq_valid(auto_out_aw_valid),.io_deq_bits_id(auto_out_aw_bits_id),.io_deq_bits_addr(auto_out_aw_bits_addr),.io_deq_bits_len(auto_out_aw_bits_len),.io_deq_bits_size(auto_out_aw_bits_size),.io_deq_bits_burst(auto_out_aw_bits_burst),.io_deq_bits_lock(auto_out_aw_bits_lock),.io_deq_bits_cache(auto_out_aw_bits_cache),.io_deq_bits_prot(auto_out_aw_bits_prot),.io_deq_bits_qos(auto_out_aw_bits_qos)); 
  Queue_1 nodeOut_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_w_ready),.io_enq_valid(auto_in_w_valid),.io_enq_bits_data(auto_in_w_bits_data),.io_enq_bits_strb(auto_in_w_bits_strb),.io_enq_bits_last(auto_in_w_bits_last),.io_deq_ready(auto_out_w_ready),.io_deq_valid(auto_out_w_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last(auto_out_w_bits_last)); 
  Queue_2 nodeIn_b_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_b_ready),.io_enq_valid(auto_out_b_valid),.io_enq_bits_id(auto_out_b_bits_id),.io_enq_bits_resp(auto_out_b_bits_resp),.io_deq_ready(auto_in_b_ready),.io_deq_valid(auto_in_b_valid),.io_deq_bits_id(auto_in_b_bits_id),.io_deq_bits_resp(auto_in_b_bits_resp)); 
  Queue nodeOut_ar_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_ar_ready),.io_enq_valid(auto_in_ar_valid),.io_enq_bits_id(auto_in_ar_bits_id),.io_enq_bits_addr(auto_in_ar_bits_addr),.io_enq_bits_len(auto_in_ar_bits_len),.io_enq_bits_size(auto_in_ar_bits_size),.io_deq_ready(auto_out_ar_ready),.io_deq_valid(auto_out_ar_valid),.io_deq_bits_id(auto_out_ar_bits_id),.io_deq_bits_addr(auto_out_ar_bits_addr),.io_deq_bits_len(auto_out_ar_bits_len),.io_deq_bits_size(auto_out_ar_bits_size),.io_deq_bits_burst(auto_out_ar_bits_burst),.io_deq_bits_lock(auto_out_ar_bits_lock),.io_deq_bits_cache(auto_out_ar_bits_cache),.io_deq_bits_prot(auto_out_ar_bits_prot),.io_deq_bits_qos(auto_out_ar_bits_qos)); 
  Queue_4 nodeIn_r_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_r_ready),.io_enq_valid(auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_last(auto_out_r_bits_last),.io_deq_ready(auto_in_r_ready),.io_deq_valid(auto_in_r_valid),.io_deq_bits_id(auto_in_r_bits_id),.io_deq_bits_data(auto_in_r_bits_data),.io_deq_bits_resp(auto_in_r_bits_resp),.io_deq_bits_last(auto_in_r_bits_last)); 
endmodule
 
module Queue_5 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_tl_state_size,
  input [4:0] io_enq_bits_tl_state_source,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_tl_state_size,
  output [4:0] io_deq_bits_tl_state_source) ; 
   reg [8:0] ram ;  
   reg full ;  
   wire do_enq=~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            ram <={io_enq_bits_tl_state_source,io_enq_bits_tl_state_size};
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(io_deq_ready&full)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=full; 
  assign io_deq_bits_tl_state_size=ram[3:0]; 
  assign io_deq_bits_tl_state_source=ram[8:4]; 
endmodule
 
module ram_8x9 (
  input [2:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [8:0] R0_data,
  input [2:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [8:0] W0_data) ; 
   reg [8:0] Memory[0:7] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:9'bx; 
endmodule
 
module Queue_6 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_tl_state_size,
  input [4:0] io_enq_bits_tl_state_source,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_tl_state_size,
  output [4:0] io_deq_bits_tl_state_source) ; 
   wire [8:0] _ram_ext_R0_data ;  
   reg [2:0] enq_ptr_value ;  
   reg [2:0] deq_ptr_value ;  
   reg maybe_full ;  
   wire ptr_match=enq_ptr_value==deq_ptr_value ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              enq_ptr_value <=3'h0;
              deq_ptr_value <=3'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 enq_ptr_value <=enq_ptr_value+3'h1;
              if (do_deq)
                 deq_ptr_value <=deq_ptr_value+3'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_8x9 ram_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(_ram_ext_R0_data),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data({io_enq_bits_tl_state_source,io_enq_bits_tl_state_size})); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
  assign io_deq_bits_tl_state_size=_ram_ext_R0_data[3:0]; 
  assign io_deq_bits_tl_state_source=_ram_ext_R0_data[8:4]; 
endmodule
 
module AXI4UserYanker (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [3:0] auto_in_aw_bits_echo_tl_state_size,
  input [4:0] auto_in_aw_bits_echo_tl_state_source,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output [3:0] auto_in_b_bits_echo_tl_state_size,
  output [4:0] auto_in_b_bits_echo_tl_state_source,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [3:0] auto_in_ar_bits_echo_tl_state_size,
  input [4:0] auto_in_ar_bits_echo_tl_state_source,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output [3:0] auto_in_r_bits_echo_tl_state_size,
  output [4:0] auto_in_r_bits_echo_tl_state_source,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_last) ; 
   wire _Queue_9_io_enq_ready ;  
   wire _Queue_9_io_deq_valid ;  
   wire [3:0] _Queue_9_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_9_io_deq_bits_tl_state_source ;  
   wire _Queue_8_io_enq_ready ;  
   wire _Queue_8_io_deq_valid ;  
   wire [3:0] _Queue_8_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_8_io_deq_bits_tl_state_source ;  
   wire _Queue_7_io_enq_ready ;  
   wire _Queue_7_io_deq_valid ;  
   wire [3:0] _Queue_7_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_7_io_deq_bits_tl_state_source ;  
   wire _Queue_6_io_enq_ready ;  
   wire _Queue_6_io_deq_valid ;  
   wire [3:0] _Queue_6_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_6_io_deq_bits_tl_state_source ;  
   wire _Queue_5_io_enq_ready ;  
   wire _Queue_5_io_deq_valid ;  
   wire [3:0] _Queue_5_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_5_io_deq_bits_tl_state_source ;  
   wire _Queue_4_io_enq_ready ;  
   wire _Queue_4_io_deq_valid ;  
   wire [3:0] _Queue_4_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_4_io_deq_bits_tl_state_source ;  
   wire _Queue_3_io_enq_ready ;  
   wire _Queue_3_io_deq_valid ;  
   wire [3:0] _Queue_3_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_3_io_deq_bits_tl_state_source ;  
   wire _Queue_2_io_enq_ready ;  
   wire _Queue_2_io_deq_valid ;  
   wire [3:0] _Queue_2_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_2_io_deq_bits_tl_state_source ;  
   wire _Queue_1_io_enq_ready ;  
   wire _Queue_1_io_deq_valid ;  
   wire [3:0] _Queue_1_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_1_io_deq_bits_tl_state_source ;  
   wire _Queue_io_enq_ready ;  
   wire _Queue_io_deq_valid ;  
   wire [3:0] _Queue_io_deq_bits_tl_state_size ;  
   wire [4:0] _Queue_io_deq_bits_tl_state_source ;  
   reg casez_tmp ;  
  always @(*)
       begin 
         casez (auto_in_ar_bits_id)
          4 'b0000:
             casez_tmp =_Queue_io_enq_ready;
          4 'b0001:
             casez_tmp =_Queue_1_io_enq_ready;
          4 'b0010:
             casez_tmp =_Queue_2_io_enq_ready;
          4 'b0011:
             casez_tmp =_Queue_3_io_enq_ready;
          4 'b0100:
             casez_tmp =_Queue_4_io_enq_ready;
          4 'b0101:
             casez_tmp =1'h0;
          4 'b0110:
             casez_tmp =1'h0;
          4 'b0111:
             casez_tmp =1'h0;
          4 'b1000:
             casez_tmp =1'h0;
          4 'b1001:
             casez_tmp =1'h0;
          4 'b1010:
             casez_tmp =1'h0;
          4 'b1011:
             casez_tmp =1'h0;
          4 'b1100:
             casez_tmp =1'h0;
          4 'b1101:
             casez_tmp =1'h0;
          4 'b1110:
             casez_tmp =1'h0;
          default :
             casez_tmp =1'h0;
         endcase 
       end
  
   reg casez_tmp_0 ;  
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp_0 =_Queue_io_deq_valid;
          4 'b0001:
             casez_tmp_0 =_Queue_1_io_deq_valid;
          4 'b0010:
             casez_tmp_0 =_Queue_2_io_deq_valid;
          4 'b0011:
             casez_tmp_0 =_Queue_3_io_deq_valid;
          4 'b0100:
             casez_tmp_0 =_Queue_4_io_deq_valid;
          4 'b0101:
             casez_tmp_0 =1'h0;
          4 'b0110:
             casez_tmp_0 =1'h0;
          4 'b0111:
             casez_tmp_0 =1'h0;
          4 'b1000:
             casez_tmp_0 =1'h0;
          4 'b1001:
             casez_tmp_0 =1'h0;
          4 'b1010:
             casez_tmp_0 =1'h0;
          4 'b1011:
             casez_tmp_0 =1'h0;
          4 'b1100:
             casez_tmp_0 =1'h0;
          4 'b1101:
             casez_tmp_0 =1'h0;
          4 'b1110:
             casez_tmp_0 =1'h0;
          default :
             casez_tmp_0 =1'h0;
         endcase 
       end
  
   reg [3:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp_1 =_Queue_io_deq_bits_tl_state_size;
          4 'b0001:
             casez_tmp_1 =_Queue_1_io_deq_bits_tl_state_size;
          4 'b0010:
             casez_tmp_1 =_Queue_2_io_deq_bits_tl_state_size;
          4 'b0011:
             casez_tmp_1 =_Queue_3_io_deq_bits_tl_state_size;
          4 'b0100:
             casez_tmp_1 =_Queue_4_io_deq_bits_tl_state_size;
          4 'b0101:
             casez_tmp_1 =4'h0;
          4 'b0110:
             casez_tmp_1 =4'h0;
          4 'b0111:
             casez_tmp_1 =4'h0;
          4 'b1000:
             casez_tmp_1 =4'h0;
          4 'b1001:
             casez_tmp_1 =4'h0;
          4 'b1010:
             casez_tmp_1 =4'h0;
          4 'b1011:
             casez_tmp_1 =4'h0;
          4 'b1100:
             casez_tmp_1 =4'h0;
          4 'b1101:
             casez_tmp_1 =4'h0;
          4 'b1110:
             casez_tmp_1 =4'h0;
          default :
             casez_tmp_1 =4'h0;
         endcase 
       end
  
   reg [4:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp_2 =_Queue_io_deq_bits_tl_state_source;
          4 'b0001:
             casez_tmp_2 =_Queue_1_io_deq_bits_tl_state_source;
          4 'b0010:
             casez_tmp_2 =_Queue_2_io_deq_bits_tl_state_source;
          4 'b0011:
             casez_tmp_2 =_Queue_3_io_deq_bits_tl_state_source;
          4 'b0100:
             casez_tmp_2 =_Queue_4_io_deq_bits_tl_state_source;
          4 'b0101:
             casez_tmp_2 =5'h0;
          4 'b0110:
             casez_tmp_2 =5'h0;
          4 'b0111:
             casez_tmp_2 =5'h0;
          4 'b1000:
             casez_tmp_2 =5'h0;
          4 'b1001:
             casez_tmp_2 =5'h0;
          4 'b1010:
             casez_tmp_2 =5'h0;
          4 'b1011:
             casez_tmp_2 =5'h0;
          4 'b1100:
             casez_tmp_2 =5'h0;
          4 'b1101:
             casez_tmp_2 =5'h0;
          4 'b1110:
             casez_tmp_2 =5'h0;
          default :
             casez_tmp_2 =5'h0;
         endcase 
       end
  
   wire _rqueues_15_deq_ready_T=auto_out_r_valid&auto_in_r_ready ;  
   wire _rqueues_15_enq_valid_T=auto_in_ar_valid&auto_out_ar_ready ;  
   reg casez_tmp_3 ;  
  always @(*)
       begin 
         casez (auto_in_aw_bits_id)
          4 'b0000:
             casez_tmp_3 =_Queue_5_io_enq_ready;
          4 'b0001:
             casez_tmp_3 =_Queue_6_io_enq_ready;
          4 'b0010:
             casez_tmp_3 =_Queue_7_io_enq_ready;
          4 'b0011:
             casez_tmp_3 =_Queue_8_io_enq_ready;
          4 'b0100:
             casez_tmp_3 =_Queue_9_io_enq_ready;
          4 'b0101:
             casez_tmp_3 =1'h0;
          4 'b0110:
             casez_tmp_3 =1'h0;
          4 'b0111:
             casez_tmp_3 =1'h0;
          4 'b1000:
             casez_tmp_3 =1'h0;
          4 'b1001:
             casez_tmp_3 =1'h0;
          4 'b1010:
             casez_tmp_3 =1'h0;
          4 'b1011:
             casez_tmp_3 =1'h0;
          4 'b1100:
             casez_tmp_3 =1'h0;
          4 'b1101:
             casez_tmp_3 =1'h0;
          4 'b1110:
             casez_tmp_3 =1'h0;
          default :
             casez_tmp_3 =1'h0;
         endcase 
       end
  
   reg casez_tmp_4 ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp_4 =_Queue_5_io_deq_valid;
          4 'b0001:
             casez_tmp_4 =_Queue_6_io_deq_valid;
          4 'b0010:
             casez_tmp_4 =_Queue_7_io_deq_valid;
          4 'b0011:
             casez_tmp_4 =_Queue_8_io_deq_valid;
          4 'b0100:
             casez_tmp_4 =_Queue_9_io_deq_valid;
          4 'b0101:
             casez_tmp_4 =1'h0;
          4 'b0110:
             casez_tmp_4 =1'h0;
          4 'b0111:
             casez_tmp_4 =1'h0;
          4 'b1000:
             casez_tmp_4 =1'h0;
          4 'b1001:
             casez_tmp_4 =1'h0;
          4 'b1010:
             casez_tmp_4 =1'h0;
          4 'b1011:
             casez_tmp_4 =1'h0;
          4 'b1100:
             casez_tmp_4 =1'h0;
          4 'b1101:
             casez_tmp_4 =1'h0;
          4 'b1110:
             casez_tmp_4 =1'h0;
          default :
             casez_tmp_4 =1'h0;
         endcase 
       end
  
  always @( posedge clock)
       begin 
         if (~reset&~(~auto_out_r_valid|casez_tmp_0))
            begin 
              if (1)$display("Assertion failed\n    at UserYanker.scala:66 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
              if (1)$display("");
            end 
         if (~reset&~(~auto_out_b_valid|casez_tmp_4))
            begin 
              if (1)$display("Assertion failed\n    at UserYanker.scala:95 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
              if (1)$display("");
            end 
       end
  
   reg [3:0] casez_tmp_5 ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp_5 =_Queue_5_io_deq_bits_tl_state_size;
          4 'b0001:
             casez_tmp_5 =_Queue_6_io_deq_bits_tl_state_size;
          4 'b0010:
             casez_tmp_5 =_Queue_7_io_deq_bits_tl_state_size;
          4 'b0011:
             casez_tmp_5 =_Queue_8_io_deq_bits_tl_state_size;
          4 'b0100:
             casez_tmp_5 =_Queue_9_io_deq_bits_tl_state_size;
          4 'b0101:
             casez_tmp_5 =4'h0;
          4 'b0110:
             casez_tmp_5 =4'h0;
          4 'b0111:
             casez_tmp_5 =4'h0;
          4 'b1000:
             casez_tmp_5 =4'h0;
          4 'b1001:
             casez_tmp_5 =4'h0;
          4 'b1010:
             casez_tmp_5 =4'h0;
          4 'b1011:
             casez_tmp_5 =4'h0;
          4 'b1100:
             casez_tmp_5 =4'h0;
          4 'b1101:
             casez_tmp_5 =4'h0;
          4 'b1110:
             casez_tmp_5 =4'h0;
          default :
             casez_tmp_5 =4'h0;
         endcase 
       end
  
   reg [4:0] casez_tmp_6 ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp_6 =_Queue_5_io_deq_bits_tl_state_source;
          4 'b0001:
             casez_tmp_6 =_Queue_6_io_deq_bits_tl_state_source;
          4 'b0010:
             casez_tmp_6 =_Queue_7_io_deq_bits_tl_state_source;
          4 'b0011:
             casez_tmp_6 =_Queue_8_io_deq_bits_tl_state_source;
          4 'b0100:
             casez_tmp_6 =_Queue_9_io_deq_bits_tl_state_source;
          4 'b0101:
             casez_tmp_6 =5'h0;
          4 'b0110:
             casez_tmp_6 =5'h0;
          4 'b0111:
             casez_tmp_6 =5'h0;
          4 'b1000:
             casez_tmp_6 =5'h0;
          4 'b1001:
             casez_tmp_6 =5'h0;
          4 'b1010:
             casez_tmp_6 =5'h0;
          4 'b1011:
             casez_tmp_6 =5'h0;
          4 'b1100:
             casez_tmp_6 =5'h0;
          4 'b1101:
             casez_tmp_6 =5'h0;
          4 'b1110:
             casez_tmp_6 =5'h0;
          default :
             casez_tmp_6 =5'h0;
         endcase 
       end
  
   wire _wqueues_15_deq_ready_T=auto_out_b_valid&auto_in_b_ready ;  
   wire _wqueues_15_enq_valid_T=auto_in_aw_valid&auto_out_aw_ready ;  
  Queue_5 Queue(.clock(clock),.reset(reset),.io_enq_ready(_Queue_io_enq_ready),.io_enq_valid(_rqueues_15_enq_valid_T&auto_in_ar_bits_id==4'h0),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_deq_ready(_rqueues_15_deq_ready_T&auto_out_r_bits_id==4'h0&auto_out_r_bits_last),.io_deq_valid(_Queue_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_io_deq_bits_tl_state_source)); 
  Queue_6 Queue_1(.clock(clock),.reset(reset),.io_enq_ready(_Queue_1_io_enq_ready),.io_enq_valid(_rqueues_15_enq_valid_T&auto_in_ar_bits_id==4'h1),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_deq_ready(_rqueues_15_deq_ready_T&auto_out_r_bits_id==4'h1&auto_out_r_bits_last),.io_deq_valid(_Queue_1_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_1_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_1_io_deq_bits_tl_state_source)); 
  Queue_6 Queue_2(.clock(clock),.reset(reset),.io_enq_ready(_Queue_2_io_enq_ready),.io_enq_valid(_rqueues_15_enq_valid_T&auto_in_ar_bits_id==4'h2),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_deq_ready(_rqueues_15_deq_ready_T&auto_out_r_bits_id==4'h2&auto_out_r_bits_last),.io_deq_valid(_Queue_2_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_2_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_2_io_deq_bits_tl_state_source)); 
  Queue_5 Queue_3(.clock(clock),.reset(reset),.io_enq_ready(_Queue_3_io_enq_ready),.io_enq_valid(_rqueues_15_enq_valid_T&auto_in_ar_bits_id==4'h3),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_deq_ready(_rqueues_15_deq_ready_T&auto_out_r_bits_id==4'h3&auto_out_r_bits_last),.io_deq_valid(_Queue_3_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_3_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_3_io_deq_bits_tl_state_source)); 
  Queue_5 Queue_4(.clock(clock),.reset(reset),.io_enq_ready(_Queue_4_io_enq_ready),.io_enq_valid(_rqueues_15_enq_valid_T&auto_in_ar_bits_id==4'h4),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_deq_ready(_rqueues_15_deq_ready_T&auto_out_r_bits_id==4'h4&auto_out_r_bits_last),.io_deq_valid(_Queue_4_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_4_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_4_io_deq_bits_tl_state_source)); 
  Queue_5 Queue_5(.clock(clock),.reset(reset),.io_enq_ready(_Queue_5_io_enq_ready),.io_enq_valid(_wqueues_15_enq_valid_T&auto_in_aw_bits_id==4'h0),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_deq_ready(_wqueues_15_deq_ready_T&auto_out_b_bits_id==4'h0),.io_deq_valid(_Queue_5_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_5_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_5_io_deq_bits_tl_state_source)); 
  Queue_6 Queue_6(.clock(clock),.reset(reset),.io_enq_ready(_Queue_6_io_enq_ready),.io_enq_valid(_wqueues_15_enq_valid_T&auto_in_aw_bits_id==4'h1),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_deq_ready(_wqueues_15_deq_ready_T&auto_out_b_bits_id==4'h1),.io_deq_valid(_Queue_6_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_6_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_6_io_deq_bits_tl_state_source)); 
  Queue_6 Queue_7(.clock(clock),.reset(reset),.io_enq_ready(_Queue_7_io_enq_ready),.io_enq_valid(_wqueues_15_enq_valid_T&auto_in_aw_bits_id==4'h2),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_deq_ready(_wqueues_15_deq_ready_T&auto_out_b_bits_id==4'h2),.io_deq_valid(_Queue_7_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_7_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_7_io_deq_bits_tl_state_source)); 
  Queue_5 Queue_8(.clock(clock),.reset(reset),.io_enq_ready(_Queue_8_io_enq_ready),.io_enq_valid(_wqueues_15_enq_valid_T&auto_in_aw_bits_id==4'h3),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_deq_ready(_wqueues_15_deq_ready_T&auto_out_b_bits_id==4'h3),.io_deq_valid(_Queue_8_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_8_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_8_io_deq_bits_tl_state_source)); 
  Queue_5 Queue_9(.clock(clock),.reset(reset),.io_enq_ready(_Queue_9_io_enq_ready),.io_enq_valid(_wqueues_15_enq_valid_T&auto_in_aw_bits_id==4'h4),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_deq_ready(_wqueues_15_deq_ready_T&auto_out_b_bits_id==4'h4),.io_deq_valid(_Queue_9_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_9_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_9_io_deq_bits_tl_state_source)); 
  assign auto_in_aw_ready=auto_out_aw_ready&casez_tmp_3; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_b_bits_echo_tl_state_size=casez_tmp_5; 
  assign auto_in_b_bits_echo_tl_state_source=casez_tmp_6; 
  assign auto_in_ar_ready=auto_out_ar_ready&casez_tmp; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_echo_tl_state_size=casez_tmp_1; 
  assign auto_in_r_bits_echo_tl_state_source=casez_tmp_2; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid&casez_tmp_3; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid&casez_tmp; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module ram_id_8x4 (
  input [2:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [3:0] R0_data,
  input [2:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [3:0] W0_data) ; 
   reg [3:0] Memory[0:7] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:4'bx; 
endmodule
 
module ram_data_8x64 (
  input [2:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [63:0] R0_data,
  input [2:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [63:0] W0_data) ; 
   reg [63:0] Memory[0:7] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:64'bx; 
endmodule
 
module ram_resp_8x2 (
  input [2:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [1:0] R0_data,
  input [2:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [1:0] W0_data) ; 
   reg [1:0] Memory[0:7] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:2'bx; 
endmodule
 
module ram_last_8x1 (
  input [2:0] R0_addr,
  input R0_en,
  input R0_clk,
  output R0_data,
  input [2:0] W0_addr,
  input W0_en,
  input W0_clk,
  input W0_data) ; 
   reg Memory[0:7] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:1'bx; 
endmodule
 
module Queue_15 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [63:0] io_enq_bits_data,
  input [1:0] io_enq_bits_resp,
  input [3:0] io_enq_bits_echo_tl_state_size,
  input [4:0] io_enq_bits_echo_tl_state_source,
  input io_enq_bits_last,
  input io_deq_ready,
  output [3:0] io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0] io_deq_bits_resp,
  output [3:0] io_deq_bits_echo_tl_state_size,
  output [4:0] io_deq_bits_echo_tl_state_source,
  output io_deq_bits_last) ; 
   wire [8:0] _ram_echo_ext_R0_data ;  
   reg [2:0] enq_ptr_value ;  
   reg [2:0] deq_ptr_value ;  
   reg maybe_full ;  
   wire ptr_match=enq_ptr_value==deq_ptr_value ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~(ptr_match&~maybe_full) ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              enq_ptr_value <=3'h0;
              deq_ptr_value <=3'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 enq_ptr_value <=enq_ptr_value+3'h1;
              if (do_deq)
                 deq_ptr_value <=deq_ptr_value+3'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_id_8x4 ram_id_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_data_8x64 ram_data_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_resp_8x2 ram_resp_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_resp),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_resp)); 
  ram_8x9 ram_echo_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(_ram_echo_ext_R0_data),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data({io_enq_bits_echo_tl_state_source,io_enq_bits_echo_tl_state_size})); 
  ram_last_8x1 ram_last_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_last),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_last)); 
  assign io_enq_ready=~full; 
  assign io_deq_bits_echo_tl_state_size=_ram_echo_ext_R0_data[3:0]; 
  assign io_deq_bits_echo_tl_state_source=_ram_echo_ext_R0_data[8:4]; 
endmodule
 
module AXI4Deinterleaver (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [3:0] auto_in_aw_bits_echo_tl_state_size,
  input [4:0] auto_in_aw_bits_echo_tl_state_source,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output [3:0] auto_in_b_bits_echo_tl_state_size,
  output [4:0] auto_in_b_bits_echo_tl_state_source,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [3:0] auto_in_ar_bits_echo_tl_state_size,
  input [4:0] auto_in_ar_bits_echo_tl_state_source,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output [3:0] auto_in_r_bits_echo_tl_state_size,
  output [4:0] auto_in_r_bits_echo_tl_state_source,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [3:0] auto_out_aw_bits_echo_tl_state_size,
  output [4:0] auto_out_aw_bits_echo_tl_state_source,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input [3:0] auto_out_b_bits_echo_tl_state_size,
  input [4:0] auto_out_b_bits_echo_tl_state_source,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [3:0] auto_out_ar_bits_echo_tl_state_size,
  output [4:0] auto_out_ar_bits_echo_tl_state_source,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input [3:0] auto_out_r_bits_echo_tl_state_size,
  input [4:0] auto_out_r_bits_echo_tl_state_source,
  input auto_out_r_bits_last) ; 
   reg casez_tmp ;  
   wire enq_OH_bools_15 ;  
   wire enq_OH_bools_14 ;  
   wire enq_OH_bools_13 ;  
   wire enq_OH_bools_12 ;  
   wire enq_OH_bools_11 ;  
   wire enq_OH_bools_10 ;  
   wire enq_OH_bools_9 ;  
   wire enq_OH_bools_8 ;  
   wire enq_OH_bools_7 ;  
   wire enq_OH_bools_6 ;  
   wire enq_OH_bools_5 ;  
   reg casez_tmp_0 ;  
   wire _qs_queue_4_io_enq_ready ;  
   wire [3:0] _qs_queue_4_io_deq_bits_id ;  
   wire [63:0] _qs_queue_4_io_deq_bits_data ;  
   wire [1:0] _qs_queue_4_io_deq_bits_resp ;  
   wire [3:0] _qs_queue_4_io_deq_bits_echo_tl_state_size ;  
   wire [4:0] _qs_queue_4_io_deq_bits_echo_tl_state_source ;  
   wire _qs_queue_4_io_deq_bits_last ;  
   wire _qs_queue_3_io_enq_ready ;  
   wire [3:0] _qs_queue_3_io_deq_bits_id ;  
   wire [63:0] _qs_queue_3_io_deq_bits_data ;  
   wire [1:0] _qs_queue_3_io_deq_bits_resp ;  
   wire [3:0] _qs_queue_3_io_deq_bits_echo_tl_state_size ;  
   wire [4:0] _qs_queue_3_io_deq_bits_echo_tl_state_source ;  
   wire _qs_queue_3_io_deq_bits_last ;  
   wire _qs_queue_2_io_enq_ready ;  
   wire [3:0] _qs_queue_2_io_deq_bits_id ;  
   wire [63:0] _qs_queue_2_io_deq_bits_data ;  
   wire [1:0] _qs_queue_2_io_deq_bits_resp ;  
   wire [3:0] _qs_queue_2_io_deq_bits_echo_tl_state_size ;  
   wire [4:0] _qs_queue_2_io_deq_bits_echo_tl_state_source ;  
   wire _qs_queue_2_io_deq_bits_last ;  
   wire _qs_queue_1_io_enq_ready ;  
   wire [3:0] _qs_queue_1_io_deq_bits_id ;  
   wire [63:0] _qs_queue_1_io_deq_bits_data ;  
   wire [1:0] _qs_queue_1_io_deq_bits_resp ;  
   wire [3:0] _qs_queue_1_io_deq_bits_echo_tl_state_size ;  
   wire [4:0] _qs_queue_1_io_deq_bits_echo_tl_state_source ;  
   wire _qs_queue_1_io_deq_bits_last ;  
   wire _qs_queue_0_io_enq_ready ;  
   wire [3:0] _qs_queue_0_io_deq_bits_id ;  
   wire [63:0] _qs_queue_0_io_deq_bits_data ;  
   wire [1:0] _qs_queue_0_io_deq_bits_resp ;  
   wire [3:0] _qs_queue_0_io_deq_bits_echo_tl_state_size ;  
   wire [4:0] _qs_queue_0_io_deq_bits_echo_tl_state_source ;  
   wire _qs_queue_0_io_deq_bits_last ;  
   reg locked ;  
   reg [3:0] deq_id ;  
   reg [3:0] pending_count ;  
   wire enq_OH_bools_0=auto_out_r_bits_id==4'h0 ;  
   wire _pending_inc_T_13=casez_tmp&auto_out_r_valid ;  
   wire pending_inc=enq_OH_bools_0&_pending_inc_T_13&auto_out_r_bits_last ;  
   wire deq_OH_bools_0=deq_id==4'h0 ;  
   wire _queue_wire_15_deq_ready_T=auto_in_r_ready&locked ;  
   wire pending_dec=deq_OH_bools_0&_queue_wire_15_deq_ready_T&casez_tmp_0 ;  
   reg [3:0] pending_count_1 ;  
   wire enq_OH_bools_1=auto_out_r_bits_id==4'h1 ;  
   wire pending_inc_1=enq_OH_bools_1&_pending_inc_T_13&auto_out_r_bits_last ;  
   wire deq_OH_bools_1=deq_id==4'h1 ;  
   wire pending_dec_1=deq_OH_bools_1&_queue_wire_15_deq_ready_T&casez_tmp_0 ;  
   reg [3:0] pending_count_2 ;  
   wire enq_OH_bools_2=auto_out_r_bits_id==4'h2 ;  
   wire pending_inc_2=enq_OH_bools_2&_pending_inc_T_13&auto_out_r_bits_last ;  
   wire deq_OH_bools_2=deq_id==4'h2 ;  
   wire pending_dec_2=deq_OH_bools_2&_queue_wire_15_deq_ready_T&casez_tmp_0 ;  
   reg [3:0] pending_count_3 ;  
   wire enq_OH_bools_3=auto_out_r_bits_id==4'h3 ;  
   wire pending_inc_3=enq_OH_bools_3&_pending_inc_T_13&auto_out_r_bits_last ;  
   wire deq_OH_bools_3=deq_id==4'h3 ;  
   wire pending_dec_3=deq_OH_bools_3&_queue_wire_15_deq_ready_T&casez_tmp_0 ;  
   reg [3:0] pending_count_4 ;  
   wire enq_OH_bools_4=auto_out_r_bits_id==4'h4 ;  
   wire pending_inc_4=enq_OH_bools_4&_pending_inc_T_13&auto_out_r_bits_last ;  
   wire deq_OH_bools_4=deq_id==4'h4 ;  
   wire pending_dec_4=deq_OH_bools_4&_queue_wire_15_deq_ready_T&casez_tmp_0 ;  
  always @( posedge clock)
       begin 
         if (~reset&enq_OH_bools_5&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 5 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_6&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 6 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_7&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 7 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_8&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 8 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_9&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 9 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_10&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 10 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_11&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 11 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_12&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 12 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_13&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 13 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_14&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 14 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&enq_OH_bools_15&auto_out_r_valid)
            begin 
              if (1)$display("Assertion failed: ID 15 should not be used\n    at Deinterleaver.scala:76 assert(!q.enq.valid, s\"ID ${i} should not be used\")\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_dec|(|pending_count)))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:100 assert (!dec || count =/= 0.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_inc|pending_count!=4'h8))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:101 assert (!inc || count =/= beats.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_dec_1|(|pending_count_1)))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:100 assert (!dec || count =/= 0.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_inc_1|pending_count_1!=4'h8))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:101 assert (!inc || count =/= beats.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_dec_2|(|pending_count_2)))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:100 assert (!dec || count =/= 0.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_inc_2|pending_count_2!=4'h8))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:101 assert (!inc || count =/= beats.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_dec_3|(|pending_count_3)))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:100 assert (!dec || count =/= 0.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_inc_3|pending_count_3!=4'h8))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:101 assert (!inc || count =/= beats.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_dec_4|(|pending_count_4)))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:100 assert (!dec || count =/= 0.U)\n");
              if (1)$display("");
            end 
         if (~reset&~(~pending_inc_4|pending_count_4!=4'h8))
            begin 
              if (1)$display("Assertion failed\n    at Deinterleaver.scala:101 assert (!inc || count =/= beats.U)\n");
              if (1)$display("");
            end 
       end
  
   reg [3:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (deq_id)
          4 'b0000:
             casez_tmp_1 =_qs_queue_0_io_deq_bits_id;
          4 'b0001:
             casez_tmp_1 =_qs_queue_1_io_deq_bits_id;
          4 'b0010:
             casez_tmp_1 =_qs_queue_2_io_deq_bits_id;
          4 'b0011:
             casez_tmp_1 =_qs_queue_3_io_deq_bits_id;
          4 'b0100:
             casez_tmp_1 =_qs_queue_4_io_deq_bits_id;
          4 'b0101:
             casez_tmp_1 =4'h0;
          4 'b0110:
             casez_tmp_1 =4'h0;
          4 'b0111:
             casez_tmp_1 =4'h0;
          4 'b1000:
             casez_tmp_1 =4'h0;
          4 'b1001:
             casez_tmp_1 =4'h0;
          4 'b1010:
             casez_tmp_1 =4'h0;
          4 'b1011:
             casez_tmp_1 =4'h0;
          4 'b1100:
             casez_tmp_1 =4'h0;
          4 'b1101:
             casez_tmp_1 =4'h0;
          4 'b1110:
             casez_tmp_1 =4'h0;
          default :
             casez_tmp_1 =4'h0;
         endcase 
       end
  
   reg [63:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (deq_id)
          4 'b0000:
             casez_tmp_2 =_qs_queue_0_io_deq_bits_data;
          4 'b0001:
             casez_tmp_2 =_qs_queue_1_io_deq_bits_data;
          4 'b0010:
             casez_tmp_2 =_qs_queue_2_io_deq_bits_data;
          4 'b0011:
             casez_tmp_2 =_qs_queue_3_io_deq_bits_data;
          4 'b0100:
             casez_tmp_2 =_qs_queue_4_io_deq_bits_data;
          4 'b0101:
             casez_tmp_2 =64'h0;
          4 'b0110:
             casez_tmp_2 =64'h0;
          4 'b0111:
             casez_tmp_2 =64'h0;
          4 'b1000:
             casez_tmp_2 =64'h0;
          4 'b1001:
             casez_tmp_2 =64'h0;
          4 'b1010:
             casez_tmp_2 =64'h0;
          4 'b1011:
             casez_tmp_2 =64'h0;
          4 'b1100:
             casez_tmp_2 =64'h0;
          4 'b1101:
             casez_tmp_2 =64'h0;
          4 'b1110:
             casez_tmp_2 =64'h0;
          default :
             casez_tmp_2 =64'h0;
         endcase 
       end
  
   reg [1:0] casez_tmp_3 ;  
  always @(*)
       begin 
         casez (deq_id)
          4 'b0000:
             casez_tmp_3 =_qs_queue_0_io_deq_bits_resp;
          4 'b0001:
             casez_tmp_3 =_qs_queue_1_io_deq_bits_resp;
          4 'b0010:
             casez_tmp_3 =_qs_queue_2_io_deq_bits_resp;
          4 'b0011:
             casez_tmp_3 =_qs_queue_3_io_deq_bits_resp;
          4 'b0100:
             casez_tmp_3 =_qs_queue_4_io_deq_bits_resp;
          4 'b0101:
             casez_tmp_3 =2'h0;
          4 'b0110:
             casez_tmp_3 =2'h0;
          4 'b0111:
             casez_tmp_3 =2'h0;
          4 'b1000:
             casez_tmp_3 =2'h0;
          4 'b1001:
             casez_tmp_3 =2'h0;
          4 'b1010:
             casez_tmp_3 =2'h0;
          4 'b1011:
             casez_tmp_3 =2'h0;
          4 'b1100:
             casez_tmp_3 =2'h0;
          4 'b1101:
             casez_tmp_3 =2'h0;
          4 'b1110:
             casez_tmp_3 =2'h0;
          default :
             casez_tmp_3 =2'h0;
         endcase 
       end
  
   reg [3:0] casez_tmp_4 ;  
  always @(*)
       begin 
         casez (deq_id)
          4 'b0000:
             casez_tmp_4 =_qs_queue_0_io_deq_bits_echo_tl_state_size;
          4 'b0001:
             casez_tmp_4 =_qs_queue_1_io_deq_bits_echo_tl_state_size;
          4 'b0010:
             casez_tmp_4 =_qs_queue_2_io_deq_bits_echo_tl_state_size;
          4 'b0011:
             casez_tmp_4 =_qs_queue_3_io_deq_bits_echo_tl_state_size;
          4 'b0100:
             casez_tmp_4 =_qs_queue_4_io_deq_bits_echo_tl_state_size;
          4 'b0101:
             casez_tmp_4 =4'h0;
          4 'b0110:
             casez_tmp_4 =4'h0;
          4 'b0111:
             casez_tmp_4 =4'h0;
          4 'b1000:
             casez_tmp_4 =4'h0;
          4 'b1001:
             casez_tmp_4 =4'h0;
          4 'b1010:
             casez_tmp_4 =4'h0;
          4 'b1011:
             casez_tmp_4 =4'h0;
          4 'b1100:
             casez_tmp_4 =4'h0;
          4 'b1101:
             casez_tmp_4 =4'h0;
          4 'b1110:
             casez_tmp_4 =4'h0;
          default :
             casez_tmp_4 =4'h0;
         endcase 
       end
  
   reg [4:0] casez_tmp_5 ;  
  always @(*)
       begin 
         casez (deq_id)
          4 'b0000:
             casez_tmp_5 =_qs_queue_0_io_deq_bits_echo_tl_state_source;
          4 'b0001:
             casez_tmp_5 =_qs_queue_1_io_deq_bits_echo_tl_state_source;
          4 'b0010:
             casez_tmp_5 =_qs_queue_2_io_deq_bits_echo_tl_state_source;
          4 'b0011:
             casez_tmp_5 =_qs_queue_3_io_deq_bits_echo_tl_state_source;
          4 'b0100:
             casez_tmp_5 =_qs_queue_4_io_deq_bits_echo_tl_state_source;
          4 'b0101:
             casez_tmp_5 =5'h0;
          4 'b0110:
             casez_tmp_5 =5'h0;
          4 'b0111:
             casez_tmp_5 =5'h0;
          4 'b1000:
             casez_tmp_5 =5'h0;
          4 'b1001:
             casez_tmp_5 =5'h0;
          4 'b1010:
             casez_tmp_5 =5'h0;
          4 'b1011:
             casez_tmp_5 =5'h0;
          4 'b1100:
             casez_tmp_5 =5'h0;
          4 'b1101:
             casez_tmp_5 =5'h0;
          4 'b1110:
             casez_tmp_5 =5'h0;
          default :
             casez_tmp_5 =5'h0;
         endcase 
       end
  
  always @(*)
       begin 
         casez (deq_id)
          4 'b0000:
             casez_tmp_0 =_qs_queue_0_io_deq_bits_last;
          4 'b0001:
             casez_tmp_0 =_qs_queue_1_io_deq_bits_last;
          4 'b0010:
             casez_tmp_0 =_qs_queue_2_io_deq_bits_last;
          4 'b0011:
             casez_tmp_0 =_qs_queue_3_io_deq_bits_last;
          4 'b0100:
             casez_tmp_0 =_qs_queue_4_io_deq_bits_last;
          4 'b0101:
             casez_tmp_0 =1'h0;
          4 'b0110:
             casez_tmp_0 =1'h0;
          4 'b0111:
             casez_tmp_0 =1'h0;
          4 'b1000:
             casez_tmp_0 =1'h0;
          4 'b1001:
             casez_tmp_0 =1'h0;
          4 'b1010:
             casez_tmp_0 =1'h0;
          4 'b1011:
             casez_tmp_0 =1'h0;
          4 'b1100:
             casez_tmp_0 =1'h0;
          4 'b1101:
             casez_tmp_0 =1'h0;
          4 'b1110:
             casez_tmp_0 =1'h0;
          default :
             casez_tmp_0 =1'h0;
         endcase 
       end
  
  assign enq_OH_bools_5=auto_out_r_bits_id==4'h5; 
  assign enq_OH_bools_6=auto_out_r_bits_id==4'h6; 
  assign enq_OH_bools_7=auto_out_r_bits_id==4'h7; 
  assign enq_OH_bools_8=auto_out_r_bits_id==4'h8; 
  assign enq_OH_bools_9=auto_out_r_bits_id==4'h9; 
  assign enq_OH_bools_10=auto_out_r_bits_id==4'hA; 
  assign enq_OH_bools_11=auto_out_r_bits_id==4'hB; 
  assign enq_OH_bools_12=auto_out_r_bits_id==4'hC; 
  assign enq_OH_bools_13=auto_out_r_bits_id==4'hD; 
  assign enq_OH_bools_14=auto_out_r_bits_id==4'hE; 
  assign enq_OH_bools_15=&auto_out_r_bits_id; 
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp =_qs_queue_0_io_enq_ready;
          4 'b0001:
             casez_tmp =_qs_queue_1_io_enq_ready;
          4 'b0010:
             casez_tmp =_qs_queue_2_io_enq_ready;
          4 'b0011:
             casez_tmp =_qs_queue_3_io_enq_ready;
          4 'b0100:
             casez_tmp =_qs_queue_4_io_enq_ready;
          4 'b0101:
             casez_tmp =1'h0;
          4 'b0110:
             casez_tmp =1'h0;
          4 'b0111:
             casez_tmp =1'h0;
          4 'b1000:
             casez_tmp =1'h0;
          4 'b1001:
             casez_tmp =1'h0;
          4 'b1010:
             casez_tmp =1'h0;
          4 'b1011:
             casez_tmp =1'h0;
          4 'b1100:
             casez_tmp =1'h0;
          4 'b1101:
             casez_tmp =1'h0;
          4 'b1110:
             casez_tmp =1'h0;
          default :
             casez_tmp =1'h0;
         endcase 
       end
  
   wire [3:0] _pending_next_T_2=pending_count+{3'h0,pending_inc}-{3'h0,pending_dec} ;  
   wire [3:0] _pending_next_T_6=pending_count_1+{3'h0,pending_inc_1}-{3'h0,pending_dec_1} ;  
   wire [3:0] _pending_next_T_10=pending_count_2+{3'h0,pending_inc_2}-{3'h0,pending_dec_2} ;  
   wire [3:0] _pending_next_T_14=pending_count_3+{3'h0,pending_inc_3}-{3'h0,pending_dec_3} ;  
   wire [3:0] _pending_next_T_18=pending_count_4+{3'h0,pending_inc_4}-{3'h0,pending_dec_4} ;  
   wire _GEN=~locked|_queue_wire_15_deq_ready_T&casez_tmp_0 ;  
   wire _GEN_0=(|_pending_next_T_18)|(|_pending_next_T_14) ;  
   wire _GEN_1=(|_pending_next_T_14)|(|_pending_next_T_10) ;  
   wire _GEN_2=(|_pending_next_T_10)|(|_pending_next_T_6) ;  
   wire _GEN_3=(|_pending_next_T_6)|(|_pending_next_T_2) ;  
   wire _GEN_4=_GEN_1|_GEN_3 ;  
   wire _GEN_5=_GEN_2|(|_pending_next_T_2) ;  
   wire _GEN_6=(|_pending_next_T_18)|_GEN_4 ;  
   wire _GEN_7=_GEN_0|_GEN_5 ;  
   wire _GEN_8=(|_pending_next_T_18)|_GEN_1|_GEN_3 ;  
   wire _GEN_9=_GEN_0|_GEN_2|(|_pending_next_T_2) ;  
   wire [14:0] deq_id_lo={~_GEN_7,~_GEN_8,~_GEN_9,~_GEN_6,~_GEN_7,~_GEN_8,~_GEN_9,~_GEN_6,~_GEN_7,~_GEN_8,~_GEN_9,~_GEN_4,~_GEN_5,~_GEN_3,~(|_pending_next_T_2)}&{11'h0,|_pending_next_T_18,|_pending_next_T_14,|_pending_next_T_10,|_pending_next_T_6} ;  
   wire [6:0] _deq_id_T_3=deq_id_lo[14:8]|deq_id_lo[6:0] ;  
   wire [2:0] _deq_id_T_5=_deq_id_T_3[6:4]|_deq_id_T_3[2:0] ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              locked <=1'h0;
              pending_count <=4'h0;
              pending_count_1 <=4'h0;
              pending_count_2 <=4'h0;
              pending_count_3 <=4'h0;
              pending_count_4 <=4'h0;
            end 
          else 
            begin 
              if (_GEN)
                 locked <=|{|_pending_next_T_18,|_pending_next_T_14,|_pending_next_T_10,|_pending_next_T_6,|_pending_next_T_2};
              pending_count <=_pending_next_T_2;
              pending_count_1 <=_pending_next_T_6;
              pending_count_2 <=_pending_next_T_10;
              pending_count_3 <=_pending_next_T_14;
              pending_count_4 <=_pending_next_T_18;
            end 
         if (_GEN)
            deq_id <={|(deq_id_lo[14:7]),|(_deq_id_T_3[6:3]),|(_deq_id_T_5[2:1]),_deq_id_T_5[2]|_deq_id_T_5[0]};
       end
  
  Queue_15 qs_queue_0(.clock(clock),.reset(reset),.io_enq_ready(_qs_queue_0_io_enq_ready),.io_enq_valid(enq_OH_bools_0&auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_echo_tl_state_size(auto_out_r_bits_echo_tl_state_size),.io_enq_bits_echo_tl_state_source(auto_out_r_bits_echo_tl_state_source),.io_enq_bits_last(auto_out_r_bits_last),.io_deq_ready(deq_OH_bools_0&_queue_wire_15_deq_ready_T),.io_deq_bits_id(_qs_queue_0_io_deq_bits_id),.io_deq_bits_data(_qs_queue_0_io_deq_bits_data),.io_deq_bits_resp(_qs_queue_0_io_deq_bits_resp),.io_deq_bits_echo_tl_state_size(_qs_queue_0_io_deq_bits_echo_tl_state_size),.io_deq_bits_echo_tl_state_source(_qs_queue_0_io_deq_bits_echo_tl_state_source),.io_deq_bits_last(_qs_queue_0_io_deq_bits_last)); 
  Queue_15 qs_queue_1(.clock(clock),.reset(reset),.io_enq_ready(_qs_queue_1_io_enq_ready),.io_enq_valid(enq_OH_bools_1&auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_echo_tl_state_size(auto_out_r_bits_echo_tl_state_size),.io_enq_bits_echo_tl_state_source(auto_out_r_bits_echo_tl_state_source),.io_enq_bits_last(auto_out_r_bits_last),.io_deq_ready(deq_OH_bools_1&_queue_wire_15_deq_ready_T),.io_deq_bits_id(_qs_queue_1_io_deq_bits_id),.io_deq_bits_data(_qs_queue_1_io_deq_bits_data),.io_deq_bits_resp(_qs_queue_1_io_deq_bits_resp),.io_deq_bits_echo_tl_state_size(_qs_queue_1_io_deq_bits_echo_tl_state_size),.io_deq_bits_echo_tl_state_source(_qs_queue_1_io_deq_bits_echo_tl_state_source),.io_deq_bits_last(_qs_queue_1_io_deq_bits_last)); 
  Queue_15 qs_queue_2(.clock(clock),.reset(reset),.io_enq_ready(_qs_queue_2_io_enq_ready),.io_enq_valid(enq_OH_bools_2&auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_echo_tl_state_size(auto_out_r_bits_echo_tl_state_size),.io_enq_bits_echo_tl_state_source(auto_out_r_bits_echo_tl_state_source),.io_enq_bits_last(auto_out_r_bits_last),.io_deq_ready(deq_OH_bools_2&_queue_wire_15_deq_ready_T),.io_deq_bits_id(_qs_queue_2_io_deq_bits_id),.io_deq_bits_data(_qs_queue_2_io_deq_bits_data),.io_deq_bits_resp(_qs_queue_2_io_deq_bits_resp),.io_deq_bits_echo_tl_state_size(_qs_queue_2_io_deq_bits_echo_tl_state_size),.io_deq_bits_echo_tl_state_source(_qs_queue_2_io_deq_bits_echo_tl_state_source),.io_deq_bits_last(_qs_queue_2_io_deq_bits_last)); 
  Queue_15 qs_queue_3(.clock(clock),.reset(reset),.io_enq_ready(_qs_queue_3_io_enq_ready),.io_enq_valid(enq_OH_bools_3&auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_echo_tl_state_size(auto_out_r_bits_echo_tl_state_size),.io_enq_bits_echo_tl_state_source(auto_out_r_bits_echo_tl_state_source),.io_enq_bits_last(auto_out_r_bits_last),.io_deq_ready(deq_OH_bools_3&_queue_wire_15_deq_ready_T),.io_deq_bits_id(_qs_queue_3_io_deq_bits_id),.io_deq_bits_data(_qs_queue_3_io_deq_bits_data),.io_deq_bits_resp(_qs_queue_3_io_deq_bits_resp),.io_deq_bits_echo_tl_state_size(_qs_queue_3_io_deq_bits_echo_tl_state_size),.io_deq_bits_echo_tl_state_source(_qs_queue_3_io_deq_bits_echo_tl_state_source),.io_deq_bits_last(_qs_queue_3_io_deq_bits_last)); 
  Queue_15 qs_queue_4(.clock(clock),.reset(reset),.io_enq_ready(_qs_queue_4_io_enq_ready),.io_enq_valid(enq_OH_bools_4&auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_echo_tl_state_size(auto_out_r_bits_echo_tl_state_size),.io_enq_bits_echo_tl_state_source(auto_out_r_bits_echo_tl_state_source),.io_enq_bits_last(auto_out_r_bits_last),.io_deq_ready(deq_OH_bools_4&_queue_wire_15_deq_ready_T),.io_deq_bits_id(_qs_queue_4_io_deq_bits_id),.io_deq_bits_data(_qs_queue_4_io_deq_bits_data),.io_deq_bits_resp(_qs_queue_4_io_deq_bits_resp),.io_deq_bits_echo_tl_state_size(_qs_queue_4_io_deq_bits_echo_tl_state_size),.io_deq_bits_echo_tl_state_source(_qs_queue_4_io_deq_bits_echo_tl_state_source),.io_deq_bits_last(_qs_queue_4_io_deq_bits_last)); 
  assign auto_in_aw_ready=auto_out_aw_ready; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_b_bits_echo_tl_state_size=auto_out_b_bits_echo_tl_state_size; 
  assign auto_in_b_bits_echo_tl_state_source=auto_out_b_bits_echo_tl_state_source; 
  assign auto_in_ar_ready=auto_out_ar_ready; 
  assign auto_in_r_valid=locked; 
  assign auto_in_r_bits_id=casez_tmp_1; 
  assign auto_in_r_bits_data=casez_tmp_2; 
  assign auto_in_r_bits_resp=casez_tmp_3; 
  assign auto_in_r_bits_echo_tl_state_size=casez_tmp_4; 
  assign auto_in_r_bits_echo_tl_state_source=casez_tmp_5; 
  assign auto_in_r_bits_last=casez_tmp_0; 
  assign auto_out_aw_valid=auto_in_aw_valid; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_aw_bits_echo_tl_state_size=auto_in_aw_bits_echo_tl_state_size; 
  assign auto_out_aw_bits_echo_tl_state_source=auto_in_aw_bits_echo_tl_state_source; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_ar_bits_echo_tl_state_size=auto_in_ar_bits_echo_tl_state_size; 
  assign auto_out_ar_bits_echo_tl_state_source=auto_in_ar_bits_echo_tl_state_source; 
  assign auto_out_r_ready=casez_tmp; 
endmodule
 
module AXI4IdIndexer (
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [2:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [3:0] auto_in_aw_bits_echo_tl_state_size,
  input [4:0] auto_in_aw_bits_echo_tl_state_source,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [2:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output [3:0] auto_in_b_bits_echo_tl_state_size,
  output [4:0] auto_in_b_bits_echo_tl_state_source,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [2:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [3:0] auto_in_ar_bits_echo_tl_state_size,
  input [4:0] auto_in_ar_bits_echo_tl_state_source,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [2:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output [3:0] auto_in_r_bits_echo_tl_state_size,
  output [4:0] auto_in_r_bits_echo_tl_state_source,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [3:0] auto_out_aw_bits_echo_tl_state_size,
  output [4:0] auto_out_aw_bits_echo_tl_state_source,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input [3:0] auto_out_b_bits_echo_tl_state_size,
  input [4:0] auto_out_b_bits_echo_tl_state_source,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [3:0] auto_out_ar_bits_echo_tl_state_size,
  output [4:0] auto_out_ar_bits_echo_tl_state_source,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input [3:0] auto_out_r_bits_echo_tl_state_size,
  input [4:0] auto_out_r_bits_echo_tl_state_source,
  input auto_out_r_bits_last) ; 
  assign auto_in_aw_ready=auto_out_aw_ready; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id=auto_out_b_bits_id[2:0]; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_b_bits_echo_tl_state_size=auto_out_b_bits_echo_tl_state_size; 
  assign auto_in_b_bits_echo_tl_state_source=auto_out_b_bits_echo_tl_state_source; 
  assign auto_in_ar_ready=auto_out_ar_ready; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id[2:0]; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_echo_tl_state_size=auto_out_r_bits_echo_tl_state_size; 
  assign auto_in_r_bits_echo_tl_state_source=auto_out_r_bits_echo_tl_state_source; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid; 
  assign auto_out_aw_bits_id={1'h0,auto_in_aw_bits_id}; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_aw_bits_echo_tl_state_size=auto_in_aw_bits_echo_tl_state_size; 
  assign auto_out_aw_bits_echo_tl_state_source=auto_in_aw_bits_echo_tl_state_source; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid; 
  assign auto_out_ar_bits_id={1'h0,auto_in_ar_bits_id}; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_ar_bits_echo_tl_state_size=auto_in_ar_bits_echo_tl_state_size; 
  assign auto_out_ar_bits_echo_tl_state_source=auto_in_ar_bits_echo_tl_state_source; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module TLMonitor_4 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [30:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [3:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [22:0] _GEN={19'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [4:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [4:0] source ;  
   reg [30:0] address ;  
   reg [4:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [3:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg denied ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [151:0] inflight_sizes ;  
   reg [4:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==5'h0 ;  
   reg [4:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==5'h0 ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>{69'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _GEN_0={27'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [31:0] _GEN_2={27'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [151:0] inflight_sizes_1 ;  
   reg [4:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==5'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [22:0] _is_aligned_mask_T_1=23'hFF<<_GEN ;  
   wire [7:0] _GEN_3=io_in_a_bits_address[7:0]&~(_is_aligned_mask_T_1[7:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=_source_ok_T_12&io_in_a_bits_size==4'h6&_GEN_4&(&(io_in_a_bits_address[30:29])) ;  
   wire _GEN_7=io_in_a_bits_param>3'h2 ;  
   wire _GEN_8=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_9=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_10=_GEN_4&(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14) ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_12=io_in_a_bits_mask!=mask ;  
   wire _GEN_13=_GEN_10&io_in_a_bits_size<4'h9&(&(io_in_a_bits_address[30:29])) ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_17=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_19=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_20=io_in_d_bits_size<4'h3 ;  
   wire _GEN_21=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_22=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_23=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_24=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_25=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_26=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_27=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_28=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [151:0] _GEN_29={144'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [31:0] _a_set_wo_ready_T=32'h1<<_GEN_0 ;  
   wire [18:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_30=io_in_d_valid&d_first_1 ;  
   wire _GEN_31=_GEN_30&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_32={14'h0,io_in_d_bits_source} ;  
   wire _GEN_33=_GEN_31&same_cycle_resp&~reset ;  
   wire _GEN_34=_GEN_31&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_35={4'h0,io_in_d_bits_size} ;  
   wire _GEN_36=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_37=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_38=inflight>>_GEN_32 ;  
   wire [151:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_29 ;  
   wire [31:0] _d_clr_wo_ready_T=32'h1<<_GEN_2 ;  
   wire [18:0] _GEN_39=inflight_1>>_GEN_32 ;  
   wire [151:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_29 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(io_in_a_bits_size<4'h7&(&(io_in_a_bits_address[30:29]))))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_37[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~reset&~(_GEN_38[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&_GEN_35!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_31 ? _d_clr_wo_ready_T[18:0]:19'h0)|a_set_wo_ready==19'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~(_GEN_39[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&_GEN_35!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:126:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [22:0] _a_first_beats1_decode_T_1=23'hFF<<_GEN ;  
   wire [22:0] _a_first_beats1_decode_T_5=23'hFF<<_GEN ;  
   wire [22:0] _GEN_40={19'h0,io_in_d_bits_size} ;  
   wire [22:0] _d_first_beats1_decode_T_1=23'hFF<<_GEN_40 ;  
   wire [22:0] _d_first_beats1_decode_T_5=23'hFF<<_GEN_40 ;  
   wire [22:0] _d_first_beats1_decode_T_9=23'hFF<<_GEN_40 ;  
   wire [270:0] _GEN_41={263'h0,io_in_d_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_2 ;  
   wire [31:0] _a_set_T=32'h1<<_GEN_0 ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<{264'h0,io_in_d_bits_source,2'h0} ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _d_sizes_clr_T_5=271'hFF<<_GEN_41 ;  
   wire [259:0] _a_sizes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{252'h0,io_in_a_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_2 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hFF<<_GEN_41 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_42=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_43=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=5'h0;
              d_first_counter <=5'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=152'h0;
              a_first_counter_1 <=5'h0;
              d_first_counter_1 <=5'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=152'h0;
              d_first_counter_2 <=5'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-5'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 5'h0:~(_a_first_beats1_decode_T_1[7:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 5'h0:~(_a_first_beats1_decode_T_5[7:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-5'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-5'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[7:3]):5'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[7:3]):5'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-5'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[7:3]):5'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-5'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[18:0]:19'h0))&~(_GEN_42 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_42 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[151:0]:152'h0))&~(_GEN_42 ? _d_sizes_clr_T_5[151:0]:152'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_43 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_43 ? _d_sizes_clr_T_11[151:0]:152'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module Queue_20 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [63:0] io_enq_bits_data,
  input [7:0] io_enq_bits_strb,
  input io_enq_bits_last,
  input io_deq_ready,
  output io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0] io_deq_bits_strb,
  output io_deq_bits_last) ; 
   reg ram_last ;  
   reg [7:0] ram_strb ;  
   reg [63:0] ram_data ;  
   reg full ;  
   wire io_enq_ready_0=io_deq_ready|~full ;  
   wire do_enq=io_enq_ready_0&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_last <=io_enq_bits_last;
              ram_strb <=io_enq_bits_strb;
              ram_data <=io_enq_bits_data;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(io_deq_ready&full)))
               full <=do_enq;
       end
  
  assign io_enq_ready=io_enq_ready_0; 
  assign io_deq_valid=full; 
  assign io_deq_bits_data=ram_data; 
  assign io_deq_bits_strb=ram_strb; 
  assign io_deq_bits_last=ram_last; 
endmodule
 
module Queue_21 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_id,
  input [30:0] io_enq_bits_addr,
  input [7:0] io_enq_bits_len,
  input [2:0] io_enq_bits_size,
  input [3:0] io_enq_bits_echo_tl_state_size,
  input [4:0] io_enq_bits_echo_tl_state_source,
  input io_enq_bits_wen,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [3:0] io_deq_bits_echo_tl_state_size,
  output [4:0] io_deq_bits_echo_tl_state_source,
  output io_deq_bits_wen) ; 
   reg ram_wen ;  
   reg [2:0] ram_size ;  
   reg [7:0] ram_len ;  
   reg [30:0] ram_addr ;  
   reg [2:0] ram_id ;  
   reg [8:0] ram_echo ;  
   reg full ;  
   wire io_enq_ready_0=io_deq_ready|~full ;  
   wire do_enq=io_enq_ready_0&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_wen <=io_enq_bits_wen;
              ram_size <=io_enq_bits_size;
              ram_len <=io_enq_bits_len;
              ram_addr <=io_enq_bits_addr;
              ram_id <=io_enq_bits_id;
              ram_echo <={io_enq_bits_echo_tl_state_source,io_enq_bits_echo_tl_state_size};
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(io_deq_ready&full)))
               full <=do_enq;
       end
  
  assign io_enq_ready=io_enq_ready_0; 
  assign io_deq_valid=full; 
  assign io_deq_bits_id=ram_id; 
  assign io_deq_bits_addr=ram_addr; 
  assign io_deq_bits_len=ram_len; 
  assign io_deq_bits_size=ram_size; 
  assign io_deq_bits_echo_tl_state_size=ram_echo[3:0]; 
  assign io_deq_bits_echo_tl_state_source=ram_echo[8:4]; 
  assign io_deq_bits_wen=ram_wen; 
endmodule
 
module TLToAXI4 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [30:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [3:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [2:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [3:0] auto_out_aw_bits_echo_tl_state_size,
  output [4:0] auto_out_aw_bits_echo_tl_state_source,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [2:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input [3:0] auto_out_b_bits_echo_tl_state_size,
  input [4:0] auto_out_b_bits_echo_tl_state_source,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [2:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [3:0] auto_out_ar_bits_echo_tl_state_size,
  output [4:0] auto_out_ar_bits_echo_tl_state_source,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [2:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input [3:0] auto_out_r_bits_echo_tl_state_size,
  input [4:0] auto_out_r_bits_echo_tl_state_source,
  input auto_out_r_bits_last) ; 
   reg count_5 ;  
   reg count_4 ;  
   reg write_2 ;  
   reg [3:0] count_3 ;  
   reg write_1 ;  
   reg [3:0] count_2 ;  
   reg count_1 ;  
   wire _queue_arw_deq_q_io_enq_ready ;  
   wire _queue_arw_deq_q_io_deq_valid ;  
   wire [2:0] _queue_arw_deq_q_io_deq_bits_id ;  
   wire [30:0] _queue_arw_deq_q_io_deq_bits_addr ;  
   wire [7:0] _queue_arw_deq_q_io_deq_bits_len ;  
   wire [2:0] _queue_arw_deq_q_io_deq_bits_size ;  
   wire [3:0] _queue_arw_deq_q_io_deq_bits_echo_tl_state_size ;  
   wire [4:0] _queue_arw_deq_q_io_deq_bits_echo_tl_state_source ;  
   wire _queue_arw_deq_q_io_deq_bits_wen ;  
   wire _nodeOut_w_deq_q_io_enq_ready ;  
   wire [22:0] _beats1_decode_T_1=23'hFF<<auto_in_a_bits_size ;  
   wire [4:0] beats1=auto_in_a_bits_opcode[2] ? 5'h0:~(_beats1_decode_T_1[7:3]) ;  
   reg [4:0] counter ;  
   wire a_first=counter==5'h0 ;  
   wire a_last=counter==5'h1|beats1==5'h0 ;  
   reg doneAW ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_source)
          5 'b00000:
             casez_tmp =3'h1;
          5 'b00001:
             casez_tmp =3'h1;
          5 'b00010:
             casez_tmp =3'h1;
          5 'b00011:
             casez_tmp =3'h1;
          5 'b00100:
             casez_tmp =3'h1;
          5 'b00101:
             casez_tmp =3'h1;
          5 'b00110:
             casez_tmp =3'h1;
          5 'b00111:
             casez_tmp =3'h1;
          5 'b01000:
             casez_tmp =3'h2;
          5 'b01001:
             casez_tmp =3'h2;
          5 'b01010:
             casez_tmp =3'h2;
          5 'b01011:
             casez_tmp =3'h2;
          5 'b01100:
             casez_tmp =3'h2;
          5 'b01101:
             casez_tmp =3'h2;
          5 'b01110:
             casez_tmp =3'h2;
          5 'b01111:
             casez_tmp =3'h2;
          5 'b10000:
             casez_tmp =3'h4;
          5 'b10001:
             casez_tmp =3'h3;
          5 'b10010:
             casez_tmp =3'h0;
          5 'b10011:
             casez_tmp =3'h1;
          5 'b10100:
             casez_tmp =3'h1;
          5 'b10101:
             casez_tmp =3'h1;
          5 'b10110:
             casez_tmp =3'h1;
          5 'b10111:
             casez_tmp =3'h1;
          5 'b11000:
             casez_tmp =3'h1;
          5 'b11001:
             casez_tmp =3'h1;
          5 'b11010:
             casez_tmp =3'h1;
          5 'b11011:
             casez_tmp =3'h1;
          5 'b11100:
             casez_tmp =3'h1;
          5 'b11101:
             casez_tmp =3'h1;
          5 'b11110:
             casez_tmp =3'h1;
          default :
             casez_tmp =3'h1;
         endcase 
       end
  
   wire [25:0] _out_arw_bits_len_T_1=26'h7FF<<auto_in_a_bits_size ;  
   reg casez_tmp_0 ;  
   wire idStall_1=(|count_2)&write_1!=~(auto_in_a_bits_opcode[2])|count_2==4'h8 ;  
   wire idStall_2=(|count_3)&write_2!=~(auto_in_a_bits_opcode[2])|count_3==4'h8 ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_source)
          5 'b00000:
             casez_tmp_0 =idStall_1;
          5 'b00001:
             casez_tmp_0 =idStall_1;
          5 'b00010:
             casez_tmp_0 =idStall_1;
          5 'b00011:
             casez_tmp_0 =idStall_1;
          5 'b00100:
             casez_tmp_0 =idStall_1;
          5 'b00101:
             casez_tmp_0 =idStall_1;
          5 'b00110:
             casez_tmp_0 =idStall_1;
          5 'b00111:
             casez_tmp_0 =idStall_1;
          5 'b01000:
             casez_tmp_0 =idStall_2;
          5 'b01001:
             casez_tmp_0 =idStall_2;
          5 'b01010:
             casez_tmp_0 =idStall_2;
          5 'b01011:
             casez_tmp_0 =idStall_2;
          5 'b01100:
             casez_tmp_0 =idStall_2;
          5 'b01101:
             casez_tmp_0 =idStall_2;
          5 'b01110:
             casez_tmp_0 =idStall_2;
          5 'b01111:
             casez_tmp_0 =idStall_2;
          5 'b10000:
             casez_tmp_0 =count_5;
          5 'b10001:
             casez_tmp_0 =count_4;
          5 'b10010:
             casez_tmp_0 =count_1;
          5 'b10011:
             casez_tmp_0 =idStall_1;
          5 'b10100:
             casez_tmp_0 =idStall_1;
          5 'b10101:
             casez_tmp_0 =idStall_1;
          5 'b10110:
             casez_tmp_0 =idStall_1;
          5 'b10111:
             casez_tmp_0 =idStall_1;
          5 'b11000:
             casez_tmp_0 =idStall_1;
          5 'b11001:
             casez_tmp_0 =idStall_1;
          5 'b11010:
             casez_tmp_0 =idStall_1;
          5 'b11011:
             casez_tmp_0 =idStall_1;
          5 'b11100:
             casez_tmp_0 =idStall_1;
          5 'b11101:
             casez_tmp_0 =idStall_1;
          5 'b11110:
             casez_tmp_0 =idStall_1;
          default :
             casez_tmp_0 =idStall_1;
         endcase 
       end
  
   wire stall=casez_tmp_0&a_first ;  
   wire _out_w_valid_T_3=doneAW|_queue_arw_deq_q_io_enq_ready ;  
   wire nodeIn_a_ready=~stall&(auto_in_a_bits_opcode[2] ? _queue_arw_deq_q_io_enq_ready:_out_w_valid_T_3&_nodeOut_w_deq_q_io_enq_ready) ;  
   wire out_arw_valid=~stall&auto_in_a_valid&(auto_in_a_bits_opcode[2]|~doneAW&_nodeOut_w_deq_q_io_enq_ready) ;  
   reg r_holds_d ;  
   reg [2:0] b_delay ;  
   wire r_wins=auto_out_r_valid&b_delay!=3'h7|r_holds_d ;  
   wire nodeOut_r_ready=auto_in_d_ready&r_wins ;  
   wire nodeOut_b_ready=auto_in_d_ready&~r_wins ;  
   wire nodeIn_d_valid=r_wins ? auto_out_r_valid:auto_out_b_valid ;  
   reg r_first ;  
   reg r_denied_r ;  
   wire r_denied=r_first ? (&auto_out_r_bits_resp):r_denied_r ;  
   wire [2:0] nodeIn_d_bits_opcode={2'h0,r_wins} ;  
   wire [3:0] nodeIn_d_bits_size=r_wins ? auto_out_r_bits_echo_tl_state_size:auto_out_b_bits_echo_tl_state_size ;  
   wire [4:0] nodeIn_d_bits_source=r_wins ? auto_out_r_bits_echo_tl_state_source:auto_out_b_bits_echo_tl_state_source ;  
   wire nodeIn_d_bits_denied=r_wins ? r_denied:(|auto_out_b_bits_resp) ;  
   wire nodeIn_d_bits_corrupt=r_wins&((|auto_out_r_bits_resp)|r_denied) ;  
   wire [2:0] d_sel_shiftAmount=r_wins ? auto_out_r_bits_id:auto_out_b_bits_id ;  
   wire d_last=~r_wins|auto_out_r_bits_last ;  
   wire _inc_T_4=_queue_arw_deq_q_io_enq_ready&out_arw_valid ;  
   wire inc=casez_tmp==3'h0&_inc_T_4 ;  
   wire _dec_T_9=auto_in_d_ready&nodeIn_d_valid ;  
   wire dec=d_sel_shiftAmount==3'h0&d_last&_dec_T_9 ;  
   wire inc_1=casez_tmp==3'h1&_inc_T_4 ;  
   wire dec_1=d_sel_shiftAmount==3'h1&d_last&_dec_T_9 ;  
   wire inc_2=casez_tmp==3'h2&_inc_T_4 ;  
   wire dec_2=d_sel_shiftAmount==3'h2&d_last&_dec_T_9 ;  
   wire inc_3=casez_tmp==3'h3&_inc_T_4 ;  
   wire dec_3=d_sel_shiftAmount==3'h3&d_last&_dec_T_9 ;  
   wire inc_4=casez_tmp==3'h4&_inc_T_4 ;  
   wire dec_4=d_sel_shiftAmount==3'h4&d_last&_dec_T_9 ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~dec|count_1))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc|~count_1))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_1|(|count_2)))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_1|count_2!=4'h8))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_2|(|count_3)))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_2|count_3!=4'h8))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_3|count_4))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_3|~count_4))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_4|count_5))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_4|~count_5))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
       end
  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              counter <=5'h0;
              doneAW <=1'h0;
              r_holds_d <=1'h0;
              r_first <=1'h1;
              count_1 <=1'h0;
              count_2 <=4'h0;
              count_3 <=4'h0;
              count_4 <=1'h0;
              count_5 <=1'h0;
            end 
          else 
            begin 
              if (nodeIn_a_ready&auto_in_a_valid)
                 begin 
                   if (a_first)
                      counter <=beats1;
                    else 
                      counter <=counter-5'h1;
                   doneAW <=~a_last;
                 end 
              if (nodeOut_r_ready&auto_out_r_valid)
                 begin 
                   r_holds_d <=~auto_out_r_bits_last;
                   r_first <=auto_out_r_bits_last;
                 end 
              count_1 <=count_1+inc-dec;
              count_2 <=count_2+{3'h0,inc_1}-{3'h0,dec_1};
              count_3 <=count_3+{3'h0,inc_2}-{3'h0,dec_2};
              count_4 <=count_4+inc_3-dec_3;
              count_5 <=count_5+inc_4-dec_4;
            end 
         if (auto_out_b_valid&~nodeOut_b_ready)
            b_delay <=b_delay+3'h1;
          else 
            b_delay <=3'h0;
         if (r_first)
            r_denied_r <=&auto_out_r_bits_resp;
         if (inc_1)
            write_1 <=~(auto_in_a_bits_opcode[2]);
         if (inc_2)
            write_2 <=~(auto_in_a_bits_opcode[2]);
       end
  
  TLMonitor_4 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(nodeIn_d_bits_opcode),.io_in_d_bits_size(nodeIn_d_bits_size),.io_in_d_bits_source(nodeIn_d_bits_source),.io_in_d_bits_denied(nodeIn_d_bits_denied),.io_in_d_bits_corrupt(nodeIn_d_bits_corrupt)); 
  Queue_20 nodeOut_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_w_deq_q_io_enq_ready),.io_enq_valid(~stall&auto_in_a_valid&~(auto_in_a_bits_opcode[2])&_out_w_valid_T_3),.io_enq_bits_data(auto_in_a_bits_data),.io_enq_bits_strb(auto_in_a_bits_mask),.io_enq_bits_last(a_last),.io_deq_ready(auto_out_w_ready),.io_deq_valid(auto_out_w_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last(auto_out_w_bits_last)); 
  Queue_21 queue_arw_deq_q(.clock(clock),.reset(reset),.io_enq_ready(_queue_arw_deq_q_io_enq_ready),.io_enq_valid(out_arw_valid),.io_enq_bits_id(casez_tmp),.io_enq_bits_addr(auto_in_a_bits_address),.io_enq_bits_len(~(_out_arw_bits_len_T_1[10:3])),.io_enq_bits_size(auto_in_a_bits_size>4'h2 ? 3'h3:auto_in_a_bits_size[2:0]),.io_enq_bits_echo_tl_state_size(auto_in_a_bits_size),.io_enq_bits_echo_tl_state_source(auto_in_a_bits_source),.io_enq_bits_wen(~(auto_in_a_bits_opcode[2])),.io_deq_ready(_queue_arw_deq_q_io_deq_bits_wen ? auto_out_aw_ready:auto_out_ar_ready),.io_deq_valid(_queue_arw_deq_q_io_deq_valid),.io_deq_bits_id(_queue_arw_deq_q_io_deq_bits_id),.io_deq_bits_addr(_queue_arw_deq_q_io_deq_bits_addr),.io_deq_bits_len(_queue_arw_deq_q_io_deq_bits_len),.io_deq_bits_size(_queue_arw_deq_q_io_deq_bits_size),.io_deq_bits_echo_tl_state_size(_queue_arw_deq_q_io_deq_bits_echo_tl_state_size),.io_deq_bits_echo_tl_state_source(_queue_arw_deq_q_io_deq_bits_echo_tl_state_source),.io_deq_bits_wen(_queue_arw_deq_q_io_deq_bits_wen)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=nodeIn_d_bits_opcode; 
  assign auto_in_d_bits_size=nodeIn_d_bits_size; 
  assign auto_in_d_bits_source=nodeIn_d_bits_source; 
  assign auto_in_d_bits_denied=nodeIn_d_bits_denied; 
  assign auto_in_d_bits_data=auto_out_r_bits_data; 
  assign auto_in_d_bits_corrupt=nodeIn_d_bits_corrupt; 
  assign auto_out_aw_valid=_queue_arw_deq_q_io_deq_valid&_queue_arw_deq_q_io_deq_bits_wen; 
  assign auto_out_aw_bits_id=_queue_arw_deq_q_io_deq_bits_id; 
  assign auto_out_aw_bits_addr=_queue_arw_deq_q_io_deq_bits_addr; 
  assign auto_out_aw_bits_len=_queue_arw_deq_q_io_deq_bits_len; 
  assign auto_out_aw_bits_size=_queue_arw_deq_q_io_deq_bits_size; 
  assign auto_out_aw_bits_echo_tl_state_size=_queue_arw_deq_q_io_deq_bits_echo_tl_state_size; 
  assign auto_out_aw_bits_echo_tl_state_source=_queue_arw_deq_q_io_deq_bits_echo_tl_state_source; 
  assign auto_out_b_ready=nodeOut_b_ready; 
  assign auto_out_ar_valid=_queue_arw_deq_q_io_deq_valid&~_queue_arw_deq_q_io_deq_bits_wen; 
  assign auto_out_ar_bits_id=_queue_arw_deq_q_io_deq_bits_id; 
  assign auto_out_ar_bits_addr=_queue_arw_deq_q_io_deq_bits_addr; 
  assign auto_out_ar_bits_len=_queue_arw_deq_q_io_deq_bits_len; 
  assign auto_out_ar_bits_size=_queue_arw_deq_q_io_deq_bits_size; 
  assign auto_out_ar_bits_echo_tl_state_size=_queue_arw_deq_q_io_deq_bits_echo_tl_state_size; 
  assign auto_out_ar_bits_echo_tl_state_source=_queue_arw_deq_q_io_deq_bits_echo_tl_state_source; 
  assign auto_out_r_ready=nodeOut_r_ready; 
endmodule
 
module TLInterconnectCoupler_4 (
  input clock,
  input reset,
  input auto_axi4buf_out_aw_ready,
  output auto_axi4buf_out_aw_valid,
  output [3:0] auto_axi4buf_out_aw_bits_id,
  output [30:0] auto_axi4buf_out_aw_bits_addr,
  output [7:0] auto_axi4buf_out_aw_bits_len,
  output [2:0] auto_axi4buf_out_aw_bits_size,
  output [1:0] auto_axi4buf_out_aw_bits_burst,
  output auto_axi4buf_out_aw_bits_lock,
  output [3:0] auto_axi4buf_out_aw_bits_cache,
  output [2:0] auto_axi4buf_out_aw_bits_prot,
  output [3:0] auto_axi4buf_out_aw_bits_qos,
  input auto_axi4buf_out_w_ready,
  output auto_axi4buf_out_w_valid,
  output [63:0] auto_axi4buf_out_w_bits_data,
  output [7:0] auto_axi4buf_out_w_bits_strb,
  output auto_axi4buf_out_w_bits_last,
  output auto_axi4buf_out_b_ready,
  input auto_axi4buf_out_b_valid,
  input [3:0] auto_axi4buf_out_b_bits_id,
  input [1:0] auto_axi4buf_out_b_bits_resp,
  input auto_axi4buf_out_ar_ready,
  output auto_axi4buf_out_ar_valid,
  output [3:0] auto_axi4buf_out_ar_bits_id,
  output [30:0] auto_axi4buf_out_ar_bits_addr,
  output [7:0] auto_axi4buf_out_ar_bits_len,
  output [2:0] auto_axi4buf_out_ar_bits_size,
  output [1:0] auto_axi4buf_out_ar_bits_burst,
  output auto_axi4buf_out_ar_bits_lock,
  output [3:0] auto_axi4buf_out_ar_bits_cache,
  output [2:0] auto_axi4buf_out_ar_bits_prot,
  output [3:0] auto_axi4buf_out_ar_bits_qos,
  output auto_axi4buf_out_r_ready,
  input auto_axi4buf_out_r_valid,
  input [3:0] auto_axi4buf_out_r_bits_id,
  input [63:0] auto_axi4buf_out_r_bits_data,
  input [1:0] auto_axi4buf_out_r_bits_resp,
  input auto_axi4buf_out_r_bits_last,
  output auto_tl_in_a_ready,
  input auto_tl_in_a_valid,
  input [2:0] auto_tl_in_a_bits_opcode,
  input [2:0] auto_tl_in_a_bits_param,
  input [3:0] auto_tl_in_a_bits_size,
  input [4:0] auto_tl_in_a_bits_source,
  input [30:0] auto_tl_in_a_bits_address,
  input [7:0] auto_tl_in_a_bits_mask,
  input [63:0] auto_tl_in_a_bits_data,
  input auto_tl_in_a_bits_corrupt,
  input auto_tl_in_d_ready,
  output auto_tl_in_d_valid,
  output [2:0] auto_tl_in_d_bits_opcode,
  output [3:0] auto_tl_in_d_bits_size,
  output [4:0] auto_tl_in_d_bits_source,
  output auto_tl_in_d_bits_denied,
  output [63:0] auto_tl_in_d_bits_data,
  output auto_tl_in_d_bits_corrupt) ; 
   wire _tl2axi4_auto_out_aw_valid ;  
   wire [2:0] _tl2axi4_auto_out_aw_bits_id ;  
   wire [30:0] _tl2axi4_auto_out_aw_bits_addr ;  
   wire [7:0] _tl2axi4_auto_out_aw_bits_len ;  
   wire [2:0] _tl2axi4_auto_out_aw_bits_size ;  
   wire [3:0] _tl2axi4_auto_out_aw_bits_echo_tl_state_size ;  
   wire [4:0] _tl2axi4_auto_out_aw_bits_echo_tl_state_source ;  
   wire _tl2axi4_auto_out_w_valid ;  
   wire [63:0] _tl2axi4_auto_out_w_bits_data ;  
   wire [7:0] _tl2axi4_auto_out_w_bits_strb ;  
   wire _tl2axi4_auto_out_w_bits_last ;  
   wire _tl2axi4_auto_out_b_ready ;  
   wire _tl2axi4_auto_out_ar_valid ;  
   wire [2:0] _tl2axi4_auto_out_ar_bits_id ;  
   wire [30:0] _tl2axi4_auto_out_ar_bits_addr ;  
   wire [7:0] _tl2axi4_auto_out_ar_bits_len ;  
   wire [2:0] _tl2axi4_auto_out_ar_bits_size ;  
   wire [3:0] _tl2axi4_auto_out_ar_bits_echo_tl_state_size ;  
   wire [4:0] _tl2axi4_auto_out_ar_bits_echo_tl_state_source ;  
   wire _tl2axi4_auto_out_r_ready ;  
   wire _axi4index_auto_in_aw_ready ;  
   wire _axi4index_auto_in_w_ready ;  
   wire _axi4index_auto_in_b_valid ;  
   wire [2:0] _axi4index_auto_in_b_bits_id ;  
   wire [1:0] _axi4index_auto_in_b_bits_resp ;  
   wire [3:0] _axi4index_auto_in_b_bits_echo_tl_state_size ;  
   wire [4:0] _axi4index_auto_in_b_bits_echo_tl_state_source ;  
   wire _axi4index_auto_in_ar_ready ;  
   wire _axi4index_auto_in_r_valid ;  
   wire [2:0] _axi4index_auto_in_r_bits_id ;  
   wire [63:0] _axi4index_auto_in_r_bits_data ;  
   wire [1:0] _axi4index_auto_in_r_bits_resp ;  
   wire [3:0] _axi4index_auto_in_r_bits_echo_tl_state_size ;  
   wire [4:0] _axi4index_auto_in_r_bits_echo_tl_state_source ;  
   wire _axi4index_auto_in_r_bits_last ;  
   wire _axi4index_auto_out_aw_valid ;  
   wire [3:0] _axi4index_auto_out_aw_bits_id ;  
   wire [30:0] _axi4index_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4index_auto_out_aw_bits_len ;  
   wire [2:0] _axi4index_auto_out_aw_bits_size ;  
   wire [3:0] _axi4index_auto_out_aw_bits_echo_tl_state_size ;  
   wire [4:0] _axi4index_auto_out_aw_bits_echo_tl_state_source ;  
   wire _axi4index_auto_out_w_valid ;  
   wire [63:0] _axi4index_auto_out_w_bits_data ;  
   wire [7:0] _axi4index_auto_out_w_bits_strb ;  
   wire _axi4index_auto_out_w_bits_last ;  
   wire _axi4index_auto_out_b_ready ;  
   wire _axi4index_auto_out_ar_valid ;  
   wire [3:0] _axi4index_auto_out_ar_bits_id ;  
   wire [30:0] _axi4index_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4index_auto_out_ar_bits_len ;  
   wire [2:0] _axi4index_auto_out_ar_bits_size ;  
   wire [3:0] _axi4index_auto_out_ar_bits_echo_tl_state_size ;  
   wire [4:0] _axi4index_auto_out_ar_bits_echo_tl_state_source ;  
   wire _axi4index_auto_out_r_ready ;  
   wire _axi4deint_auto_in_aw_ready ;  
   wire _axi4deint_auto_in_w_ready ;  
   wire _axi4deint_auto_in_b_valid ;  
   wire [3:0] _axi4deint_auto_in_b_bits_id ;  
   wire [1:0] _axi4deint_auto_in_b_bits_resp ;  
   wire [3:0] _axi4deint_auto_in_b_bits_echo_tl_state_size ;  
   wire [4:0] _axi4deint_auto_in_b_bits_echo_tl_state_source ;  
   wire _axi4deint_auto_in_ar_ready ;  
   wire _axi4deint_auto_in_r_valid ;  
   wire [3:0] _axi4deint_auto_in_r_bits_id ;  
   wire [63:0] _axi4deint_auto_in_r_bits_data ;  
   wire [1:0] _axi4deint_auto_in_r_bits_resp ;  
   wire [3:0] _axi4deint_auto_in_r_bits_echo_tl_state_size ;  
   wire [4:0] _axi4deint_auto_in_r_bits_echo_tl_state_source ;  
   wire _axi4deint_auto_in_r_bits_last ;  
   wire _axi4deint_auto_out_aw_valid ;  
   wire [3:0] _axi4deint_auto_out_aw_bits_id ;  
   wire [30:0] _axi4deint_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4deint_auto_out_aw_bits_len ;  
   wire [2:0] _axi4deint_auto_out_aw_bits_size ;  
   wire [3:0] _axi4deint_auto_out_aw_bits_echo_tl_state_size ;  
   wire [4:0] _axi4deint_auto_out_aw_bits_echo_tl_state_source ;  
   wire _axi4deint_auto_out_w_valid ;  
   wire [63:0] _axi4deint_auto_out_w_bits_data ;  
   wire [7:0] _axi4deint_auto_out_w_bits_strb ;  
   wire _axi4deint_auto_out_w_bits_last ;  
   wire _axi4deint_auto_out_b_ready ;  
   wire _axi4deint_auto_out_ar_valid ;  
   wire [3:0] _axi4deint_auto_out_ar_bits_id ;  
   wire [30:0] _axi4deint_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4deint_auto_out_ar_bits_len ;  
   wire [2:0] _axi4deint_auto_out_ar_bits_size ;  
   wire [3:0] _axi4deint_auto_out_ar_bits_echo_tl_state_size ;  
   wire [4:0] _axi4deint_auto_out_ar_bits_echo_tl_state_source ;  
   wire _axi4deint_auto_out_r_ready ;  
   wire _axi4yank_auto_in_aw_ready ;  
   wire _axi4yank_auto_in_w_ready ;  
   wire _axi4yank_auto_in_b_valid ;  
   wire [3:0] _axi4yank_auto_in_b_bits_id ;  
   wire [1:0] _axi4yank_auto_in_b_bits_resp ;  
   wire [3:0] _axi4yank_auto_in_b_bits_echo_tl_state_size ;  
   wire [4:0] _axi4yank_auto_in_b_bits_echo_tl_state_source ;  
   wire _axi4yank_auto_in_ar_ready ;  
   wire _axi4yank_auto_in_r_valid ;  
   wire [3:0] _axi4yank_auto_in_r_bits_id ;  
   wire [63:0] _axi4yank_auto_in_r_bits_data ;  
   wire [1:0] _axi4yank_auto_in_r_bits_resp ;  
   wire [3:0] _axi4yank_auto_in_r_bits_echo_tl_state_size ;  
   wire [4:0] _axi4yank_auto_in_r_bits_echo_tl_state_source ;  
   wire _axi4yank_auto_in_r_bits_last ;  
   wire _axi4yank_auto_out_aw_valid ;  
   wire [3:0] _axi4yank_auto_out_aw_bits_id ;  
   wire [30:0] _axi4yank_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4yank_auto_out_aw_bits_len ;  
   wire [2:0] _axi4yank_auto_out_aw_bits_size ;  
   wire _axi4yank_auto_out_w_valid ;  
   wire [63:0] _axi4yank_auto_out_w_bits_data ;  
   wire [7:0] _axi4yank_auto_out_w_bits_strb ;  
   wire _axi4yank_auto_out_w_bits_last ;  
   wire _axi4yank_auto_out_b_ready ;  
   wire _axi4yank_auto_out_ar_valid ;  
   wire [3:0] _axi4yank_auto_out_ar_bits_id ;  
   wire [30:0] _axi4yank_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4yank_auto_out_ar_bits_len ;  
   wire [2:0] _axi4yank_auto_out_ar_bits_size ;  
   wire _axi4yank_auto_out_r_ready ;  
   wire _axi4buf_auto_in_aw_ready ;  
   wire _axi4buf_auto_in_w_ready ;  
   wire _axi4buf_auto_in_b_valid ;  
   wire [3:0] _axi4buf_auto_in_b_bits_id ;  
   wire [1:0] _axi4buf_auto_in_b_bits_resp ;  
   wire _axi4buf_auto_in_ar_ready ;  
   wire _axi4buf_auto_in_r_valid ;  
   wire [3:0] _axi4buf_auto_in_r_bits_id ;  
   wire [63:0] _axi4buf_auto_in_r_bits_data ;  
   wire [1:0] _axi4buf_auto_in_r_bits_resp ;  
   wire _axi4buf_auto_in_r_bits_last ;  
  AXI4Buffer axi4buf(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4buf_auto_in_aw_ready),.auto_in_aw_valid(_axi4yank_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4yank_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4yank_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4yank_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4yank_auto_out_aw_bits_size),.auto_in_w_ready(_axi4buf_auto_in_w_ready),.auto_in_w_valid(_axi4yank_auto_out_w_valid),.auto_in_w_bits_data(_axi4yank_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4yank_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4yank_auto_out_w_bits_last),.auto_in_b_ready(_axi4yank_auto_out_b_ready),.auto_in_b_valid(_axi4buf_auto_in_b_valid),.auto_in_b_bits_id(_axi4buf_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4buf_auto_in_b_bits_resp),.auto_in_ar_ready(_axi4buf_auto_in_ar_ready),.auto_in_ar_valid(_axi4yank_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4yank_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4yank_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4yank_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4yank_auto_out_ar_bits_size),.auto_in_r_ready(_axi4yank_auto_out_r_ready),.auto_in_r_valid(_axi4buf_auto_in_r_valid),.auto_in_r_bits_id(_axi4buf_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4buf_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4buf_auto_in_r_bits_resp),.auto_in_r_bits_last(_axi4buf_auto_in_r_bits_last),.auto_out_aw_ready(auto_axi4buf_out_aw_ready),.auto_out_aw_valid(auto_axi4buf_out_aw_valid),.auto_out_aw_bits_id(auto_axi4buf_out_aw_bits_id),.auto_out_aw_bits_addr(auto_axi4buf_out_aw_bits_addr),.auto_out_aw_bits_len(auto_axi4buf_out_aw_bits_len),.auto_out_aw_bits_size(auto_axi4buf_out_aw_bits_size),.auto_out_aw_bits_burst(auto_axi4buf_out_aw_bits_burst),.auto_out_aw_bits_lock(auto_axi4buf_out_aw_bits_lock),.auto_out_aw_bits_cache(auto_axi4buf_out_aw_bits_cache),.auto_out_aw_bits_prot(auto_axi4buf_out_aw_bits_prot),.auto_out_aw_bits_qos(auto_axi4buf_out_aw_bits_qos),.auto_out_w_ready(auto_axi4buf_out_w_ready),.auto_out_w_valid(auto_axi4buf_out_w_valid),.auto_out_w_bits_data(auto_axi4buf_out_w_bits_data),.auto_out_w_bits_strb(auto_axi4buf_out_w_bits_strb),.auto_out_w_bits_last(auto_axi4buf_out_w_bits_last),.auto_out_b_ready(auto_axi4buf_out_b_ready),.auto_out_b_valid(auto_axi4buf_out_b_valid),.auto_out_b_bits_id(auto_axi4buf_out_b_bits_id),.auto_out_b_bits_resp(auto_axi4buf_out_b_bits_resp),.auto_out_ar_ready(auto_axi4buf_out_ar_ready),.auto_out_ar_valid(auto_axi4buf_out_ar_valid),.auto_out_ar_bits_id(auto_axi4buf_out_ar_bits_id),.auto_out_ar_bits_addr(auto_axi4buf_out_ar_bits_addr),.auto_out_ar_bits_len(auto_axi4buf_out_ar_bits_len),.auto_out_ar_bits_size(auto_axi4buf_out_ar_bits_size),.auto_out_ar_bits_burst(auto_axi4buf_out_ar_bits_burst),.auto_out_ar_bits_lock(auto_axi4buf_out_ar_bits_lock),.auto_out_ar_bits_cache(auto_axi4buf_out_ar_bits_cache),.auto_out_ar_bits_prot(auto_axi4buf_out_ar_bits_prot),.auto_out_ar_bits_qos(auto_axi4buf_out_ar_bits_qos),.auto_out_r_ready(auto_axi4buf_out_r_ready),.auto_out_r_valid(auto_axi4buf_out_r_valid),.auto_out_r_bits_id(auto_axi4buf_out_r_bits_id),.auto_out_r_bits_data(auto_axi4buf_out_r_bits_data),.auto_out_r_bits_resp(auto_axi4buf_out_r_bits_resp),.auto_out_r_bits_last(auto_axi4buf_out_r_bits_last)); 
  AXI4UserYanker axi4yank(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4yank_auto_in_aw_ready),.auto_in_aw_valid(_axi4deint_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4deint_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4deint_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4deint_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4deint_auto_out_aw_bits_size),.auto_in_aw_bits_echo_tl_state_size(_axi4deint_auto_out_aw_bits_echo_tl_state_size),.auto_in_aw_bits_echo_tl_state_source(_axi4deint_auto_out_aw_bits_echo_tl_state_source),.auto_in_w_ready(_axi4yank_auto_in_w_ready),.auto_in_w_valid(_axi4deint_auto_out_w_valid),.auto_in_w_bits_data(_axi4deint_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4deint_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4deint_auto_out_w_bits_last),.auto_in_b_ready(_axi4deint_auto_out_b_ready),.auto_in_b_valid(_axi4yank_auto_in_b_valid),.auto_in_b_bits_id(_axi4yank_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4yank_auto_in_b_bits_resp),.auto_in_b_bits_echo_tl_state_size(_axi4yank_auto_in_b_bits_echo_tl_state_size),.auto_in_b_bits_echo_tl_state_source(_axi4yank_auto_in_b_bits_echo_tl_state_source),.auto_in_ar_ready(_axi4yank_auto_in_ar_ready),.auto_in_ar_valid(_axi4deint_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4deint_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4deint_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4deint_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4deint_auto_out_ar_bits_size),.auto_in_ar_bits_echo_tl_state_size(_axi4deint_auto_out_ar_bits_echo_tl_state_size),.auto_in_ar_bits_echo_tl_state_source(_axi4deint_auto_out_ar_bits_echo_tl_state_source),.auto_in_r_ready(_axi4deint_auto_out_r_ready),.auto_in_r_valid(_axi4yank_auto_in_r_valid),.auto_in_r_bits_id(_axi4yank_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4yank_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4yank_auto_in_r_bits_resp),.auto_in_r_bits_echo_tl_state_size(_axi4yank_auto_in_r_bits_echo_tl_state_size),.auto_in_r_bits_echo_tl_state_source(_axi4yank_auto_in_r_bits_echo_tl_state_source),.auto_in_r_bits_last(_axi4yank_auto_in_r_bits_last),.auto_out_aw_ready(_axi4buf_auto_in_aw_ready),.auto_out_aw_valid(_axi4yank_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4yank_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4yank_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4yank_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4yank_auto_out_aw_bits_size),.auto_out_w_ready(_axi4buf_auto_in_w_ready),.auto_out_w_valid(_axi4yank_auto_out_w_valid),.auto_out_w_bits_data(_axi4yank_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4yank_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4yank_auto_out_w_bits_last),.auto_out_b_ready(_axi4yank_auto_out_b_ready),.auto_out_b_valid(_axi4buf_auto_in_b_valid),.auto_out_b_bits_id(_axi4buf_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4buf_auto_in_b_bits_resp),.auto_out_ar_ready(_axi4buf_auto_in_ar_ready),.auto_out_ar_valid(_axi4yank_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4yank_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4yank_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4yank_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4yank_auto_out_ar_bits_size),.auto_out_r_ready(_axi4yank_auto_out_r_ready),.auto_out_r_valid(_axi4buf_auto_in_r_valid),.auto_out_r_bits_id(_axi4buf_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4buf_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4buf_auto_in_r_bits_resp),.auto_out_r_bits_last(_axi4buf_auto_in_r_bits_last)); 
  AXI4Deinterleaver axi4deint(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4deint_auto_in_aw_ready),.auto_in_aw_valid(_axi4index_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4index_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4index_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4index_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4index_auto_out_aw_bits_size),.auto_in_aw_bits_echo_tl_state_size(_axi4index_auto_out_aw_bits_echo_tl_state_size),.auto_in_aw_bits_echo_tl_state_source(_axi4index_auto_out_aw_bits_echo_tl_state_source),.auto_in_w_ready(_axi4deint_auto_in_w_ready),.auto_in_w_valid(_axi4index_auto_out_w_valid),.auto_in_w_bits_data(_axi4index_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4index_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4index_auto_out_w_bits_last),.auto_in_b_ready(_axi4index_auto_out_b_ready),.auto_in_b_valid(_axi4deint_auto_in_b_valid),.auto_in_b_bits_id(_axi4deint_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4deint_auto_in_b_bits_resp),.auto_in_b_bits_echo_tl_state_size(_axi4deint_auto_in_b_bits_echo_tl_state_size),.auto_in_b_bits_echo_tl_state_source(_axi4deint_auto_in_b_bits_echo_tl_state_source),.auto_in_ar_ready(_axi4deint_auto_in_ar_ready),.auto_in_ar_valid(_axi4index_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4index_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4index_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4index_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4index_auto_out_ar_bits_size),.auto_in_ar_bits_echo_tl_state_size(_axi4index_auto_out_ar_bits_echo_tl_state_size),.auto_in_ar_bits_echo_tl_state_source(_axi4index_auto_out_ar_bits_echo_tl_state_source),.auto_in_r_ready(_axi4index_auto_out_r_ready),.auto_in_r_valid(_axi4deint_auto_in_r_valid),.auto_in_r_bits_id(_axi4deint_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4deint_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4deint_auto_in_r_bits_resp),.auto_in_r_bits_echo_tl_state_size(_axi4deint_auto_in_r_bits_echo_tl_state_size),.auto_in_r_bits_echo_tl_state_source(_axi4deint_auto_in_r_bits_echo_tl_state_source),.auto_in_r_bits_last(_axi4deint_auto_in_r_bits_last),.auto_out_aw_ready(_axi4yank_auto_in_aw_ready),.auto_out_aw_valid(_axi4deint_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4deint_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4deint_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4deint_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4deint_auto_out_aw_bits_size),.auto_out_aw_bits_echo_tl_state_size(_axi4deint_auto_out_aw_bits_echo_tl_state_size),.auto_out_aw_bits_echo_tl_state_source(_axi4deint_auto_out_aw_bits_echo_tl_state_source),.auto_out_w_ready(_axi4yank_auto_in_w_ready),.auto_out_w_valid(_axi4deint_auto_out_w_valid),.auto_out_w_bits_data(_axi4deint_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4deint_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4deint_auto_out_w_bits_last),.auto_out_b_ready(_axi4deint_auto_out_b_ready),.auto_out_b_valid(_axi4yank_auto_in_b_valid),.auto_out_b_bits_id(_axi4yank_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4yank_auto_in_b_bits_resp),.auto_out_b_bits_echo_tl_state_size(_axi4yank_auto_in_b_bits_echo_tl_state_size),.auto_out_b_bits_echo_tl_state_source(_axi4yank_auto_in_b_bits_echo_tl_state_source),.auto_out_ar_ready(_axi4yank_auto_in_ar_ready),.auto_out_ar_valid(_axi4deint_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4deint_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4deint_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4deint_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4deint_auto_out_ar_bits_size),.auto_out_ar_bits_echo_tl_state_size(_axi4deint_auto_out_ar_bits_echo_tl_state_size),.auto_out_ar_bits_echo_tl_state_source(_axi4deint_auto_out_ar_bits_echo_tl_state_source),.auto_out_r_ready(_axi4deint_auto_out_r_ready),.auto_out_r_valid(_axi4yank_auto_in_r_valid),.auto_out_r_bits_id(_axi4yank_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4yank_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4yank_auto_in_r_bits_resp),.auto_out_r_bits_echo_tl_state_size(_axi4yank_auto_in_r_bits_echo_tl_state_size),.auto_out_r_bits_echo_tl_state_source(_axi4yank_auto_in_r_bits_echo_tl_state_source),.auto_out_r_bits_last(_axi4yank_auto_in_r_bits_last)); 
  AXI4IdIndexer axi4index(.auto_in_aw_ready(_axi4index_auto_in_aw_ready),.auto_in_aw_valid(_tl2axi4_auto_out_aw_valid),.auto_in_aw_bits_id(_tl2axi4_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_tl2axi4_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_tl2axi4_auto_out_aw_bits_len),.auto_in_aw_bits_size(_tl2axi4_auto_out_aw_bits_size),.auto_in_aw_bits_echo_tl_state_size(_tl2axi4_auto_out_aw_bits_echo_tl_state_size),.auto_in_aw_bits_echo_tl_state_source(_tl2axi4_auto_out_aw_bits_echo_tl_state_source),.auto_in_w_ready(_axi4index_auto_in_w_ready),.auto_in_w_valid(_tl2axi4_auto_out_w_valid),.auto_in_w_bits_data(_tl2axi4_auto_out_w_bits_data),.auto_in_w_bits_strb(_tl2axi4_auto_out_w_bits_strb),.auto_in_w_bits_last(_tl2axi4_auto_out_w_bits_last),.auto_in_b_ready(_tl2axi4_auto_out_b_ready),.auto_in_b_valid(_axi4index_auto_in_b_valid),.auto_in_b_bits_id(_axi4index_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4index_auto_in_b_bits_resp),.auto_in_b_bits_echo_tl_state_size(_axi4index_auto_in_b_bits_echo_tl_state_size),.auto_in_b_bits_echo_tl_state_source(_axi4index_auto_in_b_bits_echo_tl_state_source),.auto_in_ar_ready(_axi4index_auto_in_ar_ready),.auto_in_ar_valid(_tl2axi4_auto_out_ar_valid),.auto_in_ar_bits_id(_tl2axi4_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_tl2axi4_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_tl2axi4_auto_out_ar_bits_len),.auto_in_ar_bits_size(_tl2axi4_auto_out_ar_bits_size),.auto_in_ar_bits_echo_tl_state_size(_tl2axi4_auto_out_ar_bits_echo_tl_state_size),.auto_in_ar_bits_echo_tl_state_source(_tl2axi4_auto_out_ar_bits_echo_tl_state_source),.auto_in_r_ready(_tl2axi4_auto_out_r_ready),.auto_in_r_valid(_axi4index_auto_in_r_valid),.auto_in_r_bits_id(_axi4index_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4index_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4index_auto_in_r_bits_resp),.auto_in_r_bits_echo_tl_state_size(_axi4index_auto_in_r_bits_echo_tl_state_size),.auto_in_r_bits_echo_tl_state_source(_axi4index_auto_in_r_bits_echo_tl_state_source),.auto_in_r_bits_last(_axi4index_auto_in_r_bits_last),.auto_out_aw_ready(_axi4deint_auto_in_aw_ready),.auto_out_aw_valid(_axi4index_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4index_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4index_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4index_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4index_auto_out_aw_bits_size),.auto_out_aw_bits_echo_tl_state_size(_axi4index_auto_out_aw_bits_echo_tl_state_size),.auto_out_aw_bits_echo_tl_state_source(_axi4index_auto_out_aw_bits_echo_tl_state_source),.auto_out_w_ready(_axi4deint_auto_in_w_ready),.auto_out_w_valid(_axi4index_auto_out_w_valid),.auto_out_w_bits_data(_axi4index_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4index_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4index_auto_out_w_bits_last),.auto_out_b_ready(_axi4index_auto_out_b_ready),.auto_out_b_valid(_axi4deint_auto_in_b_valid),.auto_out_b_bits_id(_axi4deint_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4deint_auto_in_b_bits_resp),.auto_out_b_bits_echo_tl_state_size(_axi4deint_auto_in_b_bits_echo_tl_state_size),.auto_out_b_bits_echo_tl_state_source(_axi4deint_auto_in_b_bits_echo_tl_state_source),.auto_out_ar_ready(_axi4deint_auto_in_ar_ready),.auto_out_ar_valid(_axi4index_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4index_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4index_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4index_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4index_auto_out_ar_bits_size),.auto_out_ar_bits_echo_tl_state_size(_axi4index_auto_out_ar_bits_echo_tl_state_size),.auto_out_ar_bits_echo_tl_state_source(_axi4index_auto_out_ar_bits_echo_tl_state_source),.auto_out_r_ready(_axi4index_auto_out_r_ready),.auto_out_r_valid(_axi4deint_auto_in_r_valid),.auto_out_r_bits_id(_axi4deint_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4deint_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4deint_auto_in_r_bits_resp),.auto_out_r_bits_echo_tl_state_size(_axi4deint_auto_in_r_bits_echo_tl_state_size),.auto_out_r_bits_echo_tl_state_source(_axi4deint_auto_in_r_bits_echo_tl_state_source),.auto_out_r_bits_last(_axi4deint_auto_in_r_bits_last)); 
  TLToAXI4 tl2axi4(.clock(clock),.reset(reset),.auto_in_a_ready(auto_tl_in_a_ready),.auto_in_a_valid(auto_tl_in_a_valid),.auto_in_a_bits_opcode(auto_tl_in_a_bits_opcode),.auto_in_a_bits_param(auto_tl_in_a_bits_param),.auto_in_a_bits_size(auto_tl_in_a_bits_size),.auto_in_a_bits_source(auto_tl_in_a_bits_source),.auto_in_a_bits_address(auto_tl_in_a_bits_address),.auto_in_a_bits_mask(auto_tl_in_a_bits_mask),.auto_in_a_bits_data(auto_tl_in_a_bits_data),.auto_in_a_bits_corrupt(auto_tl_in_a_bits_corrupt),.auto_in_d_ready(auto_tl_in_d_ready),.auto_in_d_valid(auto_tl_in_d_valid),.auto_in_d_bits_opcode(auto_tl_in_d_bits_opcode),.auto_in_d_bits_size(auto_tl_in_d_bits_size),.auto_in_d_bits_source(auto_tl_in_d_bits_source),.auto_in_d_bits_denied(auto_tl_in_d_bits_denied),.auto_in_d_bits_data(auto_tl_in_d_bits_data),.auto_in_d_bits_corrupt(auto_tl_in_d_bits_corrupt),.auto_out_aw_ready(_axi4index_auto_in_aw_ready),.auto_out_aw_valid(_tl2axi4_auto_out_aw_valid),.auto_out_aw_bits_id(_tl2axi4_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_tl2axi4_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_tl2axi4_auto_out_aw_bits_len),.auto_out_aw_bits_size(_tl2axi4_auto_out_aw_bits_size),.auto_out_aw_bits_echo_tl_state_size(_tl2axi4_auto_out_aw_bits_echo_tl_state_size),.auto_out_aw_bits_echo_tl_state_source(_tl2axi4_auto_out_aw_bits_echo_tl_state_source),.auto_out_w_ready(_axi4index_auto_in_w_ready),.auto_out_w_valid(_tl2axi4_auto_out_w_valid),.auto_out_w_bits_data(_tl2axi4_auto_out_w_bits_data),.auto_out_w_bits_strb(_tl2axi4_auto_out_w_bits_strb),.auto_out_w_bits_last(_tl2axi4_auto_out_w_bits_last),.auto_out_b_ready(_tl2axi4_auto_out_b_ready),.auto_out_b_valid(_axi4index_auto_in_b_valid),.auto_out_b_bits_id(_axi4index_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4index_auto_in_b_bits_resp),.auto_out_b_bits_echo_tl_state_size(_axi4index_auto_in_b_bits_echo_tl_state_size),.auto_out_b_bits_echo_tl_state_source(_axi4index_auto_in_b_bits_echo_tl_state_source),.auto_out_ar_ready(_axi4index_auto_in_ar_ready),.auto_out_ar_valid(_tl2axi4_auto_out_ar_valid),.auto_out_ar_bits_id(_tl2axi4_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_tl2axi4_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_tl2axi4_auto_out_ar_bits_len),.auto_out_ar_bits_size(_tl2axi4_auto_out_ar_bits_size),.auto_out_ar_bits_echo_tl_state_size(_tl2axi4_auto_out_ar_bits_echo_tl_state_size),.auto_out_ar_bits_echo_tl_state_source(_tl2axi4_auto_out_ar_bits_echo_tl_state_source),.auto_out_r_ready(_tl2axi4_auto_out_r_ready),.auto_out_r_valid(_axi4index_auto_in_r_valid),.auto_out_r_bits_id(_axi4index_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4index_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4index_auto_in_r_bits_resp),.auto_out_r_bits_echo_tl_state_size(_axi4index_auto_in_r_bits_echo_tl_state_size),.auto_out_r_bits_echo_tl_state_source(_axi4index_auto_in_r_bits_echo_tl_state_source),.auto_out_r_bits_last(_axi4index_auto_in_r_bits_last)); 
endmodule
 
module SystemBus (
  input auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_ready,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_valid,
  output [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_id,
  output [30:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_addr,
  output [7:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_len,
  output [2:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_size,
  output [1:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_burst,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_lock,
  output [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_cache,
  output [2:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_prot,
  output [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_qos,
  input auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_ready,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_valid,
  output [63:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_data,
  output [7:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_strb,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_last,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_ready,
  input auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_valid,
  input [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_bits_id,
  input [1:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_bits_resp,
  input auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_ready,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_valid,
  output [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_id,
  output [30:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_addr,
  output [7:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_len,
  output [2:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_size,
  output [1:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_burst,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_lock,
  output [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_cache,
  output [2:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_prot,
  output [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_qos,
  output auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_ready,
  input auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_valid,
  input [3:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_id,
  input [63:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_data,
  input [1:0] auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_resp,
  input auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_last,
  output auto_coupler_from_tile_tl_master_clock_xing_in_a_ready,
  input auto_coupler_from_tile_tl_master_clock_xing_in_a_valid,
  input [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode,
  input [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param,
  input [3:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size,
  input [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source,
  input [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address,
  input [7:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask,
  input [63:0] auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data,
  input auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt,
  input auto_coupler_from_tile_tl_master_clock_xing_in_b_ready,
  output auto_coupler_from_tile_tl_master_clock_xing_in_b_valid,
  output [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param,
  output [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address,
  output auto_coupler_from_tile_tl_master_clock_xing_in_c_ready,
  input auto_coupler_from_tile_tl_master_clock_xing_in_c_valid,
  input [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode,
  input [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param,
  input [3:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size,
  input [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source,
  input [31:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address,
  input [63:0] auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data,
  input auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_corrupt,
  input auto_coupler_from_tile_tl_master_clock_xing_in_d_ready,
  output auto_coupler_from_tile_tl_master_clock_xing_in_d_valid,
  output [2:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode,
  output [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param,
  output [3:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size,
  output [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source,
  output [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink,
  output auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied,
  output [63:0] auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data,
  output auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt,
  input auto_coupler_from_tile_tl_master_clock_xing_in_e_valid,
  input [1:0] auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink,
  input auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready,
  output auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid,
  output [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode,
  output [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param,
  output [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size,
  output [4:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source,
  output [31:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address,
  output [7:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask,
  output [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data,
  output auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_corrupt,
  output auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready,
  input auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid,
  input [1:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param,
  input [31:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address,
  input auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready,
  output auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid,
  output [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode,
  output [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param,
  output [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size,
  output [4:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source,
  output [31:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address,
  output [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data,
  output auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_corrupt,
  output auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready,
  input auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid,
  input [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode,
  input [1:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param,
  input [2:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size,
  input [4:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source,
  input [1:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink,
  input auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied,
  input [63:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data,
  input auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt,
  output auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid,
  output [1:0] auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink,
  output auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready,
  input auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid,
  input [2:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode,
  input [2:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param,
  input [3:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size,
  input [3:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source,
  input [31:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address,
  input [7:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask,
  input [63:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data,
  input auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt,
  input auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready,
  output auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid,
  output [2:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode,
  output [1:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param,
  output [3:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size,
  output [3:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source,
  output [1:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink,
  output auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied,
  output [63:0] auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data,
  output auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt,
  input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready,
  output auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid,
  output [2:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode,
  output [2:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param,
  output [3:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size,
  output [4:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source,
  output [27:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address,
  output [7:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask,
  output [63:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data,
  output auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt,
  output auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready,
  input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid,
  input [2:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode,
  input [1:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param,
  input [3:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size,
  input [4:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source,
  input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink,
  input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied,
  input [63:0] auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data,
  input auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt,
  output auto_fixedClockNode_out_1_clock,
  output auto_fixedClockNode_out_1_reset,
  output auto_fixedClockNode_out_0_clock,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock,
  input auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset,
  output auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock,
  output auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset,
  output auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock,
  output auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset,
  output auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock,
  output auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset,
  output auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock,
  output auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset,
  output auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock,
  output auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset) ; 
   wire _coupler_to_port_named_mmio_port_axi4_auto_tl_in_a_ready ;  
   wire _coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_valid ;  
   wire [2:0] _coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_opcode ;  
   wire [3:0] _coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_size ;  
   wire [4:0] _coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_source ;  
   wire _coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_denied ;  
   wire [63:0] _coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_data ;  
   wire _coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_corrupt ;  
   wire _fixer_auto_out_1_a_valid ;  
   wire [2:0] _fixer_auto_out_1_a_bits_opcode ;  
   wire [2:0] _fixer_auto_out_1_a_bits_param ;  
   wire [3:0] _fixer_auto_out_1_a_bits_size ;  
   wire [1:0] _fixer_auto_out_1_a_bits_source ;  
   wire [31:0] _fixer_auto_out_1_a_bits_address ;  
   wire [7:0] _fixer_auto_out_1_a_bits_mask ;  
   wire [63:0] _fixer_auto_out_1_a_bits_data ;  
   wire _fixer_auto_out_1_a_bits_corrupt ;  
   wire _fixer_auto_out_1_b_ready ;  
   wire _fixer_auto_out_1_c_valid ;  
   wire [2:0] _fixer_auto_out_1_c_bits_opcode ;  
   wire [2:0] _fixer_auto_out_1_c_bits_param ;  
   wire [3:0] _fixer_auto_out_1_c_bits_size ;  
   wire [1:0] _fixer_auto_out_1_c_bits_source ;  
   wire [31:0] _fixer_auto_out_1_c_bits_address ;  
   wire [63:0] _fixer_auto_out_1_c_bits_data ;  
   wire _fixer_auto_out_1_c_bits_corrupt ;  
   wire _fixer_auto_out_1_d_ready ;  
   wire _fixer_auto_out_1_e_valid ;  
   wire [1:0] _fixer_auto_out_1_e_bits_sink ;  
   wire _fixer_auto_out_0_a_valid ;  
   wire [2:0] _fixer_auto_out_0_a_bits_opcode ;  
   wire [2:0] _fixer_auto_out_0_a_bits_param ;  
   wire [3:0] _fixer_auto_out_0_a_bits_size ;  
   wire [3:0] _fixer_auto_out_0_a_bits_source ;  
   wire [31:0] _fixer_auto_out_0_a_bits_address ;  
   wire [7:0] _fixer_auto_out_0_a_bits_mask ;  
   wire [63:0] _fixer_auto_out_0_a_bits_data ;  
   wire _fixer_auto_out_0_a_bits_corrupt ;  
   wire _fixer_auto_out_0_d_ready ;  
   wire _system_bus_xbar_auto_in_1_a_ready ;  
   wire _system_bus_xbar_auto_in_1_b_valid ;  
   wire [1:0] _system_bus_xbar_auto_in_1_b_bits_param ;  
   wire [31:0] _system_bus_xbar_auto_in_1_b_bits_address ;  
   wire _system_bus_xbar_auto_in_1_c_ready ;  
   wire _system_bus_xbar_auto_in_1_d_valid ;  
   wire [2:0] _system_bus_xbar_auto_in_1_d_bits_opcode ;  
   wire [1:0] _system_bus_xbar_auto_in_1_d_bits_param ;  
   wire [3:0] _system_bus_xbar_auto_in_1_d_bits_size ;  
   wire [1:0] _system_bus_xbar_auto_in_1_d_bits_source ;  
   wire [1:0] _system_bus_xbar_auto_in_1_d_bits_sink ;  
   wire _system_bus_xbar_auto_in_1_d_bits_denied ;  
   wire [63:0] _system_bus_xbar_auto_in_1_d_bits_data ;  
   wire _system_bus_xbar_auto_in_1_d_bits_corrupt ;  
   wire _system_bus_xbar_auto_in_0_a_ready ;  
   wire _system_bus_xbar_auto_in_0_d_valid ;  
   wire [2:0] _system_bus_xbar_auto_in_0_d_bits_opcode ;  
   wire [1:0] _system_bus_xbar_auto_in_0_d_bits_param ;  
   wire [3:0] _system_bus_xbar_auto_in_0_d_bits_size ;  
   wire [3:0] _system_bus_xbar_auto_in_0_d_bits_source ;  
   wire [1:0] _system_bus_xbar_auto_in_0_d_bits_sink ;  
   wire _system_bus_xbar_auto_in_0_d_bits_denied ;  
   wire [63:0] _system_bus_xbar_auto_in_0_d_bits_data ;  
   wire _system_bus_xbar_auto_in_0_d_bits_corrupt ;  
   wire _system_bus_xbar_auto_out_2_a_valid ;  
   wire [2:0] _system_bus_xbar_auto_out_2_a_bits_opcode ;  
   wire [2:0] _system_bus_xbar_auto_out_2_a_bits_param ;  
   wire [3:0] _system_bus_xbar_auto_out_2_a_bits_size ;  
   wire [4:0] _system_bus_xbar_auto_out_2_a_bits_source ;  
   wire [30:0] _system_bus_xbar_auto_out_2_a_bits_address ;  
   wire [7:0] _system_bus_xbar_auto_out_2_a_bits_mask ;  
   wire [63:0] _system_bus_xbar_auto_out_2_a_bits_data ;  
   wire _system_bus_xbar_auto_out_2_a_bits_corrupt ;  
   wire _system_bus_xbar_auto_out_2_d_ready ;  
   wire _fixedClockNode_auto_out_0_clock ;  
   wire _fixedClockNode_auto_out_0_reset ;  
  FixedClockBroadcast fixedClockNode(.auto_in_clock(auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock),.auto_in_reset(auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset),.auto_out_2_clock(auto_fixedClockNode_out_1_clock),.auto_out_2_reset(auto_fixedClockNode_out_1_reset),.auto_out_1_clock(auto_fixedClockNode_out_0_clock),.auto_out_0_clock(_fixedClockNode_auto_out_0_clock),.auto_out_0_reset(_fixedClockNode_auto_out_0_reset)); 
  TLXbar system_bus_xbar(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_in_1_a_ready(_system_bus_xbar_auto_in_1_a_ready),.auto_in_1_a_valid(_fixer_auto_out_1_a_valid),.auto_in_1_a_bits_opcode(_fixer_auto_out_1_a_bits_opcode),.auto_in_1_a_bits_param(_fixer_auto_out_1_a_bits_param),.auto_in_1_a_bits_size(_fixer_auto_out_1_a_bits_size),.auto_in_1_a_bits_source(_fixer_auto_out_1_a_bits_source),.auto_in_1_a_bits_address(_fixer_auto_out_1_a_bits_address),.auto_in_1_a_bits_mask(_fixer_auto_out_1_a_bits_mask),.auto_in_1_a_bits_data(_fixer_auto_out_1_a_bits_data),.auto_in_1_a_bits_corrupt(_fixer_auto_out_1_a_bits_corrupt),.auto_in_1_b_ready(_fixer_auto_out_1_b_ready),.auto_in_1_b_valid(_system_bus_xbar_auto_in_1_b_valid),.auto_in_1_b_bits_param(_system_bus_xbar_auto_in_1_b_bits_param),.auto_in_1_b_bits_address(_system_bus_xbar_auto_in_1_b_bits_address),.auto_in_1_c_ready(_system_bus_xbar_auto_in_1_c_ready),.auto_in_1_c_valid(_fixer_auto_out_1_c_valid),.auto_in_1_c_bits_opcode(_fixer_auto_out_1_c_bits_opcode),.auto_in_1_c_bits_param(_fixer_auto_out_1_c_bits_param),.auto_in_1_c_bits_size(_fixer_auto_out_1_c_bits_size),.auto_in_1_c_bits_source(_fixer_auto_out_1_c_bits_source),.auto_in_1_c_bits_address(_fixer_auto_out_1_c_bits_address),.auto_in_1_c_bits_data(_fixer_auto_out_1_c_bits_data),.auto_in_1_c_bits_corrupt(_fixer_auto_out_1_c_bits_corrupt),.auto_in_1_d_ready(_fixer_auto_out_1_d_ready),.auto_in_1_d_valid(_system_bus_xbar_auto_in_1_d_valid),.auto_in_1_d_bits_opcode(_system_bus_xbar_auto_in_1_d_bits_opcode),.auto_in_1_d_bits_param(_system_bus_xbar_auto_in_1_d_bits_param),.auto_in_1_d_bits_size(_system_bus_xbar_auto_in_1_d_bits_size),.auto_in_1_d_bits_source(_system_bus_xbar_auto_in_1_d_bits_source),.auto_in_1_d_bits_sink(_system_bus_xbar_auto_in_1_d_bits_sink),.auto_in_1_d_bits_denied(_system_bus_xbar_auto_in_1_d_bits_denied),.auto_in_1_d_bits_data(_system_bus_xbar_auto_in_1_d_bits_data),.auto_in_1_d_bits_corrupt(_system_bus_xbar_auto_in_1_d_bits_corrupt),.auto_in_1_e_valid(_fixer_auto_out_1_e_valid),.auto_in_1_e_bits_sink(_fixer_auto_out_1_e_bits_sink),.auto_in_0_a_ready(_system_bus_xbar_auto_in_0_a_ready),.auto_in_0_a_valid(_fixer_auto_out_0_a_valid),.auto_in_0_a_bits_opcode(_fixer_auto_out_0_a_bits_opcode),.auto_in_0_a_bits_param(_fixer_auto_out_0_a_bits_param),.auto_in_0_a_bits_size(_fixer_auto_out_0_a_bits_size),.auto_in_0_a_bits_source(_fixer_auto_out_0_a_bits_source),.auto_in_0_a_bits_address(_fixer_auto_out_0_a_bits_address),.auto_in_0_a_bits_mask(_fixer_auto_out_0_a_bits_mask),.auto_in_0_a_bits_data(_fixer_auto_out_0_a_bits_data),.auto_in_0_a_bits_corrupt(_fixer_auto_out_0_a_bits_corrupt),.auto_in_0_d_ready(_fixer_auto_out_0_d_ready),.auto_in_0_d_valid(_system_bus_xbar_auto_in_0_d_valid),.auto_in_0_d_bits_opcode(_system_bus_xbar_auto_in_0_d_bits_opcode),.auto_in_0_d_bits_param(_system_bus_xbar_auto_in_0_d_bits_param),.auto_in_0_d_bits_size(_system_bus_xbar_auto_in_0_d_bits_size),.auto_in_0_d_bits_source(_system_bus_xbar_auto_in_0_d_bits_source),.auto_in_0_d_bits_sink(_system_bus_xbar_auto_in_0_d_bits_sink),.auto_in_0_d_bits_denied(_system_bus_xbar_auto_in_0_d_bits_denied),.auto_in_0_d_bits_data(_system_bus_xbar_auto_in_0_d_bits_data),.auto_in_0_d_bits_corrupt(_system_bus_xbar_auto_in_0_d_bits_corrupt),.auto_out_2_a_ready(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_a_ready),.auto_out_2_a_valid(_system_bus_xbar_auto_out_2_a_valid),.auto_out_2_a_bits_opcode(_system_bus_xbar_auto_out_2_a_bits_opcode),.auto_out_2_a_bits_param(_system_bus_xbar_auto_out_2_a_bits_param),.auto_out_2_a_bits_size(_system_bus_xbar_auto_out_2_a_bits_size),.auto_out_2_a_bits_source(_system_bus_xbar_auto_out_2_a_bits_source),.auto_out_2_a_bits_address(_system_bus_xbar_auto_out_2_a_bits_address),.auto_out_2_a_bits_mask(_system_bus_xbar_auto_out_2_a_bits_mask),.auto_out_2_a_bits_data(_system_bus_xbar_auto_out_2_a_bits_data),.auto_out_2_a_bits_corrupt(_system_bus_xbar_auto_out_2_a_bits_corrupt),.auto_out_2_d_ready(_system_bus_xbar_auto_out_2_d_ready),.auto_out_2_d_valid(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_valid),.auto_out_2_d_bits_opcode(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_opcode),.auto_out_2_d_bits_size(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_size),.auto_out_2_d_bits_source(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_source),.auto_out_2_d_bits_denied(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_denied),.auto_out_2_d_bits_data(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_data),.auto_out_2_d_bits_corrupt(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_corrupt),.auto_out_1_a_ready(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready),.auto_out_1_a_valid(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid),.auto_out_1_a_bits_opcode(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode),.auto_out_1_a_bits_param(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param),.auto_out_1_a_bits_size(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size),.auto_out_1_a_bits_source(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source),.auto_out_1_a_bits_address(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address),.auto_out_1_a_bits_mask(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask),.auto_out_1_a_bits_data(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data),.auto_out_1_a_bits_corrupt(auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_corrupt),.auto_out_1_b_ready(auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready),.auto_out_1_b_valid(auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid),.auto_out_1_b_bits_param(auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param),.auto_out_1_b_bits_address(auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address),.auto_out_1_c_ready(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready),.auto_out_1_c_valid(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid),.auto_out_1_c_bits_opcode(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode),.auto_out_1_c_bits_param(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param),.auto_out_1_c_bits_size(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size),.auto_out_1_c_bits_source(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source),.auto_out_1_c_bits_address(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address),.auto_out_1_c_bits_data(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data),.auto_out_1_c_bits_corrupt(auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_corrupt),.auto_out_1_d_ready(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready),.auto_out_1_d_valid(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid),.auto_out_1_d_bits_opcode(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode),.auto_out_1_d_bits_param(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param),.auto_out_1_d_bits_size(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size),.auto_out_1_d_bits_source(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source),.auto_out_1_d_bits_sink(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink),.auto_out_1_d_bits_denied(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied),.auto_out_1_d_bits_data(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data),.auto_out_1_d_bits_corrupt(auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt),.auto_out_1_e_valid(auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid),.auto_out_1_e_bits_sink(auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink),.auto_out_0_a_ready(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready),.auto_out_0_a_valid(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid),.auto_out_0_a_bits_opcode(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode),.auto_out_0_a_bits_param(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param),.auto_out_0_a_bits_size(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size),.auto_out_0_a_bits_source(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source),.auto_out_0_a_bits_address(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address),.auto_out_0_a_bits_mask(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask),.auto_out_0_a_bits_data(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data),.auto_out_0_a_bits_corrupt(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt),.auto_out_0_d_ready(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready),.auto_out_0_d_valid(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid),.auto_out_0_d_bits_opcode(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode),.auto_out_0_d_bits_param(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param),.auto_out_0_d_bits_size(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size),.auto_out_0_d_bits_source(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source),.auto_out_0_d_bits_sink(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink),.auto_out_0_d_bits_denied(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied),.auto_out_0_d_bits_data(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data),.auto_out_0_d_bits_corrupt(auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt)); 
  TLFIFOFixer fixer(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_in_1_a_ready(auto_coupler_from_tile_tl_master_clock_xing_in_a_ready),.auto_in_1_a_valid(auto_coupler_from_tile_tl_master_clock_xing_in_a_valid),.auto_in_1_a_bits_opcode(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode),.auto_in_1_a_bits_param(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param),.auto_in_1_a_bits_size(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size),.auto_in_1_a_bits_source(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source),.auto_in_1_a_bits_address(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address),.auto_in_1_a_bits_mask(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask),.auto_in_1_a_bits_data(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data),.auto_in_1_a_bits_corrupt(auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt),.auto_in_1_b_ready(auto_coupler_from_tile_tl_master_clock_xing_in_b_ready),.auto_in_1_b_valid(auto_coupler_from_tile_tl_master_clock_xing_in_b_valid),.auto_in_1_b_bits_param(auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param),.auto_in_1_b_bits_address(auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address),.auto_in_1_c_ready(auto_coupler_from_tile_tl_master_clock_xing_in_c_ready),.auto_in_1_c_valid(auto_coupler_from_tile_tl_master_clock_xing_in_c_valid),.auto_in_1_c_bits_opcode(auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode),.auto_in_1_c_bits_param(auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param),.auto_in_1_c_bits_size(auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size),.auto_in_1_c_bits_source(auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source),.auto_in_1_c_bits_address(auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address),.auto_in_1_c_bits_data(auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data),.auto_in_1_c_bits_corrupt(auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_corrupt),.auto_in_1_d_ready(auto_coupler_from_tile_tl_master_clock_xing_in_d_ready),.auto_in_1_d_valid(auto_coupler_from_tile_tl_master_clock_xing_in_d_valid),.auto_in_1_d_bits_opcode(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode),.auto_in_1_d_bits_param(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param),.auto_in_1_d_bits_size(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size),.auto_in_1_d_bits_source(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source),.auto_in_1_d_bits_sink(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink),.auto_in_1_d_bits_denied(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied),.auto_in_1_d_bits_data(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data),.auto_in_1_d_bits_corrupt(auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt),.auto_in_1_e_valid(auto_coupler_from_tile_tl_master_clock_xing_in_e_valid),.auto_in_1_e_bits_sink(auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink),.auto_in_0_a_ready(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready),.auto_in_0_a_valid(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid),.auto_in_0_a_bits_opcode(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode),.auto_in_0_a_bits_param(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param),.auto_in_0_a_bits_size(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size),.auto_in_0_a_bits_source(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source),.auto_in_0_a_bits_address(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address),.auto_in_0_a_bits_mask(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask),.auto_in_0_a_bits_data(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data),.auto_in_0_a_bits_corrupt(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt),.auto_in_0_d_ready(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready),.auto_in_0_d_valid(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid),.auto_in_0_d_bits_opcode(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode),.auto_in_0_d_bits_param(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param),.auto_in_0_d_bits_size(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size),.auto_in_0_d_bits_source(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source),.auto_in_0_d_bits_sink(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink),.auto_in_0_d_bits_denied(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied),.auto_in_0_d_bits_data(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data),.auto_in_0_d_bits_corrupt(auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt),.auto_out_1_a_ready(_system_bus_xbar_auto_in_1_a_ready),.auto_out_1_a_valid(_fixer_auto_out_1_a_valid),.auto_out_1_a_bits_opcode(_fixer_auto_out_1_a_bits_opcode),.auto_out_1_a_bits_param(_fixer_auto_out_1_a_bits_param),.auto_out_1_a_bits_size(_fixer_auto_out_1_a_bits_size),.auto_out_1_a_bits_source(_fixer_auto_out_1_a_bits_source),.auto_out_1_a_bits_address(_fixer_auto_out_1_a_bits_address),.auto_out_1_a_bits_mask(_fixer_auto_out_1_a_bits_mask),.auto_out_1_a_bits_data(_fixer_auto_out_1_a_bits_data),.auto_out_1_a_bits_corrupt(_fixer_auto_out_1_a_bits_corrupt),.auto_out_1_b_ready(_fixer_auto_out_1_b_ready),.auto_out_1_b_valid(_system_bus_xbar_auto_in_1_b_valid),.auto_out_1_b_bits_param(_system_bus_xbar_auto_in_1_b_bits_param),.auto_out_1_b_bits_address(_system_bus_xbar_auto_in_1_b_bits_address),.auto_out_1_c_ready(_system_bus_xbar_auto_in_1_c_ready),.auto_out_1_c_valid(_fixer_auto_out_1_c_valid),.auto_out_1_c_bits_opcode(_fixer_auto_out_1_c_bits_opcode),.auto_out_1_c_bits_param(_fixer_auto_out_1_c_bits_param),.auto_out_1_c_bits_size(_fixer_auto_out_1_c_bits_size),.auto_out_1_c_bits_source(_fixer_auto_out_1_c_bits_source),.auto_out_1_c_bits_address(_fixer_auto_out_1_c_bits_address),.auto_out_1_c_bits_data(_fixer_auto_out_1_c_bits_data),.auto_out_1_c_bits_corrupt(_fixer_auto_out_1_c_bits_corrupt),.auto_out_1_d_ready(_fixer_auto_out_1_d_ready),.auto_out_1_d_valid(_system_bus_xbar_auto_in_1_d_valid),.auto_out_1_d_bits_opcode(_system_bus_xbar_auto_in_1_d_bits_opcode),.auto_out_1_d_bits_param(_system_bus_xbar_auto_in_1_d_bits_param),.auto_out_1_d_bits_size(_system_bus_xbar_auto_in_1_d_bits_size),.auto_out_1_d_bits_source(_system_bus_xbar_auto_in_1_d_bits_source),.auto_out_1_d_bits_sink(_system_bus_xbar_auto_in_1_d_bits_sink),.auto_out_1_d_bits_denied(_system_bus_xbar_auto_in_1_d_bits_denied),.auto_out_1_d_bits_data(_system_bus_xbar_auto_in_1_d_bits_data),.auto_out_1_d_bits_corrupt(_system_bus_xbar_auto_in_1_d_bits_corrupt),.auto_out_1_e_valid(_fixer_auto_out_1_e_valid),.auto_out_1_e_bits_sink(_fixer_auto_out_1_e_bits_sink),.auto_out_0_a_ready(_system_bus_xbar_auto_in_0_a_ready),.auto_out_0_a_valid(_fixer_auto_out_0_a_valid),.auto_out_0_a_bits_opcode(_fixer_auto_out_0_a_bits_opcode),.auto_out_0_a_bits_param(_fixer_auto_out_0_a_bits_param),.auto_out_0_a_bits_size(_fixer_auto_out_0_a_bits_size),.auto_out_0_a_bits_source(_fixer_auto_out_0_a_bits_source),.auto_out_0_a_bits_address(_fixer_auto_out_0_a_bits_address),.auto_out_0_a_bits_mask(_fixer_auto_out_0_a_bits_mask),.auto_out_0_a_bits_data(_fixer_auto_out_0_a_bits_data),.auto_out_0_a_bits_corrupt(_fixer_auto_out_0_a_bits_corrupt),.auto_out_0_d_ready(_fixer_auto_out_0_d_ready),.auto_out_0_d_valid(_system_bus_xbar_auto_in_0_d_valid),.auto_out_0_d_bits_opcode(_system_bus_xbar_auto_in_0_d_bits_opcode),.auto_out_0_d_bits_param(_system_bus_xbar_auto_in_0_d_bits_param),.auto_out_0_d_bits_size(_system_bus_xbar_auto_in_0_d_bits_size),.auto_out_0_d_bits_source(_system_bus_xbar_auto_in_0_d_bits_source),.auto_out_0_d_bits_sink(_system_bus_xbar_auto_in_0_d_bits_sink),.auto_out_0_d_bits_denied(_system_bus_xbar_auto_in_0_d_bits_denied),.auto_out_0_d_bits_data(_system_bus_xbar_auto_in_0_d_bits_data),.auto_out_0_d_bits_corrupt(_system_bus_xbar_auto_in_0_d_bits_corrupt)); 
  TLInterconnectCoupler_4 coupler_to_port_named_mmio_port_axi4(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_axi4buf_out_aw_ready(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_ready),.auto_axi4buf_out_aw_valid(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_valid),.auto_axi4buf_out_aw_bits_id(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_id),.auto_axi4buf_out_aw_bits_addr(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_addr),.auto_axi4buf_out_aw_bits_len(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_len),.auto_axi4buf_out_aw_bits_size(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_size),.auto_axi4buf_out_aw_bits_burst(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_burst),.auto_axi4buf_out_aw_bits_lock(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_lock),.auto_axi4buf_out_aw_bits_cache(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_cache),.auto_axi4buf_out_aw_bits_prot(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_prot),.auto_axi4buf_out_aw_bits_qos(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_qos),.auto_axi4buf_out_w_ready(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_ready),.auto_axi4buf_out_w_valid(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_valid),.auto_axi4buf_out_w_bits_data(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_data),.auto_axi4buf_out_w_bits_strb(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_strb),.auto_axi4buf_out_w_bits_last(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_last),.auto_axi4buf_out_b_ready(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_ready),.auto_axi4buf_out_b_valid(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_valid),.auto_axi4buf_out_b_bits_id(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_bits_id),.auto_axi4buf_out_b_bits_resp(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_bits_resp),.auto_axi4buf_out_ar_ready(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_ready),.auto_axi4buf_out_ar_valid(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_valid),.auto_axi4buf_out_ar_bits_id(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_id),.auto_axi4buf_out_ar_bits_addr(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_addr),.auto_axi4buf_out_ar_bits_len(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_len),.auto_axi4buf_out_ar_bits_size(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_size),.auto_axi4buf_out_ar_bits_burst(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_burst),.auto_axi4buf_out_ar_bits_lock(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_lock),.auto_axi4buf_out_ar_bits_cache(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_cache),.auto_axi4buf_out_ar_bits_prot(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_prot),.auto_axi4buf_out_ar_bits_qos(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_qos),.auto_axi4buf_out_r_ready(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_ready),.auto_axi4buf_out_r_valid(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_valid),.auto_axi4buf_out_r_bits_id(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_id),.auto_axi4buf_out_r_bits_data(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_data),.auto_axi4buf_out_r_bits_resp(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_resp),.auto_axi4buf_out_r_bits_last(auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_last),.auto_tl_in_a_ready(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_a_ready),.auto_tl_in_a_valid(_system_bus_xbar_auto_out_2_a_valid),.auto_tl_in_a_bits_opcode(_system_bus_xbar_auto_out_2_a_bits_opcode),.auto_tl_in_a_bits_param(_system_bus_xbar_auto_out_2_a_bits_param),.auto_tl_in_a_bits_size(_system_bus_xbar_auto_out_2_a_bits_size),.auto_tl_in_a_bits_source(_system_bus_xbar_auto_out_2_a_bits_source),.auto_tl_in_a_bits_address(_system_bus_xbar_auto_out_2_a_bits_address),.auto_tl_in_a_bits_mask(_system_bus_xbar_auto_out_2_a_bits_mask),.auto_tl_in_a_bits_data(_system_bus_xbar_auto_out_2_a_bits_data),.auto_tl_in_a_bits_corrupt(_system_bus_xbar_auto_out_2_a_bits_corrupt),.auto_tl_in_d_ready(_system_bus_xbar_auto_out_2_d_ready),.auto_tl_in_d_valid(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_valid),.auto_tl_in_d_bits_opcode(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_opcode),.auto_tl_in_d_bits_size(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_size),.auto_tl_in_d_bits_source(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_source),.auto_tl_in_d_bits_denied(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_denied),.auto_tl_in_d_bits_data(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_data),.auto_tl_in_d_bits_corrupt(_coupler_to_port_named_mmio_port_axi4_auto_tl_in_d_bits_corrupt)); 
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock; 
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset; 
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock; 
  assign auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset; 
  assign auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock; 
  assign auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset; 
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock; 
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset; 
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock; 
  assign auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset=auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset; 
endmodule
 
module PeripheryBus (
  input auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock,
  input auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset,
  output clock,
  output reset) ; 
  assign clock=auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock; 
  assign reset=auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset; 
endmodule
 
module TLMonitor_5 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [3:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [3:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [3:0] source ;  
   reg [31:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [3:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [15:0] inflight ;  
   reg [63:0] inflight_opcodes ;  
   reg [127:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [63:0] _a_opcode_lookup_T_1=inflight_opcodes>>{58'h0,io_in_d_bits_source,2'h0} ;  
   wire [15:0] _GEN_0={12'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [15:0] _GEN_2={12'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [15:0] inflight_1 ;  
   reg [127:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_bits_size<4'h7 ;  
   wire _GEN_6=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_7=_GEN_4&_GEN_5&_GEN_6 ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_9=io_in_a_bits_param>3'h2 ;  
   wire _GEN_10=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_11=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_13={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_14=_GEN_4&_GEN_13 ;  
   wire _GEN_15=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_16={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_17={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_18={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_19=io_in_a_bits_mask!=mask ;  
   wire _GEN_20=_GEN_4&(_GEN_14|_GEN_5&(_GEN_15|_GEN_16|_GEN_17|_GEN_6)|io_in_a_bits_size<4'h9&_GEN_18) ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_22=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_23=_GEN_4&io_in_a_bits_size<4'h4&(_GEN_15|_GEN_13|_GEN_16|_GEN_17) ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_26=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_27=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_28=io_in_d_bits_size<4'h3 ;  
   wire _GEN_29=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_30=io_in_d_bits_param==2'h2 ;  
   wire _GEN_31=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_32=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_33=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_35=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_36=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_37=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [127:0] _GEN_38={121'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [15:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 16'h1<<_GEN_0:16'h0 ;  
   wire _GEN_39=io_in_d_valid&d_first_1 ;  
   wire _GEN_40=_GEN_39&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_41=_GEN_40&same_cycle_resp&~reset ;  
   wire _GEN_42=_GEN_40&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_43={4'h0,io_in_d_bits_size} ;  
   wire _GEN_44=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [15:0] _GEN_45=inflight>>_GEN_0 ;  
   wire [15:0] _GEN_46=inflight>>_GEN_2 ;  
   wire [127:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_38 ;  
   wire [15:0] _GEN_47=inflight_1>>_GEN_2 ;  
   wire [127:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_38 ;  
  always @( posedge clock)
       begin 
         if (_GEN_8&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~(_GEN_14|_GEN_5&(_GEN_15|{io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0|_GEN_16|_GEN_17|_GEN_18|_GEN_6)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(_GEN_4&_GEN_14))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_45[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~reset&~(_GEN_46[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_43!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_40 ? 16'h1<<_GEN_2:16'h0)|a_set_wo_ready==16'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==16'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~(_GEN_47[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&_GEN_43!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==16'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_48={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_48 ;  
   wire [142:0] _GEN_49={136'h0,io_in_d_bits_source,3'h0} ;  
   wire [142:0] _d_opcodes_clr_T_5=143'hF<<{137'h0,io_in_d_bits_source,2'h0} ;  
   wire [130:0] _a_opcodes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{125'h0,io_in_a_bits_source,2'h0} ;  
   wire [142:0] _d_sizes_clr_T_5=143'hFF<<_GEN_49 ;  
   wire [131:0] _a_sizes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{125'h0,io_in_a_bits_source,3'h0} ;  
   wire [142:0] _d_sizes_clr_T_11=143'hFF<<_GEN_49 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_50=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_51=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=16'h0;
              inflight_opcodes <=64'h0;
              inflight_sizes <=128'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=16'h0;
              inflight_sizes_1 <=128'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? 16'h1<<_GEN_0:16'h0))&~(_GEN_50 ? 16'h1<<_GEN_2:16'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[63:0]:64'h0))&~(_GEN_50 ? _d_opcodes_clr_T_5[63:0]:64'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[127:0]:128'h0))&~(_GEN_50 ? _d_sizes_clr_T_5[127:0]:128'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_51 ? 16'h1<<_GEN_2:16'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_51 ? _d_sizes_clr_T_11[127:0]:128'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module ram_addr_2x32 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [31:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [31:0] W0_data) ; 
   reg [31:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:32'bx; 
endmodule
 
module Queue_22 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [3:0] io_enq_bits_source,
  input [31:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input [63:0] io_enq_bits_data,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [3:0] io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x3 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_2x4 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_addr_2x32 ram_address_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_address),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_address)); 
  ram_2x8 ram_mask_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_mask),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_mask)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_corrupt)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_23 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [1:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [3:0] io_enq_bits_source,
  input [1:0] io_enq_bits_sink,
  input io_enq_bits_denied,
  input [63:0] io_enq_bits_data,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [1:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [3:0] io_deq_bits_source,
  output [1:0] io_deq_bits_sink,
  output io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x2 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_2x4 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_2x2 ram_sink_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_sink),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_sink)); 
  ram_2x1 ram_denied_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_denied),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_denied)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_corrupt)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module TLBuffer_2 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [3:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [3:0] auto_in_d_bits_source,
  output [1:0] auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [3:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [3:0] auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   wire _nodeIn_d_q_io_deq_valid ;  
   wire [2:0] _nodeIn_d_q_io_deq_bits_opcode ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_param ;  
   wire [3:0] _nodeIn_d_q_io_deq_bits_size ;  
   wire [3:0] _nodeIn_d_q_io_deq_bits_source ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_sink ;  
   wire _nodeIn_d_q_io_deq_bits_denied ;  
   wire _nodeIn_d_q_io_deq_bits_corrupt ;  
   wire _nodeOut_a_q_io_enq_ready ;  
  TLMonitor_5 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_nodeOut_a_q_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(_nodeIn_d_q_io_deq_valid),.io_in_d_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_in_d_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_in_d_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_in_d_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_in_d_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_in_d_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_in_d_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  Queue_22 nodeOut_a_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_a_q_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_data(auto_in_a_bits_data),.io_enq_bits_corrupt(auto_in_a_bits_corrupt),.io_deq_ready(auto_out_a_ready),.io_deq_valid(auto_out_a_valid),.io_deq_bits_opcode(auto_out_a_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(auto_out_a_bits_size),.io_deq_bits_source(auto_out_a_bits_source),.io_deq_bits_address(auto_out_a_bits_address),.io_deq_bits_mask(auto_out_a_bits_mask),.io_deq_bits_data(auto_out_a_bits_data),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  Queue_23 nodeIn_d_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_d_ready),.io_enq_valid(auto_out_d_valid),.io_enq_bits_opcode(auto_out_d_bits_opcode),.io_enq_bits_param(auto_out_d_bits_param),.io_enq_bits_size(auto_out_d_bits_size),.io_enq_bits_source(auto_out_d_bits_source),.io_enq_bits_sink(auto_out_d_bits_sink),.io_enq_bits_denied(auto_out_d_bits_denied),.io_enq_bits_data(auto_out_d_bits_data),.io_enq_bits_corrupt(auto_out_d_bits_corrupt),.io_deq_ready(auto_in_d_ready),.io_deq_valid(_nodeIn_d_q_io_deq_valid),.io_deq_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_deq_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_deq_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_deq_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_deq_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_deq_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_deq_bits_data(auto_in_d_bits_data),.io_deq_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  assign auto_in_a_ready=_nodeOut_a_q_io_enq_ready; 
  assign auto_in_d_valid=_nodeIn_d_q_io_deq_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_q_io_deq_bits_opcode; 
  assign auto_in_d_bits_param=_nodeIn_d_q_io_deq_bits_param; 
  assign auto_in_d_bits_size=_nodeIn_d_q_io_deq_bits_size; 
  assign auto_in_d_bits_source=_nodeIn_d_q_io_deq_bits_source; 
  assign auto_in_d_bits_sink=_nodeIn_d_q_io_deq_bits_sink; 
  assign auto_in_d_bits_denied=_nodeIn_d_q_io_deq_bits_denied; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_q_io_deq_bits_corrupt; 
endmodule
 
module TLMonitor_6 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [3:0] io_in_a_bits_size,
  input [3:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [3:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [3:0] size ;  
   reg [3:0] source ;  
   reg [31:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [3:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [15:0] inflight ;  
   reg [63:0] inflight_opcodes ;  
   reg [127:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [63:0] _a_opcode_lookup_T_1=inflight_opcodes>>{58'h0,io_in_d_bits_source,2'h0} ;  
   wire [15:0] _GEN_0={12'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [15:0] _GEN_2={12'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [15:0] inflight_1 ;  
   reg [127:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_bits_size<4'h7 ;  
   wire _GEN_6=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_7=_GEN_4&_GEN_5&_GEN_6 ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_9=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_10=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_12={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_13=_GEN_4&_GEN_12 ;  
   wire _GEN_14=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_15={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_16={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_17={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_18=io_in_a_bits_mask!=mask ;  
   wire _GEN_19=_GEN_4&(_GEN_13|_GEN_5&(_GEN_14|_GEN_15|_GEN_16|_GEN_6)|io_in_a_bits_size<4'h9&_GEN_17) ;  
   wire _GEN_20=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_22=_GEN_4&io_in_a_bits_size<4'h4&(_GEN_14|_GEN_12|_GEN_15|_GEN_16) ;  
   wire _GEN_23=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_26=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_27=io_in_d_bits_size<4'h3 ;  
   wire _GEN_28=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_29=io_in_d_bits_param==2'h2 ;  
   wire _GEN_30=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_31=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_32=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_33=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_35=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_36=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [127:0] _GEN_37={121'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [15:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 16'h1<<_GEN_0:16'h0 ;  
   wire _GEN_38=io_in_d_valid&d_first_1 ;  
   wire _GEN_39=_GEN_38&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_40=_GEN_39&same_cycle_resp&~reset ;  
   wire _GEN_41=_GEN_39&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_42={4'h0,io_in_d_bits_size} ;  
   wire _GEN_43=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [15:0] _GEN_44=inflight>>_GEN_0 ;  
   wire [15:0] _GEN_45=inflight>>_GEN_2 ;  
   wire [127:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_37 ;  
   wire [15:0] _GEN_46=inflight_1>>_GEN_2 ;  
   wire [127:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_37 ;  
  always @( posedge clock)
       begin 
         if (_GEN_8&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(_GEN_13|_GEN_5&(_GEN_14|{io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0|_GEN_15|_GEN_16|_GEN_17|_GEN_6)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~(_GEN_4&_GEN_13))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_44[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&~reset&~(_GEN_45[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&_GEN_42!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_39 ? 16'h1<<_GEN_2:16'h0)|a_set_wo_ready==16'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 5 (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==16'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&~(_GEN_46[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&_GEN_42!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==16'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:151:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_47={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_47 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_47 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_47 ;  
   wire [142:0] _GEN_48={136'h0,io_in_d_bits_source,3'h0} ;  
   wire [142:0] _d_opcodes_clr_T_5=143'hF<<{137'h0,io_in_d_bits_source,2'h0} ;  
   wire [130:0] _a_opcodes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{125'h0,io_in_a_bits_source,2'h0} ;  
   wire [142:0] _d_sizes_clr_T_5=143'hFF<<_GEN_48 ;  
   wire [131:0] _a_sizes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{125'h0,io_in_a_bits_source,3'h0} ;  
   wire [142:0] _d_sizes_clr_T_11=143'hFF<<_GEN_48 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_49=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_50=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=16'h0;
              inflight_opcodes <=64'h0;
              inflight_sizes <=128'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=16'h0;
              inflight_sizes_1 <=128'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? 16'h1<<_GEN_0:16'h0))&~(_GEN_49 ? 16'h1<<_GEN_2:16'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[63:0]:64'h0))&~(_GEN_49 ? _d_opcodes_clr_T_5[63:0]:64'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[127:0]:128'h0))&~(_GEN_49 ? _d_sizes_clr_T_5[127:0]:128'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_50 ? 16'h1<<_GEN_2:16'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_50 ? _d_sizes_clr_T_11[127:0]:128'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLBuffer_3 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [3:0] auto_in_a_bits_size,
  input [3:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [3:0] auto_in_d_bits_source,
  output [1:0] auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [3:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [3:0] auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   wire _nodeIn_d_q_io_deq_valid ;  
   wire [2:0] _nodeIn_d_q_io_deq_bits_opcode ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_param ;  
   wire [3:0] _nodeIn_d_q_io_deq_bits_size ;  
   wire [3:0] _nodeIn_d_q_io_deq_bits_source ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_sink ;  
   wire _nodeIn_d_q_io_deq_bits_denied ;  
   wire _nodeIn_d_q_io_deq_bits_corrupt ;  
   wire _nodeOut_a_q_io_enq_ready ;  
  TLMonitor_6 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_nodeOut_a_q_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(_nodeIn_d_q_io_deq_valid),.io_in_d_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_in_d_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_in_d_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_in_d_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_in_d_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_in_d_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_in_d_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  Queue_22 nodeOut_a_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_a_q_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(3'h0),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_data(auto_in_a_bits_data),.io_enq_bits_corrupt(1'h0),.io_deq_ready(auto_out_a_ready),.io_deq_valid(auto_out_a_valid),.io_deq_bits_opcode(auto_out_a_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(auto_out_a_bits_size),.io_deq_bits_source(auto_out_a_bits_source),.io_deq_bits_address(auto_out_a_bits_address),.io_deq_bits_mask(auto_out_a_bits_mask),.io_deq_bits_data(auto_out_a_bits_data),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  Queue_23 nodeIn_d_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_d_ready),.io_enq_valid(auto_out_d_valid),.io_enq_bits_opcode(auto_out_d_bits_opcode),.io_enq_bits_param(auto_out_d_bits_param),.io_enq_bits_size(auto_out_d_bits_size),.io_enq_bits_source(auto_out_d_bits_source),.io_enq_bits_sink(auto_out_d_bits_sink),.io_enq_bits_denied(auto_out_d_bits_denied),.io_enq_bits_data(auto_out_d_bits_data),.io_enq_bits_corrupt(auto_out_d_bits_corrupt),.io_deq_ready(auto_in_d_ready),.io_deq_valid(_nodeIn_d_q_io_deq_valid),.io_deq_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_deq_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_deq_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_deq_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_deq_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_deq_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_deq_bits_data(auto_in_d_bits_data),.io_deq_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  assign auto_in_a_ready=_nodeOut_a_q_io_enq_ready; 
  assign auto_in_d_valid=_nodeIn_d_q_io_deq_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_q_io_deq_bits_opcode; 
  assign auto_in_d_bits_param=_nodeIn_d_q_io_deq_bits_param; 
  assign auto_in_d_bits_size=_nodeIn_d_q_io_deq_bits_size; 
  assign auto_in_d_bits_source=_nodeIn_d_q_io_deq_bits_source; 
  assign auto_in_d_bits_sink=_nodeIn_d_q_io_deq_bits_sink; 
  assign auto_in_d_bits_denied=_nodeIn_d_q_io_deq_bits_denied; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_q_io_deq_bits_corrupt; 
endmodule
 
module TLMonitor_7 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [3:0] io_in_a_bits_size,
  input [3:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [3:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [3:0] size ;  
   reg [3:0] source ;  
   reg [31:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [3:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [15:0] inflight ;  
   reg [63:0] inflight_opcodes ;  
   reg [127:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [63:0] _a_opcode_lookup_T_1=inflight_opcodes>>{58'h0,io_in_d_bits_source,2'h0} ;  
   wire [15:0] _GEN_0={12'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [15:0] _GEN_2={12'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [15:0] inflight_1 ;  
   reg [127:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_bits_size<4'h7 ;  
   wire _GEN_6=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_7=_GEN_4&_GEN_5&_GEN_6 ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_9=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_10=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_12={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_13=_GEN_4&_GEN_12 ;  
   wire _GEN_14=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_15={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_16={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_17={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_18=io_in_a_bits_mask!=mask ;  
   wire _GEN_19=_GEN_4&(_GEN_13|_GEN_5&(_GEN_14|_GEN_15|_GEN_16|_GEN_6)|io_in_a_bits_size<4'h9&_GEN_17) ;  
   wire _GEN_20=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_22=_GEN_4&io_in_a_bits_size<4'h4&(_GEN_14|_GEN_12|_GEN_15|_GEN_16) ;  
   wire _GEN_23=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_26=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_27=io_in_d_bits_size<4'h3 ;  
   wire _GEN_28=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_29=io_in_d_bits_param==2'h2 ;  
   wire _GEN_30=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_31=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_32=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_33=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_35=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_36=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [127:0] _GEN_37={121'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [15:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 16'h1<<_GEN_0:16'h0 ;  
   wire _GEN_38=io_in_d_valid&d_first_1 ;  
   wire _GEN_39=_GEN_38&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_40=_GEN_39&same_cycle_resp&~reset ;  
   wire _GEN_41=_GEN_39&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_42={4'h0,io_in_d_bits_size} ;  
   wire _GEN_43=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [15:0] _GEN_44=inflight>>_GEN_0 ;  
   wire [15:0] _GEN_45=inflight>>_GEN_2 ;  
   wire [127:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_37 ;  
   wire [15:0] _GEN_46=inflight_1>>_GEN_2 ;  
   wire [127:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_37 ;  
  always @( posedge clock)
       begin 
         if (_GEN_8&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(_GEN_13|_GEN_5&(_GEN_14|{io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0|_GEN_15|_GEN_16|_GEN_17|_GEN_6)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~(_GEN_4&_GEN_13))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_44[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&~reset&~(_GEN_45[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&_GEN_42!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_39 ? 16'h1<<_GEN_2:16'h0)|a_set_wo_ready==16'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 5 (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==16'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&~(_GEN_46[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&_GEN_42!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==16'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:152:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_47={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_47 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_47 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_47 ;  
   wire [142:0] _GEN_48={136'h0,io_in_d_bits_source,3'h0} ;  
   wire [142:0] _d_opcodes_clr_T_5=143'hF<<{137'h0,io_in_d_bits_source,2'h0} ;  
   wire [130:0] _a_opcodes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{125'h0,io_in_a_bits_source,2'h0} ;  
   wire [142:0] _d_sizes_clr_T_5=143'hFF<<_GEN_48 ;  
   wire [131:0] _a_sizes_set_T_1={127'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{125'h0,io_in_a_bits_source,3'h0} ;  
   wire [142:0] _d_sizes_clr_T_11=143'hFF<<_GEN_48 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_49=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_50=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=16'h0;
              inflight_opcodes <=64'h0;
              inflight_sizes <=128'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=16'h0;
              inflight_sizes_1 <=128'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? 16'h1<<_GEN_0:16'h0))&~(_GEN_49 ? 16'h1<<_GEN_2:16'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[63:0]:64'h0))&~(_GEN_49 ? _d_opcodes_clr_T_5[63:0]:64'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[127:0]:128'h0))&~(_GEN_49 ? _d_sizes_clr_T_5[127:0]:128'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_50 ? 16'h1<<_GEN_2:16'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_50 ? _d_sizes_clr_T_11[127:0]:128'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLFIFOFixer_2 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [3:0] auto_in_a_bits_size,
  input [3:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [3:0] auto_in_d_bits_size,
  output [3:0] auto_in_d_bits_source,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [3:0] auto_out_a_bits_size,
  output [3:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [3:0] auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   reg [8:0] a_first_counter ;  
   wire a_first=a_first_counter==9'h0 ;  
   reg [8:0] d_first_counter ;  
   reg flight_0 ;  
   reg flight_1 ;  
   reg flight_2 ;  
   reg flight_3 ;  
   reg flight_4 ;  
   reg flight_5 ;  
   reg flight_6 ;  
   reg flight_7 ;  
   reg flight_8 ;  
   reg flight_9 ;  
   reg flight_10 ;  
   reg flight_11 ;  
   reg flight_12 ;  
   reg flight_13 ;  
   reg flight_14 ;  
   reg flight_15 ;  
   reg stalls_id ;  
   reg stalls_id_1 ;  
   wire stall=~(auto_in_a_bits_source[3])&a_first&(flight_0|flight_1|flight_2|flight_3|flight_4|flight_5|flight_6|flight_7)&(auto_in_a_bits_address[31]|stalls_id!=~(auto_in_a_bits_address[31]))|auto_in_a_bits_source[3]&a_first&(flight_8|flight_9|flight_10|flight_11|flight_12|flight_13|flight_14|flight_15)&(auto_in_a_bits_address[31]|stalls_id_1!=~(auto_in_a_bits_address[31])) ;  
   wire nodeIn_a_ready=auto_out_a_ready&~stall ;  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<auto_in_a_bits_size ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<auto_out_d_bits_size ;  
   wire d_first_first=d_first_counter==9'h0 ;  
   wire _GEN=d_first_first&auto_out_d_bits_opcode!=3'h6&auto_in_d_ready&auto_out_d_valid ;  
   wire _stalls_id_T_4=nodeIn_a_ready&auto_in_a_valid ;  
   wire _GEN_0=a_first&_stalls_id_T_4 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              flight_0 <=1'h0;
              flight_1 <=1'h0;
              flight_2 <=1'h0;
              flight_3 <=1'h0;
              flight_4 <=1'h0;
              flight_5 <=1'h0;
              flight_6 <=1'h0;
              flight_7 <=1'h0;
              flight_8 <=1'h0;
              flight_9 <=1'h0;
              flight_10 <=1'h0;
              flight_11 <=1'h0;
              flight_12 <=1'h0;
              flight_13 <=1'h0;
              flight_14 <=1'h0;
              flight_15 <=1'h0;
            end 
          else 
            begin 
              if (_stalls_id_T_4)
                 begin 
                   if (a_first)
                      a_first_counter <=auto_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                    else 
                      a_first_counter <=a_first_counter-9'h1;
                 end 
              if (auto_in_d_ready&auto_out_d_valid)
                 begin 
                   if (d_first_first)
                      d_first_counter <=auto_out_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                    else 
                      d_first_counter <=d_first_counter-9'h1;
                 end 
              flight_0 <=~(_GEN&auto_out_d_bits_source==4'h0)&(_GEN_0&auto_in_a_bits_source==4'h0|flight_0);
              flight_1 <=~(_GEN&auto_out_d_bits_source==4'h1)&(_GEN_0&auto_in_a_bits_source==4'h1|flight_1);
              flight_2 <=~(_GEN&auto_out_d_bits_source==4'h2)&(_GEN_0&auto_in_a_bits_source==4'h2|flight_2);
              flight_3 <=~(_GEN&auto_out_d_bits_source==4'h3)&(_GEN_0&auto_in_a_bits_source==4'h3|flight_3);
              flight_4 <=~(_GEN&auto_out_d_bits_source==4'h4)&(_GEN_0&auto_in_a_bits_source==4'h4|flight_4);
              flight_5 <=~(_GEN&auto_out_d_bits_source==4'h5)&(_GEN_0&auto_in_a_bits_source==4'h5|flight_5);
              flight_6 <=~(_GEN&auto_out_d_bits_source==4'h6)&(_GEN_0&auto_in_a_bits_source==4'h6|flight_6);
              flight_7 <=~(_GEN&auto_out_d_bits_source==4'h7)&(_GEN_0&auto_in_a_bits_source==4'h7|flight_7);
              flight_8 <=~(_GEN&auto_out_d_bits_source==4'h8)&(_GEN_0&auto_in_a_bits_source==4'h8|flight_8);
              flight_9 <=~(_GEN&auto_out_d_bits_source==4'h9)&(_GEN_0&auto_in_a_bits_source==4'h9|flight_9);
              flight_10 <=~(_GEN&auto_out_d_bits_source==4'hA)&(_GEN_0&auto_in_a_bits_source==4'hA|flight_10);
              flight_11 <=~(_GEN&auto_out_d_bits_source==4'hB)&(_GEN_0&auto_in_a_bits_source==4'hB|flight_11);
              flight_12 <=~(_GEN&auto_out_d_bits_source==4'hC)&(_GEN_0&auto_in_a_bits_source==4'hC|flight_12);
              flight_13 <=~(_GEN&auto_out_d_bits_source==4'hD)&(_GEN_0&auto_in_a_bits_source==4'hD|flight_13);
              flight_14 <=~(_GEN&auto_out_d_bits_source==4'hE)&(_GEN_0&auto_in_a_bits_source==4'hE|flight_14);
              flight_15 <=~(_GEN&(&auto_out_d_bits_source))&(_GEN_0&(&auto_in_a_bits_source)|flight_15);
            end 
         if (_stalls_id_T_4&~(auto_in_a_bits_source[3]))
            stalls_id <=~(auto_in_a_bits_address[31]);
         if (_stalls_id_T_4&auto_in_a_bits_source[3])
            stalls_id_1 <=~(auto_in_a_bits_address[31]);
       end
  
  TLMonitor_7 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_out_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_param(auto_out_d_bits_param),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source),.io_in_d_bits_sink(auto_out_d_bits_sink),.io_in_d_bits_denied(auto_out_d_bits_denied),.io_in_d_bits_corrupt(auto_out_d_bits_corrupt)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_d_valid=auto_out_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source; 
  assign auto_in_d_bits_denied=auto_out_d_bits_denied; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign auto_out_a_valid=auto_in_a_valid&~stall; 
  assign auto_out_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_a_bits_size=auto_in_a_bits_size; 
  assign auto_out_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_d_ready=auto_in_d_ready; 
endmodule
 
module Queue_26 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input io_enq_bits_id,
  input [63:0] io_enq_bits_data,
  input [1:0] io_enq_bits_resp,
  input io_enq_bits_last,
  input io_deq_ready,
  output io_deq_valid,
  output io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0] io_deq_bits_resp,
  output io_deq_bits_last) ; 
   reg ram_last ;  
   reg [1:0] ram_resp ;  
   reg [63:0] ram_data ;  
   reg ram_id ;  
   reg full ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire do_enq=~(~full&io_deq_ready)&~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_last <=io_enq_bits_last;
              ram_resp <=io_enq_bits_resp;
              ram_data <=io_enq_bits_data;
              ram_id <=io_enq_bits_id;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(full&io_deq_ready&io_deq_valid_0)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_id=full ? ram_id:io_enq_bits_id; 
  assign io_deq_bits_data=full ? ram_data:io_enq_bits_data; 
  assign io_deq_bits_resp=full ? ram_resp:io_enq_bits_resp; 
  assign io_deq_bits_last=full ? ram_last:io_enq_bits_last; 
endmodule
 
module Queue_27 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input io_enq_bits_id,
  input [1:0] io_enq_bits_resp,
  input io_deq_ready,
  output io_deq_valid,
  output io_deq_bits_id,
  output [1:0] io_deq_bits_resp) ; 
   reg [1:0] ram_resp ;  
   reg ram_id ;  
   reg full ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire do_enq=~(~full&io_deq_ready)&~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_resp <=io_enq_bits_resp;
              ram_id <=io_enq_bits_id;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(full&io_deq_ready&io_deq_valid_0)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_id=full ? ram_id:io_enq_bits_id; 
  assign io_deq_bits_resp=full ? ram_resp:io_enq_bits_resp; 
endmodule
 
module AXI4ToTL (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_last,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [3:0] auto_out_a_bits_size,
  output [3:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [3:0] auto_out_d_bits_size,
  input [3:0] auto_out_d_bits_source,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   wire w_out_ready ;  
   wire _q_b_deq_q_io_enq_ready ;  
   wire _q_b_deq_q_io_deq_valid ;  
   wire _q_b_deq_q_io_deq_bits_id ;  
   wire _nodeIn_r_deq_q_io_enq_ready ;  
   wire [22:0] _r_size1_T_1={7'h0,auto_in_ar_bits_len,8'hFF}<<auto_in_ar_bits_size ;  
   wire [13:0] _GEN=~(_r_size1_T_1[22:9]) ;  
   wire [7:0] r_size_hi=_r_size1_T_1[22:15]&{1'h1,_GEN[13:7]} ;  
   wire [6:0] _r_size_T_6=r_size_hi[7:1]|_r_size1_T_1[14:8]&_GEN[6:0] ;  
   wire [2:0] _r_size_T_8=_r_size_T_6[6:4]|_r_size_T_6[2:0] ;  
   wire _r_size_T_10=_r_size_T_8[2]|_r_size_T_8[0] ;  
   wire [3:0] r_size={|r_size_hi,|(_r_size_T_6[6:3]),|(_r_size_T_8[2:1]),_r_size_T_10} ;  
   wire [31:0] r_addr=r_size<4'hD&{auto_in_ar_bits_addr[31:14],~(auto_in_ar_bits_addr[13:12])}==20'h0|r_size<4'h7&(auto_in_ar_bits_addr[31:12]==20'h0|{auto_in_ar_bits_addr[31:17],~(auto_in_ar_bits_addr[16])}==16'h0|{auto_in_ar_bits_addr[31:26],auto_in_ar_bits_addr[25:16]^10'h200}==16'h0|{auto_in_ar_bits_addr[31:28],~(auto_in_ar_bits_addr[27:26])}==6'h0|{auto_in_ar_bits_addr[31],~(auto_in_ar_bits_addr[30:29])}==3'h0|auto_in_ar_bits_addr[31:28]==4'h8) ? auto_in_ar_bits_addr:{29'h600,auto_in_ar_bits_addr[2:0]} ;  
   reg [2:0] r_count_0 ;  
   reg [2:0] r_count_1 ;  
   wire _r_out_bits_a_mask_T=r_size>4'h2 ;  
   wire [1:0] _GEN_0={|(_r_size_T_8[2:1]),_r_size_T_10} ;  
   wire r_out_bits_a_mask_size=_GEN_0==2'h2 ;  
   wire r_out_bits_a_mask_acc=_r_out_bits_a_mask_T|r_out_bits_a_mask_size&~(r_addr[2]) ;  
   wire r_out_bits_a_mask_acc_1=_r_out_bits_a_mask_T|r_out_bits_a_mask_size&r_addr[2] ;  
   wire r_out_bits_a_mask_size_1=_GEN_0==2'h1 ;  
   wire r_out_bits_a_mask_eq_2=~(r_addr[2])&~(r_addr[1]) ;  
   wire r_out_bits_a_mask_acc_2=r_out_bits_a_mask_acc|r_out_bits_a_mask_size_1&r_out_bits_a_mask_eq_2 ;  
   wire r_out_bits_a_mask_eq_3=~(r_addr[2])&r_addr[1] ;  
   wire r_out_bits_a_mask_acc_3=r_out_bits_a_mask_acc|r_out_bits_a_mask_size_1&r_out_bits_a_mask_eq_3 ;  
   wire r_out_bits_a_mask_eq_4=r_addr[2]&~(r_addr[1]) ;  
   wire r_out_bits_a_mask_acc_4=r_out_bits_a_mask_acc_1|r_out_bits_a_mask_size_1&r_out_bits_a_mask_eq_4 ;  
   wire r_out_bits_a_mask_eq_5=r_addr[2]&r_addr[1] ;  
   wire r_out_bits_a_mask_acc_5=r_out_bits_a_mask_acc_1|r_out_bits_a_mask_size_1&r_out_bits_a_mask_eq_5 ;  
   wire [22:0] _w_size1_T_1={7'h0,auto_in_aw_bits_len,8'hFF}<<auto_in_aw_bits_size ;  
   wire [13:0] _GEN_1=~(_w_size1_T_1[22:9]) ;  
   wire [7:0] w_size_hi=_w_size1_T_1[22:15]&{1'h1,_GEN_1[13:7]} ;  
   wire [6:0] _w_size_T_6=w_size_hi[7:1]|_w_size1_T_1[14:8]&_GEN_1[6:0] ;  
   wire [2:0] _w_size_T_8=_w_size_T_6[6:4]|_w_size_T_6[2:0] ;  
   wire _w_size_T_10=_w_size_T_8[2]|_w_size_T_8[0] ;  
   wire [3:0] w_size={|w_size_hi,|(_w_size_T_6[6:3]),|(_w_size_T_8[2:1]),_w_size_T_10} ;  
   reg [2:0] w_count_0 ;  
   reg [2:0] w_count_1 ;  
   wire nodeIn_aw_ready=w_out_ready&auto_in_w_valid&auto_in_w_bits_last ;  
   wire w_out_valid=auto_in_aw_valid&auto_in_w_valid ;  
   reg [7:0] beatsLeft ;  
   wire idle=beatsLeft==8'h0 ;  
   wire [1:0] readys_valid={w_out_valid,auto_in_ar_valid} ;  
   reg [1:0] readys_mask ;  
   wire [1:0] _readys_filter_T_1=readys_valid&~readys_mask ;  
   wire [1:0] readys_readys=~({readys_mask[1],_readys_filter_T_1[1]|readys_mask[0]}&({_readys_filter_T_1[0],w_out_valid}|_readys_filter_T_1)) ;  
   wire winner_0=readys_readys[0]&auto_in_ar_valid ;  
   wire winner_1=readys_readys[1]&w_out_valid ;  
   wire _nodeOut_a_valid_T=auto_in_ar_valid|w_out_valid ;  
   wire [29:0] _GEN_2=30'h7FFF<<{26'h0,|r_size_hi,|(_r_size_T_6[6:3]),|(_r_size_T_8[2:1]),_r_size_T_10} ;  
   wire [29:0] _GEN_3=30'h7FFF<<{26'h0,|w_size_hi,|(_w_size_T_6[6:3]),|(_w_size_T_8[2:1]),_w_size_T_10} ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~auto_in_ar_valid|_r_size1_T_1[22:8]==~(_GEN_2[14:0])))
            begin 
              if (1)$display("Assertion failed\n    at ToTL.scala:108 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n");
              if (1)$display("");
            end 
         if (~reset&~(~auto_in_aw_valid|_w_size1_T_1[22:8]==~(_GEN_3[14:0])))
            begin 
              if (1)$display("Assertion failed\n    at ToTL.scala:144 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n");
              if (1)$display("");
            end 
         if (~reset&~(~auto_in_aw_valid|auto_in_aw_bits_len==8'h0|auto_in_aw_bits_size==3'h3))
            begin 
              if (1)$display("Assertion failed\n    at ToTL.scala:145 assert (!in.aw.valid || in.aw.bits.len === 0.U || in.aw.bits.size === log2Ceil(beatBytes).U) // because aligned\n");
              if (1)$display("");
            end 
         if (~reset&~(~winner_0|~winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_nodeOut_a_valid_T|winner_0|winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg state_0 ;  
   reg state_1 ;  
   wire muxState_0=idle ? winner_0:state_0 ;  
   wire muxState_1=idle ? winner_1:state_1 ;  
   wire r_out_ready=auto_out_a_ready&(idle ? readys_readys[0]:state_0) ;  
  assign w_out_ready=auto_out_a_ready&(idle ? readys_readys[1]:state_1); 
   wire nodeOut_a_valid=idle ? _nodeOut_a_valid_T:state_0&auto_in_ar_valid|state_1&w_out_valid ;  
   wire [1:0] d_resp={auto_out_d_bits_denied|auto_out_d_bits_corrupt,1'h0} ;  
   wire [26:0] _d_last_beats1_decode_T_1=27'hFFF<<auto_out_d_bits_size ;  
   wire [8:0] d_last_beats1=auto_out_d_bits_opcode[0] ? ~(_d_last_beats1_decode_T_1[11:3]):9'h0 ;  
   reg [8:0] d_last_counter ;  
   wire nodeOut_d_ready=auto_out_d_bits_opcode[0] ? _nodeIn_r_deq_q_io_enq_ready:_q_b_deq_q_io_enq_ready ;  
   reg [2:0] b_count_0 ;  
   reg [2:0] b_count_1 ;  
   wire b_allow=(_q_b_deq_q_io_deq_bits_id ? b_count_1:b_count_0)!=(_q_b_deq_q_io_deq_bits_id ? w_count_1:w_count_0) ;  
   wire nodeIn_b_valid=_q_b_deq_q_io_deq_valid&b_allow ;  
   wire [1:0] _readys_mask_T=readys_readys&readys_valid ;  
   wire _GEN_4=r_out_ready&auto_in_ar_valid ;  
   wire _GEN_5=nodeIn_aw_ready&auto_in_aw_valid ;  
   wire latch=idle&auto_out_a_ready ;  
   wire _GEN_6=auto_in_b_ready&nodeIn_b_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              r_count_0 <=3'h0;
              r_count_1 <=3'h0;
              w_count_0 <=3'h0;
              w_count_1 <=3'h0;
              beatsLeft <=8'h0;
              readys_mask <=2'h3;
              state_0 <=1'h0;
              state_1 <=1'h0;
              d_last_counter <=9'h0;
              b_count_0 <=3'h0;
              b_count_1 <=3'h0;
            end 
          else 
            begin 
              if (_GEN_4&~auto_in_ar_bits_id)
                 r_count_0 <=r_count_0+3'h1;
              if (_GEN_4&auto_in_ar_bits_id)
                 r_count_1 <=r_count_1+3'h1;
              if (_GEN_5&~auto_in_aw_bits_id)
                 w_count_0 <=w_count_0+3'h1;
              if (_GEN_5&auto_in_aw_bits_id)
                 w_count_1 <=w_count_1+3'h1;
              if (latch)
                 beatsLeft <=winner_1 ? auto_in_aw_bits_len:8'h0;
               else 
                 beatsLeft <=beatsLeft-{7'h0,auto_out_a_ready&nodeOut_a_valid};
              if (latch&(|readys_valid))
                 readys_mask <=_readys_mask_T|{_readys_mask_T[0],1'h0};
              if (idle)
                 begin 
                   state_0 <=winner_0;
                   state_1 <=winner_1;
                 end 
              if (nodeOut_d_ready&auto_out_d_valid)
                 begin 
                   if (d_last_counter==9'h0)
                      d_last_counter <=d_last_beats1;
                    else 
                      d_last_counter <=d_last_counter-9'h1;
                 end 
              if (_GEN_6&~_q_b_deq_q_io_deq_bits_id)
                 b_count_0 <=b_count_0+3'h1;
              if (_GEN_6&_q_b_deq_q_io_deq_bits_id)
                 b_count_1 <=b_count_1+3'h1;
            end 
       end
  
  Queue_26 nodeIn_r_deq_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeIn_r_deq_q_io_enq_ready),.io_enq_valid(auto_out_d_valid&auto_out_d_bits_opcode[0]),.io_enq_bits_id(auto_out_d_bits_source[3]),.io_enq_bits_data(auto_out_d_bits_data),.io_enq_bits_resp(d_resp),.io_enq_bits_last(d_last_counter==9'h1|d_last_beats1==9'h0),.io_deq_ready(auto_in_r_ready),.io_deq_valid(auto_in_r_valid),.io_deq_bits_id(auto_in_r_bits_id),.io_deq_bits_data(auto_in_r_bits_data),.io_deq_bits_resp(auto_in_r_bits_resp),.io_deq_bits_last(auto_in_r_bits_last)); 
  Queue_27 q_b_deq_q(.clock(clock),.reset(reset),.io_enq_ready(_q_b_deq_q_io_enq_ready),.io_enq_valid(auto_out_d_valid&~(auto_out_d_bits_opcode[0])),.io_enq_bits_id(auto_out_d_bits_source[3]),.io_enq_bits_resp(d_resp),.io_deq_ready(auto_in_b_ready&b_allow),.io_deq_valid(_q_b_deq_q_io_deq_valid),.io_deq_bits_id(_q_b_deq_q_io_deq_bits_id),.io_deq_bits_resp(auto_in_b_bits_resp)); 
  assign auto_in_aw_ready=nodeIn_aw_ready; 
  assign auto_in_w_ready=w_out_ready&auto_in_aw_valid; 
  assign auto_in_b_valid=nodeIn_b_valid; 
  assign auto_in_b_bits_id=_q_b_deq_q_io_deq_bits_id; 
  assign auto_in_ar_ready=r_out_ready; 
  assign auto_out_a_valid=nodeOut_a_valid; 
  assign auto_out_a_bits_opcode={muxState_0,1'h0,muxState_1}; 
  assign auto_out_a_bits_size=(muxState_0 ? r_size:4'h0)|(muxState_1 ? w_size:4'h0); 
  assign auto_out_a_bits_source=(muxState_0 ? {auto_in_ar_bits_id,auto_in_ar_bits_id ? r_count_1[1:0]:r_count_0[1:0],1'h0}:4'h0)|(muxState_1 ? {auto_in_aw_bits_id,auto_in_aw_bits_id ? w_count_1[1:0]:w_count_0[1:0],1'h1}:4'h0); 
  assign auto_out_a_bits_address=(muxState_0 ? r_addr:32'h0)|(muxState_1 ? (w_size<4'hD&{auto_in_aw_bits_addr[31:14],~(auto_in_aw_bits_addr[13:12])}==20'h0|w_size<4'h7&(auto_in_aw_bits_addr[31:12]==20'h0|{auto_in_aw_bits_addr[31:26],auto_in_aw_bits_addr[25:16]^10'h200}==16'h0|{auto_in_aw_bits_addr[31:28],~(auto_in_aw_bits_addr[27:26])}==6'h0|auto_in_aw_bits_addr[31:28]==4'h8)|w_size<4'h9&{auto_in_aw_bits_addr[31],~(auto_in_aw_bits_addr[30:29])}==3'h0 ? auto_in_aw_bits_addr:{29'h600,auto_in_aw_bits_addr[2:0]}):32'h0); 
  assign auto_out_a_bits_mask=(muxState_0 ? {r_out_bits_a_mask_acc_5|r_out_bits_a_mask_eq_5&r_addr[0],r_out_bits_a_mask_acc_5|r_out_bits_a_mask_eq_5&~(r_addr[0]),r_out_bits_a_mask_acc_4|r_out_bits_a_mask_eq_4&r_addr[0],r_out_bits_a_mask_acc_4|r_out_bits_a_mask_eq_4&~(r_addr[0]),r_out_bits_a_mask_acc_3|r_out_bits_a_mask_eq_3&r_addr[0],r_out_bits_a_mask_acc_3|r_out_bits_a_mask_eq_3&~(r_addr[0]),r_out_bits_a_mask_acc_2|r_out_bits_a_mask_eq_2&r_addr[0],r_out_bits_a_mask_acc_2|r_out_bits_a_mask_eq_2&~(r_addr[0])}:8'h0)|(muxState_1 ? auto_in_w_bits_strb:8'h0); 
  assign auto_out_a_bits_data=muxState_1 ? auto_in_w_bits_data:64'h0; 
  assign auto_out_d_ready=nodeOut_d_ready; 
endmodule
 
module ram_4x8 (
  input [1:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [7:0] R0_data,
  input [1:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [7:0] W0_data) ; 
   reg [7:0] Memory[0:3] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:8'bx; 
endmodule
 
module Queue_28 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [6:0] io_enq_bits_extra_id,
  input io_enq_bits_real_last,
  input io_deq_ready,
  output io_deq_valid,
  output [6:0] io_deq_bits_extra_id,
  output io_deq_bits_real_last) ; 
   wire [7:0] _ram_ext_R0_data ;  
   reg [1:0] enq_ptr_value ;  
   reg [1:0] deq_ptr_value ;  
   reg maybe_full ;  
   wire ptr_match=enq_ptr_value==deq_ptr_value ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              enq_ptr_value <=2'h0;
              deq_ptr_value <=2'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 enq_ptr_value <=enq_ptr_value+2'h1;
              if (do_deq)
                 deq_ptr_value <=deq_ptr_value+2'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_4x8 ram_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(_ram_ext_R0_data),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data({io_enq_bits_real_last,io_enq_bits_extra_id})); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
  assign io_deq_bits_extra_id=_ram_ext_R0_data[6:0]; 
  assign io_deq_bits_real_last=_ram_ext_R0_data[7]; 
endmodule
 
module AXI4UserYanker_1 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [6:0] auto_in_aw_bits_echo_extra_id,
  input auto_in_aw_bits_echo_real_last,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output [6:0] auto_in_b_bits_echo_extra_id,
  output auto_in_b_bits_echo_real_last,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [6:0] auto_in_ar_bits_echo_extra_id,
  input auto_in_ar_bits_echo_real_last,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output [6:0] auto_in_r_bits_echo_extra_id,
  output auto_in_r_bits_echo_real_last,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_last) ; 
   wire _Queue_3_io_enq_ready ;  
   wire _Queue_3_io_deq_valid ;  
   wire [6:0] _Queue_3_io_deq_bits_extra_id ;  
   wire _Queue_3_io_deq_bits_real_last ;  
   wire _Queue_2_io_enq_ready ;  
   wire _Queue_2_io_deq_valid ;  
   wire [6:0] _Queue_2_io_deq_bits_extra_id ;  
   wire _Queue_2_io_deq_bits_real_last ;  
   wire _Queue_1_io_enq_ready ;  
   wire _Queue_1_io_deq_valid ;  
   wire [6:0] _Queue_1_io_deq_bits_extra_id ;  
   wire _Queue_1_io_deq_bits_real_last ;  
   wire _Queue_io_enq_ready ;  
   wire _Queue_io_deq_valid ;  
   wire [6:0] _Queue_io_deq_bits_extra_id ;  
   wire _Queue_io_deq_bits_real_last ;  
   wire _GEN=auto_in_ar_bits_id ? _Queue_1_io_enq_ready:_Queue_io_enq_ready ;  
   wire _GEN_0=auto_out_r_valid&auto_in_r_ready ;  
   wire _GEN_1=auto_in_ar_valid&auto_out_ar_ready ;  
   wire _GEN_2=auto_in_aw_bits_id ? _Queue_3_io_enq_ready:_Queue_2_io_enq_ready ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~auto_out_r_valid|(auto_out_r_bits_id ? _Queue_1_io_deq_valid:_Queue_io_deq_valid)))
            begin 
              if (1)$display("Assertion failed\n    at UserYanker.scala:66 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
              if (1)$display("");
            end 
         if (~reset&~(~auto_out_b_valid|(auto_out_b_bits_id ? _Queue_3_io_deq_valid:_Queue_2_io_deq_valid)))
            begin 
              if (1)$display("Assertion failed\n    at UserYanker.scala:95 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
              if (1)$display("");
            end 
       end
  
   wire _GEN_3=auto_out_b_valid&auto_in_b_ready ;  
   wire _GEN_4=auto_in_aw_valid&auto_out_aw_ready ;  
  Queue_28 Queue(.clock(clock),.reset(reset),.io_enq_ready(_Queue_io_enq_ready),.io_enq_valid(_GEN_1&~auto_in_ar_bits_id),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),.io_deq_ready(_GEN_0&~auto_out_r_bits_id&auto_out_r_bits_last),.io_deq_valid(_Queue_io_deq_valid),.io_deq_bits_extra_id(_Queue_io_deq_bits_extra_id),.io_deq_bits_real_last(_Queue_io_deq_bits_real_last)); 
  Queue_28 Queue_1(.clock(clock),.reset(reset),.io_enq_ready(_Queue_1_io_enq_ready),.io_enq_valid(_GEN_1&auto_in_ar_bits_id),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),.io_deq_ready(_GEN_0&auto_out_r_bits_id&auto_out_r_bits_last),.io_deq_valid(_Queue_1_io_deq_valid),.io_deq_bits_extra_id(_Queue_1_io_deq_bits_extra_id),.io_deq_bits_real_last(_Queue_1_io_deq_bits_real_last)); 
  Queue_28 Queue_2(.clock(clock),.reset(reset),.io_enq_ready(_Queue_2_io_enq_ready),.io_enq_valid(_GEN_4&~auto_in_aw_bits_id),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),.io_deq_ready(_GEN_3&~auto_out_b_bits_id),.io_deq_valid(_Queue_2_io_deq_valid),.io_deq_bits_extra_id(_Queue_2_io_deq_bits_extra_id),.io_deq_bits_real_last(_Queue_2_io_deq_bits_real_last)); 
  Queue_28 Queue_3(.clock(clock),.reset(reset),.io_enq_ready(_Queue_3_io_enq_ready),.io_enq_valid(_GEN_4&auto_in_aw_bits_id),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),.io_deq_ready(_GEN_3&auto_out_b_bits_id),.io_deq_valid(_Queue_3_io_deq_valid),.io_deq_bits_extra_id(_Queue_3_io_deq_bits_extra_id),.io_deq_bits_real_last(_Queue_3_io_deq_bits_real_last)); 
  assign auto_in_aw_ready=auto_out_aw_ready&_GEN_2; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_b_bits_echo_extra_id=auto_out_b_bits_id ? _Queue_3_io_deq_bits_extra_id:_Queue_2_io_deq_bits_extra_id; 
  assign auto_in_b_bits_echo_real_last=auto_out_b_bits_id ? _Queue_3_io_deq_bits_real_last:_Queue_2_io_deq_bits_real_last; 
  assign auto_in_ar_ready=auto_out_ar_ready&_GEN; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_echo_extra_id=auto_out_r_bits_id ? _Queue_1_io_deq_bits_extra_id:_Queue_io_deq_bits_extra_id; 
  assign auto_in_r_bits_echo_real_last=auto_out_r_bits_id ? _Queue_1_io_deq_bits_real_last:_Queue_io_deq_bits_real_last; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid&_GEN_2; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid&_GEN; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module Queue_32 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input io_enq_bits_id,
  input [31:0] io_enq_bits_addr,
  input [7:0] io_enq_bits_len,
  input [2:0] io_enq_bits_size,
  input [1:0] io_enq_bits_burst,
  input [6:0] io_enq_bits_echo_extra_id,
  input io_deq_ready,
  output io_deq_valid,
  output io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst,
  output [6:0] io_deq_bits_echo_extra_id) ; 
   reg [1:0] ram_burst ;  
   reg [2:0] ram_size ;  
   reg [7:0] ram_len ;  
   reg [31:0] ram_addr ;  
   reg ram_id ;  
   reg [6:0] ram_echo_extra_id ;  
   reg full ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire do_enq=~(~full&io_deq_ready)&~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_burst <=io_enq_bits_burst;
              ram_size <=io_enq_bits_size;
              ram_len <=io_enq_bits_len;
              ram_addr <=io_enq_bits_addr;
              ram_id <=io_enq_bits_id;
              ram_echo_extra_id <=io_enq_bits_echo_extra_id;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(full&io_deq_ready&io_deq_valid_0)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_id=full ? ram_id:io_enq_bits_id; 
  assign io_deq_bits_addr=full ? ram_addr:io_enq_bits_addr; 
  assign io_deq_bits_len=full ? ram_len:io_enq_bits_len; 
  assign io_deq_bits_size=full ? ram_size:io_enq_bits_size; 
  assign io_deq_bits_burst=full ? ram_burst:io_enq_bits_burst; 
  assign io_deq_bits_echo_extra_id=full ? ram_echo_extra_id:io_enq_bits_echo_extra_id; 
endmodule
 
module Queue_34 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [63:0] io_enq_bits_data,
  input [7:0] io_enq_bits_strb,
  input io_enq_bits_last,
  input io_deq_ready,
  output io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0] io_deq_bits_strb,
  output io_deq_bits_last) ; 
   reg ram_last ;  
   reg [7:0] ram_strb ;  
   reg [63:0] ram_data ;  
   reg full ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire do_enq=~(~full&io_deq_ready)&~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_last <=io_enq_bits_last;
              ram_strb <=io_enq_bits_strb;
              ram_data <=io_enq_bits_data;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(full&io_deq_ready&io_deq_valid_0)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_data=full ? ram_data:io_enq_bits_data; 
  assign io_deq_bits_strb=full ? ram_strb:io_enq_bits_strb; 
  assign io_deq_bits_last=full ? ram_last:io_enq_bits_last; 
endmodule
 
module AXI4Fragmenter (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [1:0] auto_in_aw_bits_burst,
  input [6:0] auto_in_aw_bits_echo_extra_id,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output [6:0] auto_in_b_bits_echo_extra_id,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [1:0] auto_in_ar_bits_burst,
  input [6:0] auto_in_ar_bits_echo_extra_id,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output [6:0] auto_in_r_bits_echo_extra_id,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [6:0] auto_out_aw_bits_echo_extra_id,
  output auto_out_aw_bits_echo_real_last,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input [6:0] auto_out_b_bits_echo_extra_id,
  input auto_out_b_bits_echo_real_last,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [6:0] auto_out_ar_bits_echo_extra_id,
  output auto_out_ar_bits_echo_real_last,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input [6:0] auto_out_r_bits_echo_extra_id,
  input auto_out_r_bits_echo_real_last,
  input auto_out_r_bits_last) ; 
   wire nodeOut_w_valid ;  
   wire w_idle ;  
   wire in_aw_ready ;  
   wire _in_w_deq_q_io_deq_valid ;  
   wire _in_w_deq_q_io_deq_bits_last ;  
   wire _deq_q_1_io_deq_valid ;  
   wire [31:0] _deq_q_1_io_deq_bits_addr ;  
   wire [7:0] _deq_q_1_io_deq_bits_len ;  
   wire [2:0] _deq_q_1_io_deq_bits_size ;  
   wire [1:0] _deq_q_1_io_deq_bits_burst ;  
   wire _deq_q_io_deq_valid ;  
   wire [31:0] _deq_q_io_deq_bits_addr ;  
   wire [7:0] _deq_q_io_deq_bits_len ;  
   wire [2:0] _deq_q_io_deq_bits_size ;  
   wire [1:0] _deq_q_io_deq_bits_burst ;  
   reg busy ;  
   reg [31:0] r_addr ;  
   reg [7:0] r_len ;  
   wire [7:0] len=busy ? r_len:_deq_q_io_deq_bits_len ;  
   wire [31:0] addr=busy ? r_addr:_deq_q_io_deq_bits_addr ;  
   wire [5:0] _GEN=len[6:1]|len[7:2] ;  
   wire [4:0] _GEN_0=_GEN[4:0]|{len[7],_GEN[5:2]} ;  
   wire [7:0] _wipeHigh_T=~len ;  
   wire [7:0] _wipeHigh_T_3=_wipeHigh_T|{_wipeHigh_T[6:0],1'h0} ;  
   wire [7:0] _wipeHigh_T_6=_wipeHigh_T_3|{_wipeHigh_T_3[5:0],2'h0} ;  
   wire [7:0] _align1_T_2=addr[10:3]|{addr[9:3],1'h0} ;  
   wire [7:0] _align1_T_5=_align1_T_2|{_align1_T_2[5:0],2'h0} ;  
   wire fixed=_deq_q_io_deq_bits_burst==2'h0 ;  
   wire [7:0] beats1=fixed|_deq_q_io_deq_bits_size!=3'h3 ? 8'h0:({1'h0,len[7],_GEN[5],_GEN_0[4:3],_GEN_0[2:0]|{len[7],_GEN[5],_GEN_0[4]}}|~(_wipeHigh_T_6|{_wipeHigh_T_6[3:0],4'h0}))&~(_align1_T_5|{_align1_T_5[3:0],4'h0})&({5'h0,{3{{addr[31:30],addr[27],addr[25],addr[16],addr[13]}==6'h0|{addr[31:30],addr[27],addr[25],~(addr[16])}==5'h0|{addr[31:30],addr[27],~(addr[25]),addr[16]}==5'h0|{addr[31:30],~(addr[27])}==3'h0|{addr[31],~(addr[30])}==2'h0|addr[31:30]==2'h2}}}|{8{{addr[31:30],addr[27],addr[25],addr[16],~(addr[13])}==6'h0}}) ;  
   wire ar_last=beats1==len ;  
   wire [31:0] _out_bits_addr_T=~addr ;  
   wire [9:0] _out_bits_addr_T_2=10'h7<<_deq_q_io_deq_bits_size ;  
   reg busy_1 ;  
   reg [31:0] r_addr_1 ;  
   reg [7:0] r_len_1 ;  
   wire [7:0] len_1=busy_1 ? r_len_1:_deq_q_1_io_deq_bits_len ;  
   wire [31:0] addr_1=busy_1 ? r_addr_1:_deq_q_1_io_deq_bits_addr ;  
   wire [7:0] _support1_T_79={5'h0,{3{{addr_1[31:30],addr_1[27],addr_1[25],addr_1[13]}==5'h0|{addr_1[31:30],addr_1[27],~(addr_1[25])}==4'h0|{addr_1[31:30],~(addr_1[27])}==3'h0|addr_1[31:30]==2'h2}}}|{8{{addr_1[31:30],addr_1[27],addr_1[25],~(addr_1[13])}==5'h0}} ;  
   wire [5:0] _GEN_1=len_1[6:1]|len_1[7:2] ;  
   wire [4:0] _GEN_2=_GEN_1[4:0]|{len_1[7],_GEN_1[5:2]} ;  
   wire [7:0] _wipeHigh_T_11=~len_1 ;  
   wire [7:0] _wipeHigh_T_14=_wipeHigh_T_11|{_wipeHigh_T_11[6:0],1'h0} ;  
   wire [7:0] _wipeHigh_T_17=_wipeHigh_T_14|{_wipeHigh_T_14[5:0],2'h0} ;  
   wire [7:0] _align1_T_12=addr_1[10:3]|{addr_1[9:3],1'h0} ;  
   wire [7:0] _align1_T_15=_align1_T_12|{_align1_T_12[5:0],2'h0} ;  
   wire fixed_1=_deq_q_1_io_deq_bits_burst==2'h0 ;  
   wire [7:0] beats1_1=fixed_1|_deq_q_1_io_deq_bits_size!=3'h3 ? 8'h0:({1'h0,len_1[7],_GEN_1[5],_GEN_2[4:3],_GEN_2[2:0]|{len_1[7],_GEN_1[5],_GEN_2[4]}}|~(_wipeHigh_T_17|{_wipeHigh_T_17[3:0],4'h0}))&~(_align1_T_15|{_align1_T_15[3:0],4'h0})&{_support1_T_79[7:5],_support1_T_79[4:0]|{5{{addr_1[31],~(addr_1[30])}==2'h0}}} ;  
   wire [8:0] w_beats={beats1_1,1'h1}&{1'h1,~beats1_1} ;  
   wire aw_last=beats1_1==len_1 ;  
   wire [31:0] _out_bits_addr_T_7=~addr_1 ;  
   wire [9:0] _out_bits_addr_T_9=10'h7<<_deq_q_1_io_deq_bits_size ;  
   reg wbeats_latched ;  
   wire _in_aw_ready_T=w_idle|wbeats_latched ;  
   wire nodeOut_aw_valid=_deq_q_1_io_deq_valid&_in_aw_ready_T ;  
  assign in_aw_ready=auto_out_aw_ready&_in_aw_ready_T; 
   wire wbeats_valid=_deq_q_1_io_deq_valid&~wbeats_latched ;  
   reg [8:0] w_counter ;  
  assign w_idle=w_counter==9'h0; 
   wire [8:0] w_todo=w_idle ? (wbeats_valid ? w_beats:9'h0):w_counter ;  
   wire w_last=w_todo==9'h1 ;  
   wire _w_counter_T=auto_out_w_ready&nodeOut_w_valid ;  
  assign nodeOut_w_valid=_in_w_deq_q_io_deq_valid&(~w_idle|wbeats_valid); 
  always @( posedge clock)
       begin 
         if (~reset&~(~_w_counter_T|(|w_todo)))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:177 assert (!out.w.fire || w_todo =/= 0.U) // underflow impossible\n");
              if (1)$display("");
            end 
         if (~reset&~(~nodeOut_w_valid|~_in_w_deq_q_io_deq_bits_last|w_last))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:186 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
              if (1)$display("");
            end 
       end
  
   wire nodeOut_b_ready=auto_in_b_ready|~auto_out_b_bits_echo_real_last ;  
   reg [1:0] error_0 ;  
   reg [1:0] error_1 ;  
   wire _GEN_3=nodeOut_b_ready&auto_out_b_valid ;  
   wire [22:0] _wrapMask_T_1={7'h0,_deq_q_io_deq_bits_len,8'hFF}<<_deq_q_io_deq_bits_size ;  
   wire [31:0] _mux_addr_T_1=~_deq_q_io_deq_bits_addr ;  
   wire [8:0] beats={beats1,1'h1}&{1'h1,~beats1} ;  
   wire [31:0] _inc_addr_T_1=addr+{16'h0,{7'h0,beats}<<_deq_q_io_deq_bits_size} ;  
   wire [22:0] _wrapMask_T_3={7'h0,_deq_q_1_io_deq_bits_len,8'hFF}<<_deq_q_1_io_deq_bits_size ;  
   wire [31:0] _mux_addr_T_6=~_deq_q_1_io_deq_bits_addr ;  
   wire [31:0] _inc_addr_T_3=addr_1+{16'h0,{7'h0,w_beats}<<_deq_q_1_io_deq_bits_size} ;  
   wire _GEN_4=auto_out_ar_ready&_deq_q_io_deq_valid ;  
   wire _GEN_5=in_aw_ready&_deq_q_1_io_deq_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              busy <=1'h0;
              busy_1 <=1'h0;
              wbeats_latched <=1'h0;
              w_counter <=9'h0;
              error_0 <=2'h0;
              error_1 <=2'h0;
            end 
          else 
            begin 
              if (_GEN_4)
                 busy <=~ar_last;
              if (_GEN_5)
                 busy_1 <=~aw_last;
              wbeats_latched <=~(auto_out_aw_ready&nodeOut_aw_valid)&(wbeats_valid&w_idle|wbeats_latched);
              w_counter <=w_todo-{8'h0,_w_counter_T};
              if (~auto_out_b_bits_id&_GEN_3)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_0 <=2'h0;
                    else 
                      error_0 <=error_0|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id&_GEN_3)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_1 <=2'h0;
                    else 
                      error_1 <=error_1|auto_out_b_bits_resp;
                 end 
            end 
         if (_GEN_4)
            begin 
              if (fixed)
                 r_addr <=_deq_q_io_deq_bits_addr;
               else 
                 if (_deq_q_io_deq_bits_burst==2'h2)
                    r_addr <={17'h0,_inc_addr_T_1[14:0]&_wrapMask_T_1[22:8]}|~{_mux_addr_T_1[31:15],_mux_addr_T_1[14:0]|_wrapMask_T_1[22:8]};
                  else 
                    r_addr <=_inc_addr_T_1;
              r_len <=len-beats[7:0];
            end 
         if (_GEN_5)
            begin 
              if (fixed_1)
                 r_addr_1 <=_deq_q_1_io_deq_bits_addr;
               else 
                 if (_deq_q_1_io_deq_bits_burst==2'h2)
                    r_addr_1 <={17'h0,_inc_addr_T_3[14:0]&_wrapMask_T_3[22:8]}|~{_mux_addr_T_6[31:15],_mux_addr_T_6[14:0]|_wrapMask_T_3[22:8]};
                  else 
                    r_addr_1 <=_inc_addr_T_3;
              r_len_1 <=len_1-w_beats[7:0];
            end 
       end
  
  Queue_32 deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_ar_ready),.io_enq_valid(auto_in_ar_valid),.io_enq_bits_id(auto_in_ar_bits_id),.io_enq_bits_addr(auto_in_ar_bits_addr),.io_enq_bits_len(auto_in_ar_bits_len),.io_enq_bits_size(auto_in_ar_bits_size),.io_enq_bits_burst(auto_in_ar_bits_burst),.io_enq_bits_echo_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(auto_out_ar_ready&ar_last),.io_deq_valid(_deq_q_io_deq_valid),.io_deq_bits_id(auto_out_ar_bits_id),.io_deq_bits_addr(_deq_q_io_deq_bits_addr),.io_deq_bits_len(_deq_q_io_deq_bits_len),.io_deq_bits_size(_deq_q_io_deq_bits_size),.io_deq_bits_burst(_deq_q_io_deq_bits_burst),.io_deq_bits_echo_extra_id(auto_out_ar_bits_echo_extra_id)); 
  Queue_32 deq_q_1(.clock(clock),.reset(reset),.io_enq_ready(auto_in_aw_ready),.io_enq_valid(auto_in_aw_valid),.io_enq_bits_id(auto_in_aw_bits_id),.io_enq_bits_addr(auto_in_aw_bits_addr),.io_enq_bits_len(auto_in_aw_bits_len),.io_enq_bits_size(auto_in_aw_bits_size),.io_enq_bits_burst(auto_in_aw_bits_burst),.io_enq_bits_echo_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(in_aw_ready&aw_last),.io_deq_valid(_deq_q_1_io_deq_valid),.io_deq_bits_id(auto_out_aw_bits_id),.io_deq_bits_addr(_deq_q_1_io_deq_bits_addr),.io_deq_bits_len(_deq_q_1_io_deq_bits_len),.io_deq_bits_size(_deq_q_1_io_deq_bits_size),.io_deq_bits_burst(_deq_q_1_io_deq_bits_burst),.io_deq_bits_echo_extra_id(auto_out_aw_bits_echo_extra_id)); 
  Queue_34 in_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_w_ready),.io_enq_valid(auto_in_w_valid),.io_enq_bits_data(auto_in_w_bits_data),.io_enq_bits_strb(auto_in_w_bits_strb),.io_enq_bits_last(auto_in_w_bits_last),.io_deq_ready(auto_out_w_ready&(~w_idle|wbeats_valid)),.io_deq_valid(_in_w_deq_q_io_deq_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last(_in_w_deq_q_io_deq_bits_last)); 
  assign auto_in_b_valid=auto_out_b_valid&auto_out_b_bits_echo_real_last; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp|(auto_out_b_bits_id ? error_1:error_0); 
  assign auto_in_b_bits_echo_extra_id=auto_out_b_bits_echo_extra_id; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_echo_extra_id=auto_out_r_bits_echo_extra_id; 
  assign auto_in_r_bits_last=auto_out_r_bits_last&auto_out_r_bits_echo_real_last; 
  assign auto_out_aw_valid=nodeOut_aw_valid; 
  assign auto_out_aw_bits_addr=~{_out_bits_addr_T_7[31:3],_out_bits_addr_T_7[2:0]|~(_out_bits_addr_T_9[2:0])}; 
  assign auto_out_aw_bits_len=beats1_1; 
  assign auto_out_aw_bits_size=_deq_q_1_io_deq_bits_size; 
  assign auto_out_aw_bits_echo_real_last=aw_last; 
  assign auto_out_w_valid=nodeOut_w_valid; 
  assign auto_out_w_bits_last=w_last; 
  assign auto_out_b_ready=nodeOut_b_ready; 
  assign auto_out_ar_valid=_deq_q_io_deq_valid; 
  assign auto_out_ar_bits_addr=~{_out_bits_addr_T[31:3],_out_bits_addr_T[2:0]|~(_out_bits_addr_T_2[2:0])}; 
  assign auto_out_ar_bits_len=beats1; 
  assign auto_out_ar_bits_size=_deq_q_io_deq_bits_size; 
  assign auto_out_ar_bits_echo_real_last=ar_last; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module AXI4IdIndexer_1 (
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [7:0] auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [1:0] auto_in_aw_bits_burst,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [7:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [7:0] auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [1:0] auto_in_ar_bits_burst,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [7:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [1:0] auto_out_aw_bits_burst,
  output [6:0] auto_out_aw_bits_echo_extra_id,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input [6:0] auto_out_b_bits_echo_extra_id,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [1:0] auto_out_ar_bits_burst,
  output [6:0] auto_out_ar_bits_echo_extra_id,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input [6:0] auto_out_r_bits_echo_extra_id,
  input auto_out_r_bits_last) ; 
  assign auto_in_aw_ready=auto_out_aw_ready; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id={auto_out_b_bits_echo_extra_id,auto_out_b_bits_id}; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_ar_ready=auto_out_ar_ready; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id={auto_out_r_bits_echo_extra_id,auto_out_r_bits_id}; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id[0]; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_aw_bits_burst=auto_in_aw_bits_burst; 
  assign auto_out_aw_bits_echo_extra_id=auto_in_aw_bits_id[7:1]; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id[0]; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_ar_bits_burst=auto_in_ar_bits_burst; 
  assign auto_out_ar_bits_echo_extra_id=auto_in_ar_bits_id[7:1]; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module TLInterconnectCoupler_5 (
  input clock,
  input reset,
  output auto_axi4index_in_aw_ready,
  input auto_axi4index_in_aw_valid,
  input [7:0] auto_axi4index_in_aw_bits_id,
  input [31:0] auto_axi4index_in_aw_bits_addr,
  input [7:0] auto_axi4index_in_aw_bits_len,
  input [2:0] auto_axi4index_in_aw_bits_size,
  input [1:0] auto_axi4index_in_aw_bits_burst,
  output auto_axi4index_in_w_ready,
  input auto_axi4index_in_w_valid,
  input [63:0] auto_axi4index_in_w_bits_data,
  input [7:0] auto_axi4index_in_w_bits_strb,
  input auto_axi4index_in_w_bits_last,
  input auto_axi4index_in_b_ready,
  output auto_axi4index_in_b_valid,
  output [7:0] auto_axi4index_in_b_bits_id,
  output [1:0] auto_axi4index_in_b_bits_resp,
  output auto_axi4index_in_ar_ready,
  input auto_axi4index_in_ar_valid,
  input [7:0] auto_axi4index_in_ar_bits_id,
  input [31:0] auto_axi4index_in_ar_bits_addr,
  input [7:0] auto_axi4index_in_ar_bits_len,
  input [2:0] auto_axi4index_in_ar_bits_size,
  input [1:0] auto_axi4index_in_ar_bits_burst,
  input auto_axi4index_in_r_ready,
  output auto_axi4index_in_r_valid,
  output [7:0] auto_axi4index_in_r_bits_id,
  output [63:0] auto_axi4index_in_r_bits_data,
  output [1:0] auto_axi4index_in_r_bits_resp,
  output auto_axi4index_in_r_bits_last,
  input auto_tl_out_a_ready,
  output auto_tl_out_a_valid,
  output [2:0] auto_tl_out_a_bits_opcode,
  output [2:0] auto_tl_out_a_bits_param,
  output [3:0] auto_tl_out_a_bits_size,
  output [3:0] auto_tl_out_a_bits_source,
  output [31:0] auto_tl_out_a_bits_address,
  output [7:0] auto_tl_out_a_bits_mask,
  output [63:0] auto_tl_out_a_bits_data,
  output auto_tl_out_a_bits_corrupt,
  output auto_tl_out_d_ready,
  input auto_tl_out_d_valid,
  input [2:0] auto_tl_out_d_bits_opcode,
  input [1:0] auto_tl_out_d_bits_param,
  input [3:0] auto_tl_out_d_bits_size,
  input [3:0] auto_tl_out_d_bits_source,
  input [1:0] auto_tl_out_d_bits_sink,
  input auto_tl_out_d_bits_denied,
  input [63:0] auto_tl_out_d_bits_data,
  input auto_tl_out_d_bits_corrupt) ; 
   wire _axi4index_auto_out_aw_valid ;  
   wire _axi4index_auto_out_aw_bits_id ;  
   wire [31:0] _axi4index_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4index_auto_out_aw_bits_len ;  
   wire [2:0] _axi4index_auto_out_aw_bits_size ;  
   wire [1:0] _axi4index_auto_out_aw_bits_burst ;  
   wire [6:0] _axi4index_auto_out_aw_bits_echo_extra_id ;  
   wire _axi4index_auto_out_w_valid ;  
   wire [63:0] _axi4index_auto_out_w_bits_data ;  
   wire [7:0] _axi4index_auto_out_w_bits_strb ;  
   wire _axi4index_auto_out_w_bits_last ;  
   wire _axi4index_auto_out_b_ready ;  
   wire _axi4index_auto_out_ar_valid ;  
   wire _axi4index_auto_out_ar_bits_id ;  
   wire [31:0] _axi4index_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4index_auto_out_ar_bits_len ;  
   wire [2:0] _axi4index_auto_out_ar_bits_size ;  
   wire [1:0] _axi4index_auto_out_ar_bits_burst ;  
   wire [6:0] _axi4index_auto_out_ar_bits_echo_extra_id ;  
   wire _axi4index_auto_out_r_ready ;  
   wire _axi4frag_auto_in_aw_ready ;  
   wire _axi4frag_auto_in_w_ready ;  
   wire _axi4frag_auto_in_b_valid ;  
   wire _axi4frag_auto_in_b_bits_id ;  
   wire [1:0] _axi4frag_auto_in_b_bits_resp ;  
   wire [6:0] _axi4frag_auto_in_b_bits_echo_extra_id ;  
   wire _axi4frag_auto_in_ar_ready ;  
   wire _axi4frag_auto_in_r_valid ;  
   wire _axi4frag_auto_in_r_bits_id ;  
   wire [63:0] _axi4frag_auto_in_r_bits_data ;  
   wire [1:0] _axi4frag_auto_in_r_bits_resp ;  
   wire [6:0] _axi4frag_auto_in_r_bits_echo_extra_id ;  
   wire _axi4frag_auto_in_r_bits_last ;  
   wire _axi4frag_auto_out_aw_valid ;  
   wire _axi4frag_auto_out_aw_bits_id ;  
   wire [31:0] _axi4frag_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4frag_auto_out_aw_bits_len ;  
   wire [2:0] _axi4frag_auto_out_aw_bits_size ;  
   wire [6:0] _axi4frag_auto_out_aw_bits_echo_extra_id ;  
   wire _axi4frag_auto_out_aw_bits_echo_real_last ;  
   wire _axi4frag_auto_out_w_valid ;  
   wire [63:0] _axi4frag_auto_out_w_bits_data ;  
   wire [7:0] _axi4frag_auto_out_w_bits_strb ;  
   wire _axi4frag_auto_out_w_bits_last ;  
   wire _axi4frag_auto_out_b_ready ;  
   wire _axi4frag_auto_out_ar_valid ;  
   wire _axi4frag_auto_out_ar_bits_id ;  
   wire [31:0] _axi4frag_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4frag_auto_out_ar_bits_len ;  
   wire [2:0] _axi4frag_auto_out_ar_bits_size ;  
   wire [6:0] _axi4frag_auto_out_ar_bits_echo_extra_id ;  
   wire _axi4frag_auto_out_ar_bits_echo_real_last ;  
   wire _axi4frag_auto_out_r_ready ;  
   wire _axi4yank_auto_in_aw_ready ;  
   wire _axi4yank_auto_in_w_ready ;  
   wire _axi4yank_auto_in_b_valid ;  
   wire _axi4yank_auto_in_b_bits_id ;  
   wire [1:0] _axi4yank_auto_in_b_bits_resp ;  
   wire [6:0] _axi4yank_auto_in_b_bits_echo_extra_id ;  
   wire _axi4yank_auto_in_b_bits_echo_real_last ;  
   wire _axi4yank_auto_in_ar_ready ;  
   wire _axi4yank_auto_in_r_valid ;  
   wire _axi4yank_auto_in_r_bits_id ;  
   wire [63:0] _axi4yank_auto_in_r_bits_data ;  
   wire [1:0] _axi4yank_auto_in_r_bits_resp ;  
   wire [6:0] _axi4yank_auto_in_r_bits_echo_extra_id ;  
   wire _axi4yank_auto_in_r_bits_echo_real_last ;  
   wire _axi4yank_auto_in_r_bits_last ;  
   wire _axi4yank_auto_out_aw_valid ;  
   wire _axi4yank_auto_out_aw_bits_id ;  
   wire [31:0] _axi4yank_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4yank_auto_out_aw_bits_len ;  
   wire [2:0] _axi4yank_auto_out_aw_bits_size ;  
   wire _axi4yank_auto_out_w_valid ;  
   wire [63:0] _axi4yank_auto_out_w_bits_data ;  
   wire [7:0] _axi4yank_auto_out_w_bits_strb ;  
   wire _axi4yank_auto_out_w_bits_last ;  
   wire _axi4yank_auto_out_b_ready ;  
   wire _axi4yank_auto_out_ar_valid ;  
   wire _axi4yank_auto_out_ar_bits_id ;  
   wire [31:0] _axi4yank_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4yank_auto_out_ar_bits_len ;  
   wire [2:0] _axi4yank_auto_out_ar_bits_size ;  
   wire _axi4yank_auto_out_r_ready ;  
   wire _axi42tl_auto_in_aw_ready ;  
   wire _axi42tl_auto_in_w_ready ;  
   wire _axi42tl_auto_in_b_valid ;  
   wire _axi42tl_auto_in_b_bits_id ;  
   wire [1:0] _axi42tl_auto_in_b_bits_resp ;  
   wire _axi42tl_auto_in_ar_ready ;  
   wire _axi42tl_auto_in_r_valid ;  
   wire _axi42tl_auto_in_r_bits_id ;  
   wire [63:0] _axi42tl_auto_in_r_bits_data ;  
   wire [1:0] _axi42tl_auto_in_r_bits_resp ;  
   wire _axi42tl_auto_in_r_bits_last ;  
   wire _axi42tl_auto_out_a_valid ;  
   wire [2:0] _axi42tl_auto_out_a_bits_opcode ;  
   wire [3:0] _axi42tl_auto_out_a_bits_size ;  
   wire [3:0] _axi42tl_auto_out_a_bits_source ;  
   wire [31:0] _axi42tl_auto_out_a_bits_address ;  
   wire [7:0] _axi42tl_auto_out_a_bits_mask ;  
   wire [63:0] _axi42tl_auto_out_a_bits_data ;  
   wire _axi42tl_auto_out_d_ready ;  
   wire _fixer_auto_in_a_ready ;  
   wire _fixer_auto_in_d_valid ;  
   wire [2:0] _fixer_auto_in_d_bits_opcode ;  
   wire [3:0] _fixer_auto_in_d_bits_size ;  
   wire [3:0] _fixer_auto_in_d_bits_source ;  
   wire _fixer_auto_in_d_bits_denied ;  
   wire [63:0] _fixer_auto_in_d_bits_data ;  
   wire _fixer_auto_in_d_bits_corrupt ;  
   wire _fixer_auto_out_a_valid ;  
   wire [2:0] _fixer_auto_out_a_bits_opcode ;  
   wire [3:0] _fixer_auto_out_a_bits_size ;  
   wire [3:0] _fixer_auto_out_a_bits_source ;  
   wire [31:0] _fixer_auto_out_a_bits_address ;  
   wire [7:0] _fixer_auto_out_a_bits_mask ;  
   wire [63:0] _fixer_auto_out_a_bits_data ;  
   wire _fixer_auto_out_d_ready ;  
   wire _buffer_auto_in_a_ready ;  
   wire _buffer_auto_in_d_valid ;  
   wire [2:0] _buffer_auto_in_d_bits_opcode ;  
   wire [1:0] _buffer_auto_in_d_bits_param ;  
   wire [3:0] _buffer_auto_in_d_bits_size ;  
   wire [3:0] _buffer_auto_in_d_bits_source ;  
   wire [1:0] _buffer_auto_in_d_bits_sink ;  
   wire _buffer_auto_in_d_bits_denied ;  
   wire [63:0] _buffer_auto_in_d_bits_data ;  
   wire _buffer_auto_in_d_bits_corrupt ;  
  TLBuffer_3 buffer(.clock(clock),.reset(reset),.auto_in_a_ready(_buffer_auto_in_a_ready),.auto_in_a_valid(_fixer_auto_out_a_valid),.auto_in_a_bits_opcode(_fixer_auto_out_a_bits_opcode),.auto_in_a_bits_size(_fixer_auto_out_a_bits_size),.auto_in_a_bits_source(_fixer_auto_out_a_bits_source),.auto_in_a_bits_address(_fixer_auto_out_a_bits_address),.auto_in_a_bits_mask(_fixer_auto_out_a_bits_mask),.auto_in_a_bits_data(_fixer_auto_out_a_bits_data),.auto_in_d_ready(_fixer_auto_out_d_ready),.auto_in_d_valid(_buffer_auto_in_d_valid),.auto_in_d_bits_opcode(_buffer_auto_in_d_bits_opcode),.auto_in_d_bits_param(_buffer_auto_in_d_bits_param),.auto_in_d_bits_size(_buffer_auto_in_d_bits_size),.auto_in_d_bits_source(_buffer_auto_in_d_bits_source),.auto_in_d_bits_sink(_buffer_auto_in_d_bits_sink),.auto_in_d_bits_denied(_buffer_auto_in_d_bits_denied),.auto_in_d_bits_data(_buffer_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt),.auto_out_a_ready(auto_tl_out_a_ready),.auto_out_a_valid(auto_tl_out_a_valid),.auto_out_a_bits_opcode(auto_tl_out_a_bits_opcode),.auto_out_a_bits_param(auto_tl_out_a_bits_param),.auto_out_a_bits_size(auto_tl_out_a_bits_size),.auto_out_a_bits_source(auto_tl_out_a_bits_source),.auto_out_a_bits_address(auto_tl_out_a_bits_address),.auto_out_a_bits_mask(auto_tl_out_a_bits_mask),.auto_out_a_bits_data(auto_tl_out_a_bits_data),.auto_out_a_bits_corrupt(auto_tl_out_a_bits_corrupt),.auto_out_d_ready(auto_tl_out_d_ready),.auto_out_d_valid(auto_tl_out_d_valid),.auto_out_d_bits_opcode(auto_tl_out_d_bits_opcode),.auto_out_d_bits_param(auto_tl_out_d_bits_param),.auto_out_d_bits_size(auto_tl_out_d_bits_size),.auto_out_d_bits_source(auto_tl_out_d_bits_source),.auto_out_d_bits_sink(auto_tl_out_d_bits_sink),.auto_out_d_bits_denied(auto_tl_out_d_bits_denied),.auto_out_d_bits_data(auto_tl_out_d_bits_data),.auto_out_d_bits_corrupt(auto_tl_out_d_bits_corrupt)); 
  TLFIFOFixer_2 fixer(.clock(clock),.reset(reset),.auto_in_a_ready(_fixer_auto_in_a_ready),.auto_in_a_valid(_axi42tl_auto_out_a_valid),.auto_in_a_bits_opcode(_axi42tl_auto_out_a_bits_opcode),.auto_in_a_bits_size(_axi42tl_auto_out_a_bits_size),.auto_in_a_bits_source(_axi42tl_auto_out_a_bits_source),.auto_in_a_bits_address(_axi42tl_auto_out_a_bits_address),.auto_in_a_bits_mask(_axi42tl_auto_out_a_bits_mask),.auto_in_a_bits_data(_axi42tl_auto_out_a_bits_data),.auto_in_d_ready(_axi42tl_auto_out_d_ready),.auto_in_d_valid(_fixer_auto_in_d_valid),.auto_in_d_bits_opcode(_fixer_auto_in_d_bits_opcode),.auto_in_d_bits_size(_fixer_auto_in_d_bits_size),.auto_in_d_bits_source(_fixer_auto_in_d_bits_source),.auto_in_d_bits_denied(_fixer_auto_in_d_bits_denied),.auto_in_d_bits_data(_fixer_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_fixer_auto_in_d_bits_corrupt),.auto_out_a_ready(_buffer_auto_in_a_ready),.auto_out_a_valid(_fixer_auto_out_a_valid),.auto_out_a_bits_opcode(_fixer_auto_out_a_bits_opcode),.auto_out_a_bits_size(_fixer_auto_out_a_bits_size),.auto_out_a_bits_source(_fixer_auto_out_a_bits_source),.auto_out_a_bits_address(_fixer_auto_out_a_bits_address),.auto_out_a_bits_mask(_fixer_auto_out_a_bits_mask),.auto_out_a_bits_data(_fixer_auto_out_a_bits_data),.auto_out_d_ready(_fixer_auto_out_d_ready),.auto_out_d_valid(_buffer_auto_in_d_valid),.auto_out_d_bits_opcode(_buffer_auto_in_d_bits_opcode),.auto_out_d_bits_param(_buffer_auto_in_d_bits_param),.auto_out_d_bits_size(_buffer_auto_in_d_bits_size),.auto_out_d_bits_source(_buffer_auto_in_d_bits_source),.auto_out_d_bits_sink(_buffer_auto_in_d_bits_sink),.auto_out_d_bits_denied(_buffer_auto_in_d_bits_denied),.auto_out_d_bits_data(_buffer_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt)); 
  AXI4ToTL axi42tl(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi42tl_auto_in_aw_ready),.auto_in_aw_valid(_axi4yank_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4yank_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4yank_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4yank_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4yank_auto_out_aw_bits_size),.auto_in_w_ready(_axi42tl_auto_in_w_ready),.auto_in_w_valid(_axi4yank_auto_out_w_valid),.auto_in_w_bits_data(_axi4yank_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4yank_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4yank_auto_out_w_bits_last),.auto_in_b_ready(_axi4yank_auto_out_b_ready),.auto_in_b_valid(_axi42tl_auto_in_b_valid),.auto_in_b_bits_id(_axi42tl_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi42tl_auto_in_b_bits_resp),.auto_in_ar_ready(_axi42tl_auto_in_ar_ready),.auto_in_ar_valid(_axi4yank_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4yank_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4yank_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4yank_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4yank_auto_out_ar_bits_size),.auto_in_r_ready(_axi4yank_auto_out_r_ready),.auto_in_r_valid(_axi42tl_auto_in_r_valid),.auto_in_r_bits_id(_axi42tl_auto_in_r_bits_id),.auto_in_r_bits_data(_axi42tl_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi42tl_auto_in_r_bits_resp),.auto_in_r_bits_last(_axi42tl_auto_in_r_bits_last),.auto_out_a_ready(_fixer_auto_in_a_ready),.auto_out_a_valid(_axi42tl_auto_out_a_valid),.auto_out_a_bits_opcode(_axi42tl_auto_out_a_bits_opcode),.auto_out_a_bits_size(_axi42tl_auto_out_a_bits_size),.auto_out_a_bits_source(_axi42tl_auto_out_a_bits_source),.auto_out_a_bits_address(_axi42tl_auto_out_a_bits_address),.auto_out_a_bits_mask(_axi42tl_auto_out_a_bits_mask),.auto_out_a_bits_data(_axi42tl_auto_out_a_bits_data),.auto_out_d_ready(_axi42tl_auto_out_d_ready),.auto_out_d_valid(_fixer_auto_in_d_valid),.auto_out_d_bits_opcode(_fixer_auto_in_d_bits_opcode),.auto_out_d_bits_size(_fixer_auto_in_d_bits_size),.auto_out_d_bits_source(_fixer_auto_in_d_bits_source),.auto_out_d_bits_denied(_fixer_auto_in_d_bits_denied),.auto_out_d_bits_data(_fixer_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_fixer_auto_in_d_bits_corrupt)); 
  AXI4UserYanker_1 axi4yank(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4yank_auto_in_aw_ready),.auto_in_aw_valid(_axi4frag_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4frag_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4frag_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4frag_auto_out_aw_bits_size),.auto_in_aw_bits_echo_extra_id(_axi4frag_auto_out_aw_bits_echo_extra_id),.auto_in_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),.auto_in_w_ready(_axi4yank_auto_in_w_ready),.auto_in_w_valid(_axi4frag_auto_out_w_valid),.auto_in_w_bits_data(_axi4frag_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4frag_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4frag_auto_out_w_bits_last),.auto_in_b_ready(_axi4frag_auto_out_b_ready),.auto_in_b_valid(_axi4yank_auto_in_b_valid),.auto_in_b_bits_id(_axi4yank_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4yank_auto_in_b_bits_resp),.auto_in_b_bits_echo_extra_id(_axi4yank_auto_in_b_bits_echo_extra_id),.auto_in_b_bits_echo_real_last(_axi4yank_auto_in_b_bits_echo_real_last),.auto_in_ar_ready(_axi4yank_auto_in_ar_ready),.auto_in_ar_valid(_axi4frag_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4frag_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4frag_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4frag_auto_out_ar_bits_size),.auto_in_ar_bits_echo_extra_id(_axi4frag_auto_out_ar_bits_echo_extra_id),.auto_in_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),.auto_in_r_ready(_axi4frag_auto_out_r_ready),.auto_in_r_valid(_axi4yank_auto_in_r_valid),.auto_in_r_bits_id(_axi4yank_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4yank_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4yank_auto_in_r_bits_resp),.auto_in_r_bits_echo_extra_id(_axi4yank_auto_in_r_bits_echo_extra_id),.auto_in_r_bits_echo_real_last(_axi4yank_auto_in_r_bits_echo_real_last),.auto_in_r_bits_last(_axi4yank_auto_in_r_bits_last),.auto_out_aw_ready(_axi42tl_auto_in_aw_ready),.auto_out_aw_valid(_axi4yank_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4yank_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4yank_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4yank_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4yank_auto_out_aw_bits_size),.auto_out_w_ready(_axi42tl_auto_in_w_ready),.auto_out_w_valid(_axi4yank_auto_out_w_valid),.auto_out_w_bits_data(_axi4yank_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4yank_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4yank_auto_out_w_bits_last),.auto_out_b_ready(_axi4yank_auto_out_b_ready),.auto_out_b_valid(_axi42tl_auto_in_b_valid),.auto_out_b_bits_id(_axi42tl_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi42tl_auto_in_b_bits_resp),.auto_out_ar_ready(_axi42tl_auto_in_ar_ready),.auto_out_ar_valid(_axi4yank_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4yank_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4yank_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4yank_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4yank_auto_out_ar_bits_size),.auto_out_r_ready(_axi4yank_auto_out_r_ready),.auto_out_r_valid(_axi42tl_auto_in_r_valid),.auto_out_r_bits_id(_axi42tl_auto_in_r_bits_id),.auto_out_r_bits_data(_axi42tl_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi42tl_auto_in_r_bits_resp),.auto_out_r_bits_last(_axi42tl_auto_in_r_bits_last)); 
  AXI4Fragmenter axi4frag(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4frag_auto_in_aw_ready),.auto_in_aw_valid(_axi4index_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4index_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4index_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4index_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4index_auto_out_aw_bits_size),.auto_in_aw_bits_burst(_axi4index_auto_out_aw_bits_burst),.auto_in_aw_bits_echo_extra_id(_axi4index_auto_out_aw_bits_echo_extra_id),.auto_in_w_ready(_axi4frag_auto_in_w_ready),.auto_in_w_valid(_axi4index_auto_out_w_valid),.auto_in_w_bits_data(_axi4index_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4index_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4index_auto_out_w_bits_last),.auto_in_b_ready(_axi4index_auto_out_b_ready),.auto_in_b_valid(_axi4frag_auto_in_b_valid),.auto_in_b_bits_id(_axi4frag_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4frag_auto_in_b_bits_resp),.auto_in_b_bits_echo_extra_id(_axi4frag_auto_in_b_bits_echo_extra_id),.auto_in_ar_ready(_axi4frag_auto_in_ar_ready),.auto_in_ar_valid(_axi4index_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4index_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4index_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4index_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4index_auto_out_ar_bits_size),.auto_in_ar_bits_burst(_axi4index_auto_out_ar_bits_burst),.auto_in_ar_bits_echo_extra_id(_axi4index_auto_out_ar_bits_echo_extra_id),.auto_in_r_ready(_axi4index_auto_out_r_ready),.auto_in_r_valid(_axi4frag_auto_in_r_valid),.auto_in_r_bits_id(_axi4frag_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4frag_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4frag_auto_in_r_bits_resp),.auto_in_r_bits_echo_extra_id(_axi4frag_auto_in_r_bits_echo_extra_id),.auto_in_r_bits_last(_axi4frag_auto_in_r_bits_last),.auto_out_aw_ready(_axi4yank_auto_in_aw_ready),.auto_out_aw_valid(_axi4frag_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4frag_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4frag_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4frag_auto_out_aw_bits_size),.auto_out_aw_bits_echo_extra_id(_axi4frag_auto_out_aw_bits_echo_extra_id),.auto_out_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),.auto_out_w_ready(_axi4yank_auto_in_w_ready),.auto_out_w_valid(_axi4frag_auto_out_w_valid),.auto_out_w_bits_data(_axi4frag_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4frag_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4frag_auto_out_w_bits_last),.auto_out_b_ready(_axi4frag_auto_out_b_ready),.auto_out_b_valid(_axi4yank_auto_in_b_valid),.auto_out_b_bits_id(_axi4yank_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4yank_auto_in_b_bits_resp),.auto_out_b_bits_echo_extra_id(_axi4yank_auto_in_b_bits_echo_extra_id),.auto_out_b_bits_echo_real_last(_axi4yank_auto_in_b_bits_echo_real_last),.auto_out_ar_ready(_axi4yank_auto_in_ar_ready),.auto_out_ar_valid(_axi4frag_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4frag_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4frag_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4frag_auto_out_ar_bits_size),.auto_out_ar_bits_echo_extra_id(_axi4frag_auto_out_ar_bits_echo_extra_id),.auto_out_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),.auto_out_r_ready(_axi4frag_auto_out_r_ready),.auto_out_r_valid(_axi4yank_auto_in_r_valid),.auto_out_r_bits_id(_axi4yank_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4yank_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4yank_auto_in_r_bits_resp),.auto_out_r_bits_echo_extra_id(_axi4yank_auto_in_r_bits_echo_extra_id),.auto_out_r_bits_echo_real_last(_axi4yank_auto_in_r_bits_echo_real_last),.auto_out_r_bits_last(_axi4yank_auto_in_r_bits_last)); 
  AXI4IdIndexer_1 axi4index(.auto_in_aw_ready(auto_axi4index_in_aw_ready),.auto_in_aw_valid(auto_axi4index_in_aw_valid),.auto_in_aw_bits_id(auto_axi4index_in_aw_bits_id),.auto_in_aw_bits_addr(auto_axi4index_in_aw_bits_addr),.auto_in_aw_bits_len(auto_axi4index_in_aw_bits_len),.auto_in_aw_bits_size(auto_axi4index_in_aw_bits_size),.auto_in_aw_bits_burst(auto_axi4index_in_aw_bits_burst),.auto_in_w_ready(auto_axi4index_in_w_ready),.auto_in_w_valid(auto_axi4index_in_w_valid),.auto_in_w_bits_data(auto_axi4index_in_w_bits_data),.auto_in_w_bits_strb(auto_axi4index_in_w_bits_strb),.auto_in_w_bits_last(auto_axi4index_in_w_bits_last),.auto_in_b_ready(auto_axi4index_in_b_ready),.auto_in_b_valid(auto_axi4index_in_b_valid),.auto_in_b_bits_id(auto_axi4index_in_b_bits_id),.auto_in_b_bits_resp(auto_axi4index_in_b_bits_resp),.auto_in_ar_ready(auto_axi4index_in_ar_ready),.auto_in_ar_valid(auto_axi4index_in_ar_valid),.auto_in_ar_bits_id(auto_axi4index_in_ar_bits_id),.auto_in_ar_bits_addr(auto_axi4index_in_ar_bits_addr),.auto_in_ar_bits_len(auto_axi4index_in_ar_bits_len),.auto_in_ar_bits_size(auto_axi4index_in_ar_bits_size),.auto_in_ar_bits_burst(auto_axi4index_in_ar_bits_burst),.auto_in_r_ready(auto_axi4index_in_r_ready),.auto_in_r_valid(auto_axi4index_in_r_valid),.auto_in_r_bits_id(auto_axi4index_in_r_bits_id),.auto_in_r_bits_data(auto_axi4index_in_r_bits_data),.auto_in_r_bits_resp(auto_axi4index_in_r_bits_resp),.auto_in_r_bits_last(auto_axi4index_in_r_bits_last),.auto_out_aw_ready(_axi4frag_auto_in_aw_ready),.auto_out_aw_valid(_axi4index_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4index_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4index_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4index_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4index_auto_out_aw_bits_size),.auto_out_aw_bits_burst(_axi4index_auto_out_aw_bits_burst),.auto_out_aw_bits_echo_extra_id(_axi4index_auto_out_aw_bits_echo_extra_id),.auto_out_w_ready(_axi4frag_auto_in_w_ready),.auto_out_w_valid(_axi4index_auto_out_w_valid),.auto_out_w_bits_data(_axi4index_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4index_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4index_auto_out_w_bits_last),.auto_out_b_ready(_axi4index_auto_out_b_ready),.auto_out_b_valid(_axi4frag_auto_in_b_valid),.auto_out_b_bits_id(_axi4frag_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4frag_auto_in_b_bits_resp),.auto_out_b_bits_echo_extra_id(_axi4frag_auto_in_b_bits_echo_extra_id),.auto_out_ar_ready(_axi4frag_auto_in_ar_ready),.auto_out_ar_valid(_axi4index_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4index_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4index_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4index_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4index_auto_out_ar_bits_size),.auto_out_ar_bits_burst(_axi4index_auto_out_ar_bits_burst),.auto_out_ar_bits_echo_extra_id(_axi4index_auto_out_ar_bits_echo_extra_id),.auto_out_r_ready(_axi4index_auto_out_r_ready),.auto_out_r_valid(_axi4frag_auto_in_r_valid),.auto_out_r_bits_id(_axi4frag_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4frag_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4frag_auto_in_r_bits_resp),.auto_out_r_bits_echo_extra_id(_axi4frag_auto_in_r_bits_echo_extra_id),.auto_out_r_bits_last(_axi4frag_auto_in_r_bits_last)); 
endmodule
 
module FixedClockBroadcast_3 (
  input auto_in_clock,
  input auto_in_reset,
  output auto_out_3_clock,
  output auto_out_3_reset,
  output auto_out_1_clock,
  output auto_out_1_reset,
  output auto_out_0_clock,
  output auto_out_0_reset) ; 
  assign auto_out_3_clock=auto_in_clock; 
  assign auto_out_3_reset=auto_in_reset; 
  assign auto_out_1_clock=auto_in_clock; 
  assign auto_out_1_reset=auto_in_reset; 
  assign auto_out_0_clock=auto_in_clock; 
  assign auto_out_0_reset=auto_in_reset; 
endmodule
 
module TLMonitor_8 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [27:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [4:0] source ;  
   reg [27:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg sink ;  
   reg denied ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [151:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>{69'h0,io_in_d_bits_source,2'h0} ;  
   wire _GEN_0=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [151:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_1=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_2=io_in_a_bits_size<4'hD ;  
   wire _GEN_3=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_4=io_in_a_bits_address[27:12]==16'h0 ;  
   wire _GEN_5={io_in_a_bits_address[27:14],~(io_in_a_bits_address[13:12])}==16'h0 ;  
   wire _GEN_6={io_in_a_bits_address[27:17],~(io_in_a_bits_address[16])}==12'h0 ;  
   wire _GEN_7={io_in_a_bits_address[27:26],io_in_a_bits_address[25:16]^10'h200}==12'h0 ;  
   wire _GEN_8=_source_ok_T_12&io_in_a_bits_size==4'h6&_GEN_2&(_GEN_4|_GEN_5|_GEN_6|_GEN_7|(&(io_in_a_bits_address[27:26]))) ;  
   wire _GEN_9=io_in_a_bits_param>3'h2 ;  
   wire _GEN_10=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_11=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_12=_GEN_2&(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14) ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_14=_GEN_2&_GEN_5 ;  
   wire _GEN_15=io_in_a_bits_size<4'h7 ;  
   wire _GEN_16=io_in_a_bits_mask!=mask ;  
   wire _GEN_17=_GEN_12&(_GEN_14|_GEN_15&(_GEN_4|_GEN_7|(&(io_in_a_bits_address[27:26])))) ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_19=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_20=_GEN_12&io_in_a_bits_size<4'h4&_GEN_5 ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_22=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_23=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_24=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_25=io_in_d_bits_size<4'h3 ;  
   wire _GEN_26=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_27=io_in_d_bits_param==2'h2 ;  
   wire _GEN_28=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_29=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_30=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_31=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_32=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_33=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_34=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [151:0] _GEN_35={144'h0,io_in_d_bits_source,3'h0} ;  
   wire _GEN_36=io_in_d_valid&d_first_1 ;  
   wire _GEN_37=_GEN_36&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&a_first_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_38={14'h0,io_in_d_bits_source} ;  
   wire _GEN_39=_GEN_37&same_cycle_resp&~reset ;  
   wire _GEN_40=_GEN_37&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_41={4'h0,io_in_d_bits_size} ;  
   wire _GEN_42=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_43=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_44=inflight>>_GEN_38 ;  
   wire [151:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_35 ;  
   wire [18:0] _GEN_45=inflight_1>>_GEN_38 ;  
   wire [151:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_35 ;  
  always @( posedge clock)
       begin 
         if (_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~(_GEN_14|_GEN_15&(_GEN_4|_GEN_6|_GEN_7|(&(io_in_a_bits_address[27:26])))))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~(_GEN_12&_GEN_14))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&_GEN_43[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~reset&~(_GEN_44[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_41!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~(_GEN_45[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_41!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:54:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_46={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_46 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_46 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_46 ;  
   wire [31:0] _GEN_47={27'h0,io_in_d_bits_source} ;  
   wire [270:0] _GEN_48={263'h0,io_in_d_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_47 ;  
   wire [31:0] _a_set_T=32'h1<<io_in_a_bits_source ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<{264'h0,io_in_d_bits_source,2'h0} ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_0 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _d_sizes_clr_T_5=271'hFF<<_GEN_48 ;  
   wire [259:0] _a_sizes_set_T_1={255'h0,_GEN_0 ? {io_in_a_bits_size,1'h1}:5'h0}<<{252'h0,io_in_a_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_47 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hFF<<_GEN_48 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_49=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_50=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=152'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=152'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_0 ? _a_set_T[18:0]:19'h0))&~(_GEN_49 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_0 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_49 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_0 ? _a_sizes_set_T_1[151:0]:152'h0))&~(_GEN_49 ? _d_sizes_clr_T_5[151:0]:152'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_50 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_50 ? _d_sizes_clr_T_11[151:0]:152'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLFIFOFixer_3 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [27:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [4:0] auto_out_a_bits_source,
  output [27:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [4:0] auto_out_d_bits_source,
  input auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   wire [2:0] a_id={{auto_in_a_bits_address[27],auto_in_a_bits_address[25],auto_in_a_bits_address[16],auto_in_a_bits_address[13]}==4'h0,{auto_in_a_bits_address[27],{auto_in_a_bits_address[27],auto_in_a_bits_address[25],auto_in_a_bits_address[16],~(auto_in_a_bits_address[13])}==4'h0}|{2{{auto_in_a_bits_address[27],~(auto_in_a_bits_address[25]),auto_in_a_bits_address[16]}==3'h0}}}|({auto_in_a_bits_address[27],auto_in_a_bits_address[25],~(auto_in_a_bits_address[16])}==3'h0 ? 3'h5:3'h0) ;  
   wire a_noDomain=a_id==3'h0 ;  
   reg [8:0] a_first_counter ;  
   wire a_first=a_first_counter==9'h0 ;  
   reg [8:0] d_first_counter ;  
   reg flight_0 ;  
   reg flight_1 ;  
   reg flight_2 ;  
   reg flight_3 ;  
   reg flight_4 ;  
   reg flight_5 ;  
   reg flight_6 ;  
   reg flight_7 ;  
   reg flight_8 ;  
   reg flight_9 ;  
   reg flight_10 ;  
   reg flight_11 ;  
   reg flight_12 ;  
   reg flight_13 ;  
   reg flight_14 ;  
   reg flight_15 ;  
   wire stalls_a_sel=auto_in_a_bits_source[4:3]==2'h0 ;  
   reg [2:0] stalls_id ;  
   wire stalls_a_sel_1=auto_in_a_bits_source[4:3]==2'h1 ;  
   reg [2:0] stalls_id_1 ;  
   wire stall=stalls_a_sel&a_first&(flight_0|flight_1|flight_2|flight_3|flight_4|flight_5|flight_6|flight_7)&(a_noDomain|stalls_id!=a_id)|stalls_a_sel_1&a_first&(flight_8|flight_9|flight_10|flight_11|flight_12|flight_13|flight_14|flight_15)&(a_noDomain|stalls_id_1!=a_id) ;  
   wire nodeIn_a_ready=auto_out_a_ready&~stall ;  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<auto_in_a_bits_size ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<auto_out_d_bits_size ;  
   wire d_first_first=d_first_counter==9'h0 ;  
   wire _GEN=d_first_first&auto_out_d_bits_opcode!=3'h6&auto_in_d_ready&auto_out_d_valid ;  
   wire _stalls_id_T_4=nodeIn_a_ready&auto_in_a_valid ;  
   wire _GEN_0=a_first&_stalls_id_T_4 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              flight_0 <=1'h0;
              flight_1 <=1'h0;
              flight_2 <=1'h0;
              flight_3 <=1'h0;
              flight_4 <=1'h0;
              flight_5 <=1'h0;
              flight_6 <=1'h0;
              flight_7 <=1'h0;
              flight_8 <=1'h0;
              flight_9 <=1'h0;
              flight_10 <=1'h0;
              flight_11 <=1'h0;
              flight_12 <=1'h0;
              flight_13 <=1'h0;
              flight_14 <=1'h0;
              flight_15 <=1'h0;
            end 
          else 
            begin 
              if (_stalls_id_T_4)
                 begin 
                   if (a_first)
                      a_first_counter <=auto_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                    else 
                      a_first_counter <=a_first_counter-9'h1;
                 end 
              if (auto_in_d_ready&auto_out_d_valid)
                 begin 
                   if (d_first_first)
                      d_first_counter <=auto_out_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                    else 
                      d_first_counter <=d_first_counter-9'h1;
                 end 
              flight_0 <=~(_GEN&auto_out_d_bits_source==5'h0)&(_GEN_0&auto_in_a_bits_source==5'h0|flight_0);
              flight_1 <=~(_GEN&auto_out_d_bits_source==5'h1)&(_GEN_0&auto_in_a_bits_source==5'h1|flight_1);
              flight_2 <=~(_GEN&auto_out_d_bits_source==5'h2)&(_GEN_0&auto_in_a_bits_source==5'h2|flight_2);
              flight_3 <=~(_GEN&auto_out_d_bits_source==5'h3)&(_GEN_0&auto_in_a_bits_source==5'h3|flight_3);
              flight_4 <=~(_GEN&auto_out_d_bits_source==5'h4)&(_GEN_0&auto_in_a_bits_source==5'h4|flight_4);
              flight_5 <=~(_GEN&auto_out_d_bits_source==5'h5)&(_GEN_0&auto_in_a_bits_source==5'h5|flight_5);
              flight_6 <=~(_GEN&auto_out_d_bits_source==5'h6)&(_GEN_0&auto_in_a_bits_source==5'h6|flight_6);
              flight_7 <=~(_GEN&auto_out_d_bits_source==5'h7)&(_GEN_0&auto_in_a_bits_source==5'h7|flight_7);
              flight_8 <=~(_GEN&auto_out_d_bits_source==5'h8)&(_GEN_0&auto_in_a_bits_source==5'h8|flight_8);
              flight_9 <=~(_GEN&auto_out_d_bits_source==5'h9)&(_GEN_0&auto_in_a_bits_source==5'h9|flight_9);
              flight_10 <=~(_GEN&auto_out_d_bits_source==5'hA)&(_GEN_0&auto_in_a_bits_source==5'hA|flight_10);
              flight_11 <=~(_GEN&auto_out_d_bits_source==5'hB)&(_GEN_0&auto_in_a_bits_source==5'hB|flight_11);
              flight_12 <=~(_GEN&auto_out_d_bits_source==5'hC)&(_GEN_0&auto_in_a_bits_source==5'hC|flight_12);
              flight_13 <=~(_GEN&auto_out_d_bits_source==5'hD)&(_GEN_0&auto_in_a_bits_source==5'hD|flight_13);
              flight_14 <=~(_GEN&auto_out_d_bits_source==5'hE)&(_GEN_0&auto_in_a_bits_source==5'hE|flight_14);
              flight_15 <=~(_GEN&auto_out_d_bits_source==5'hF)&(_GEN_0&auto_in_a_bits_source==5'hF|flight_15);
            end 
         if (_stalls_id_T_4&stalls_a_sel)
            stalls_id <=a_id;
         if (_stalls_id_T_4&stalls_a_sel_1)
            stalls_id_1 <=a_id;
       end
  
  TLMonitor_8 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_out_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_param(auto_out_d_bits_param),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source),.io_in_d_bits_sink(auto_out_d_bits_sink),.io_in_d_bits_denied(auto_out_d_bits_denied),.io_in_d_bits_corrupt(auto_out_d_bits_corrupt)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_d_valid=auto_out_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_param=auto_out_d_bits_param; 
  assign auto_in_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source; 
  assign auto_in_d_bits_sink=auto_out_d_bits_sink; 
  assign auto_in_d_bits_denied=auto_out_d_bits_denied; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign auto_out_a_valid=auto_in_a_valid&~stall; 
  assign auto_out_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_a_bits_size=auto_in_a_bits_size; 
  assign auto_out_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_a_bits_corrupt=auto_in_a_bits_corrupt; 
  assign auto_out_d_ready=auto_in_d_ready; 
endmodule
 
module TLMonitor_9 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [27:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [4:0] source ;  
   reg [27:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg sink ;  
   reg denied ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [151:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>{69'h0,io_in_d_bits_source,2'h0} ;  
   wire _GEN_0=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [151:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_1=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_2=io_in_a_bits_size<4'hD ;  
   wire _GEN_3=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_4=io_in_a_bits_address[27:12]==16'h0 ;  
   wire _GEN_5={io_in_a_bits_address[27:14],~(io_in_a_bits_address[13:12])}==16'h0 ;  
   wire _GEN_6={io_in_a_bits_address[27:17],~(io_in_a_bits_address[16])}==12'h0 ;  
   wire _GEN_7={io_in_a_bits_address[27:26],io_in_a_bits_address[25:16]^10'h200}==12'h0 ;  
   wire _GEN_8=_source_ok_T_12&io_in_a_bits_size==4'h6&_GEN_2&(_GEN_4|_GEN_5|_GEN_6|_GEN_7|(&(io_in_a_bits_address[27:26]))) ;  
   wire _GEN_9=io_in_a_bits_param>3'h2 ;  
   wire _GEN_10=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_11=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_12=_GEN_2&(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14) ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_14=_GEN_2&_GEN_5 ;  
   wire _GEN_15=io_in_a_bits_size<4'h7 ;  
   wire _GEN_16=io_in_a_bits_mask!=mask ;  
   wire _GEN_17=_GEN_12&(_GEN_14|_GEN_15&(_GEN_4|_GEN_7|(&(io_in_a_bits_address[27:26])))) ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_19=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_20=_GEN_12&io_in_a_bits_size<4'h4&_GEN_5 ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_22=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_23=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_24=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_25=io_in_d_bits_size<4'h3 ;  
   wire _GEN_26=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_27=io_in_d_bits_param==2'h2 ;  
   wire _GEN_28=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_29=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_30=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_31=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_32=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_33=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_34=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [151:0] _GEN_35={144'h0,io_in_d_bits_source,3'h0} ;  
   wire _GEN_36=io_in_d_valid&d_first_1 ;  
   wire _GEN_37=_GEN_36&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&a_first_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_38={14'h0,io_in_d_bits_source} ;  
   wire _GEN_39=_GEN_37&same_cycle_resp&~reset ;  
   wire _GEN_40=_GEN_37&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_41={4'h0,io_in_d_bits_size} ;  
   wire _GEN_42=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_43=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_44=inflight>>_GEN_38 ;  
   wire [151:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_35 ;  
   wire [18:0] _GEN_45=inflight_1>>_GEN_38 ;  
   wire [151:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_35 ;  
  always @( posedge clock)
       begin 
         if (_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~(_GEN_14|_GEN_15&(_GEN_4|_GEN_6|_GEN_7|(&(io_in_a_bits_address[27:26])))))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~(_GEN_12&_GEN_14))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&_GEN_43[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~reset&~(_GEN_44[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_41!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~(_GEN_45[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_41!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:53:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_46={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_46 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_46 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_46 ;  
   wire [31:0] _GEN_47={27'h0,io_in_d_bits_source} ;  
   wire [270:0] _GEN_48={263'h0,io_in_d_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_47 ;  
   wire [31:0] _a_set_T=32'h1<<io_in_a_bits_source ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<{264'h0,io_in_d_bits_source,2'h0} ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_0 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _d_sizes_clr_T_5=271'hFF<<_GEN_48 ;  
   wire [259:0] _a_sizes_set_T_1={255'h0,_GEN_0 ? {io_in_a_bits_size,1'h1}:5'h0}<<{252'h0,io_in_a_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_47 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hFF<<_GEN_48 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_49=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_50=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=152'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=152'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_0 ? _a_set_T[18:0]:19'h0))&~(_GEN_49 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_0 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_49 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_0 ? _a_sizes_set_T_1[151:0]:152'h0))&~(_GEN_49 ? _d_sizes_clr_T_5[151:0]:152'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_50 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_50 ? _d_sizes_clr_T_11[151:0]:152'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLXbar_5 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [27:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_4_a_ready,
  output auto_out_4_a_valid,
  output [2:0] auto_out_4_a_bits_opcode,
  output [2:0] auto_out_4_a_bits_param,
  output [2:0] auto_out_4_a_bits_size,
  output [4:0] auto_out_4_a_bits_source,
  output [16:0] auto_out_4_a_bits_address,
  output [7:0] auto_out_4_a_bits_mask,
  output auto_out_4_a_bits_corrupt,
  output auto_out_4_d_ready,
  input auto_out_4_d_valid,
  input [2:0] auto_out_4_d_bits_size,
  input [4:0] auto_out_4_d_bits_source,
  input [63:0] auto_out_4_d_bits_data,
  input auto_out_3_a_ready,
  output auto_out_3_a_valid,
  output [2:0] auto_out_3_a_bits_opcode,
  output [2:0] auto_out_3_a_bits_param,
  output [2:0] auto_out_3_a_bits_size,
  output [4:0] auto_out_3_a_bits_source,
  output [11:0] auto_out_3_a_bits_address,
  output [7:0] auto_out_3_a_bits_mask,
  output [63:0] auto_out_3_a_bits_data,
  output auto_out_3_a_bits_corrupt,
  output auto_out_3_d_ready,
  input auto_out_3_d_valid,
  input [2:0] auto_out_3_d_bits_opcode,
  input [2:0] auto_out_3_d_bits_size,
  input [4:0] auto_out_3_d_bits_source,
  input [63:0] auto_out_3_d_bits_data,
  input auto_out_2_a_ready,
  output auto_out_2_a_valid,
  output [2:0] auto_out_2_a_bits_opcode,
  output [2:0] auto_out_2_a_bits_param,
  output [2:0] auto_out_2_a_bits_size,
  output [4:0] auto_out_2_a_bits_source,
  output [25:0] auto_out_2_a_bits_address,
  output [7:0] auto_out_2_a_bits_mask,
  output [63:0] auto_out_2_a_bits_data,
  output auto_out_2_a_bits_corrupt,
  output auto_out_2_d_ready,
  input auto_out_2_d_valid,
  input [2:0] auto_out_2_d_bits_opcode,
  input [2:0] auto_out_2_d_bits_size,
  input [4:0] auto_out_2_d_bits_source,
  input [63:0] auto_out_2_d_bits_data,
  input auto_out_1_a_ready,
  output auto_out_1_a_valid,
  output [2:0] auto_out_1_a_bits_opcode,
  output [2:0] auto_out_1_a_bits_param,
  output [2:0] auto_out_1_a_bits_size,
  output [4:0] auto_out_1_a_bits_source,
  output [27:0] auto_out_1_a_bits_address,
  output [7:0] auto_out_1_a_bits_mask,
  output [63:0] auto_out_1_a_bits_data,
  output auto_out_1_a_bits_corrupt,
  output auto_out_1_d_ready,
  input auto_out_1_d_valid,
  input [2:0] auto_out_1_d_bits_opcode,
  input [2:0] auto_out_1_d_bits_size,
  input [4:0] auto_out_1_d_bits_source,
  input [63:0] auto_out_1_d_bits_data,
  input auto_out_0_a_ready,
  output auto_out_0_a_valid,
  output [2:0] auto_out_0_a_bits_opcode,
  output [2:0] auto_out_0_a_bits_param,
  output [3:0] auto_out_0_a_bits_size,
  output [4:0] auto_out_0_a_bits_source,
  output [13:0] auto_out_0_a_bits_address,
  output [7:0] auto_out_0_a_bits_mask,
  output auto_out_0_a_bits_corrupt,
  output auto_out_0_d_ready,
  input auto_out_0_d_valid,
  input [2:0] auto_out_0_d_bits_opcode,
  input [1:0] auto_out_0_d_bits_param,
  input [3:0] auto_out_0_d_bits_size,
  input [4:0] auto_out_0_d_bits_source,
  input auto_out_0_d_bits_sink,
  input auto_out_0_d_bits_denied,
  input [63:0] auto_out_0_d_bits_data,
  input auto_out_0_d_bits_corrupt) ; 
   wire requestAIO_0_0={auto_in_a_bits_address[27],auto_in_a_bits_address[25],auto_in_a_bits_address[16],~(auto_in_a_bits_address[13])}==4'h0 ;  
   wire requestAIO_0_2={auto_in_a_bits_address[27],~(auto_in_a_bits_address[25]),auto_in_a_bits_address[16]}==3'h0 ;  
   wire requestAIO_0_3={auto_in_a_bits_address[27],auto_in_a_bits_address[25],auto_in_a_bits_address[16],auto_in_a_bits_address[13]}==4'h0 ;  
   wire requestAIO_0_4={auto_in_a_bits_address[27],auto_in_a_bits_address[25],~(auto_in_a_bits_address[16])}==3'h0 ;  
   wire _portsAOI_in_0_a_ready_T_8=requestAIO_0_0&auto_out_0_a_ready|auto_in_a_bits_address[27]&auto_out_1_a_ready|requestAIO_0_2&auto_out_2_a_ready|requestAIO_0_3&auto_out_3_a_ready|requestAIO_0_4&auto_out_4_a_ready ;  
   reg [8:0] beatsLeft ;  
   wire idle=beatsLeft==9'h0 ;  
   wire [4:0] readys_valid={auto_out_4_d_valid,auto_out_3_d_valid,auto_out_2_d_valid,auto_out_1_d_valid,auto_out_0_d_valid} ;  
   reg [4:0] readys_mask ;  
   wire [4:0] _readys_filter_T_1=readys_valid&~readys_mask ;  
   wire [7:0] _GEN={_readys_filter_T_1[3:0],auto_out_4_d_valid,auto_out_3_d_valid,auto_out_2_d_valid,auto_out_1_d_valid}|{_readys_filter_T_1,auto_out_4_d_valid,auto_out_3_d_valid,auto_out_2_d_valid} ;  
   wire [6:0] _GEN_0=_GEN[6:0]|{_readys_filter_T_1[4],_GEN[7:2]} ;  
   wire [4:0] readys_readys=~({readys_mask[4],_readys_filter_T_1[4]|readys_mask[3],_GEN[7]|readys_mask[2],_GEN_0[6:5]|readys_mask[1:0]}&(_GEN_0[4:0]|{_readys_filter_T_1[4],_GEN[7],_GEN_0[6:4]})) ;  
   wire winner_0=readys_readys[0]&auto_out_0_d_valid ;  
   wire winner_1=readys_readys[1]&auto_out_1_d_valid ;  
   wire winner_2=readys_readys[2]&auto_out_2_d_valid ;  
   wire winner_3=readys_readys[3]&auto_out_3_d_valid ;  
   wire winner_4=readys_readys[4]&auto_out_4_d_valid ;  
   wire _in_0_d_valid_T=auto_out_0_d_valid|auto_out_1_d_valid ;  
   wire prefixOR_2=winner_0|winner_1 ;  
   wire prefixOR_3=prefixOR_2|winner_2 ;  
  always @( posedge clock)
       begin 
         if (~reset&~((~winner_0|~winner_1)&(~prefixOR_2|~winner_2)&(~prefixOR_3|~winner_3)&(~(prefixOR_3|winner_3)|~winner_4)))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~(_in_0_d_valid_T|auto_out_2_d_valid|auto_out_3_d_valid|auto_out_4_d_valid)|winner_0|winner_1|winner_2|winner_3|winner_4))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg state_0 ;  
   reg state_1 ;  
   reg state_2 ;  
   reg state_3 ;  
   reg state_4 ;  
   wire muxState_0=idle ? winner_0:state_0 ;  
   wire muxState_1=idle ? winner_1:state_1 ;  
   wire muxState_2=idle ? winner_2:state_2 ;  
   wire muxState_3=idle ? winner_3:state_3 ;  
   wire muxState_4=idle ? winner_4:state_4 ;  
   wire in_0_d_valid=idle ? _in_0_d_valid_T|auto_out_2_d_valid|auto_out_3_d_valid|auto_out_4_d_valid:state_0&auto_out_0_d_valid|state_1&auto_out_1_d_valid|state_2&auto_out_2_d_valid|state_3&auto_out_3_d_valid|state_4&auto_out_4_d_valid ;  
   wire _in_0_d_bits_T=muxState_0&auto_out_0_d_bits_corrupt ;  
   wire _in_0_d_bits_T_18=muxState_0&auto_out_0_d_bits_denied ;  
   wire _in_0_d_bits_T_27=muxState_0&auto_out_0_d_bits_sink ;  
   wire [4:0] _in_0_d_bits_T_44=(muxState_0 ? auto_out_0_d_bits_source:5'h0)|(muxState_1 ? auto_out_1_d_bits_source:5'h0)|(muxState_2 ? auto_out_2_d_bits_source:5'h0)|(muxState_3 ? auto_out_3_d_bits_source:5'h0)|(muxState_4 ? auto_out_4_d_bits_source:5'h0) ;  
   wire [3:0] _in_0_d_bits_T_53=(muxState_0 ? auto_out_0_d_bits_size:4'h0)|(muxState_1 ? {1'h0,auto_out_1_d_bits_size}:4'h0)|(muxState_2 ? {1'h0,auto_out_2_d_bits_size}:4'h0)|(muxState_3 ? {1'h0,auto_out_3_d_bits_size}:4'h0)|(muxState_4 ? {1'h0,auto_out_4_d_bits_size}:4'h0) ;  
   wire [1:0] _in_0_d_bits_T_54=muxState_0 ? auto_out_0_d_bits_param:2'h0 ;  
   wire [2:0] _in_0_d_bits_T_71=(muxState_0 ? auto_out_0_d_bits_opcode:3'h0)|(muxState_1 ? auto_out_1_d_bits_opcode:3'h0)|(muxState_2 ? auto_out_2_d_bits_opcode:3'h0)|(muxState_3 ? auto_out_3_d_bits_opcode:3'h0)|{2'h0,muxState_4} ;  
   wire [26:0] _beatsDO_decode_T_1=27'hFFF<<auto_out_0_d_bits_size ;  
   wire [8:0] maskedBeats_0=winner_0&auto_out_0_d_bits_opcode[0] ? ~(_beatsDO_decode_T_1[11:3]):9'h0 ;  
   wire [20:0] _beatsDO_decode_T_17=21'h3F<<auto_out_4_d_bits_size ;  
   wire [20:0] _beatsDO_decode_T_13=21'h3F<<auto_out_3_d_bits_size ;  
   wire [20:0] _beatsDO_decode_T_9=21'h3F<<auto_out_2_d_bits_size ;  
   wire [20:0] _beatsDO_decode_T_5=21'h3F<<auto_out_1_d_bits_size ;  
   wire [4:0] _readys_mask_T=readys_readys&readys_valid ;  
   wire [4:0] _readys_mask_T_3=_readys_mask_T|{_readys_mask_T[3:0],1'h0} ;  
   wire [4:0] _readys_mask_T_6=_readys_mask_T_3|{_readys_mask_T_3[2:0],2'h0} ;  
   wire latch=idle&auto_in_d_ready ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              beatsLeft <=9'h0;
              readys_mask <=5'h1F;
              state_0 <=1'h0;
              state_1 <=1'h0;
              state_2 <=1'h0;
              state_3 <=1'h0;
              state_4 <=1'h0;
            end 
          else 
            begin 
              if (latch)
                 beatsLeft <={maskedBeats_0[8:3],maskedBeats_0[2:0]|(winner_1&auto_out_1_d_bits_opcode[0] ? ~(_beatsDO_decode_T_5[5:3]):3'h0)|(winner_2&auto_out_2_d_bits_opcode[0] ? ~(_beatsDO_decode_T_9[5:3]):3'h0)|(winner_3&auto_out_3_d_bits_opcode[0] ? ~(_beatsDO_decode_T_13[5:3]):3'h0)|(winner_4 ? ~(_beatsDO_decode_T_17[5:3]):3'h0)};
               else 
                 beatsLeft <=beatsLeft-{8'h0,auto_in_d_ready&in_0_d_valid};
              if (latch&(|readys_valid))
                 readys_mask <=_readys_mask_T_6|{_readys_mask_T_6[0],4'h0};
              if (idle)
                 begin 
                   state_0 <=winner_0;
                   state_1 <=winner_1;
                   state_2 <=winner_2;
                   state_3 <=winner_3;
                   state_4 <=winner_4;
                 end 
            end 
       end
  
  TLMonitor_9 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_portsAOI_in_0_a_ready_T_8),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(in_0_d_valid),.io_in_d_bits_opcode(_in_0_d_bits_T_71),.io_in_d_bits_param(_in_0_d_bits_T_54),.io_in_d_bits_size(_in_0_d_bits_T_53),.io_in_d_bits_source(_in_0_d_bits_T_44),.io_in_d_bits_sink(_in_0_d_bits_T_27),.io_in_d_bits_denied(_in_0_d_bits_T_18),.io_in_d_bits_corrupt(_in_0_d_bits_T)); 
  assign auto_in_a_ready=_portsAOI_in_0_a_ready_T_8; 
  assign auto_in_d_valid=in_0_d_valid; 
  assign auto_in_d_bits_opcode=_in_0_d_bits_T_71; 
  assign auto_in_d_bits_param=_in_0_d_bits_T_54; 
  assign auto_in_d_bits_size=_in_0_d_bits_T_53; 
  assign auto_in_d_bits_source=_in_0_d_bits_T_44; 
  assign auto_in_d_bits_sink=_in_0_d_bits_T_27; 
  assign auto_in_d_bits_denied=_in_0_d_bits_T_18; 
  assign auto_in_d_bits_data=(muxState_0 ? auto_out_0_d_bits_data:64'h0)|(muxState_1 ? auto_out_1_d_bits_data:64'h0)|(muxState_2 ? auto_out_2_d_bits_data:64'h0)|(muxState_3 ? auto_out_3_d_bits_data:64'h0)|(muxState_4 ? auto_out_4_d_bits_data:64'h0); 
  assign auto_in_d_bits_corrupt=_in_0_d_bits_T; 
  assign auto_out_4_a_valid=auto_in_a_valid&requestAIO_0_4; 
  assign auto_out_4_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_4_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_4_a_bits_size=auto_in_a_bits_size[2:0]; 
  assign auto_out_4_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_4_a_bits_address=auto_in_a_bits_address[16:0]; 
  assign auto_out_4_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_4_a_bits_corrupt=auto_in_a_bits_corrupt; 
  assign auto_out_4_d_ready=auto_in_d_ready&(idle ? readys_readys[4]:state_4); 
  assign auto_out_3_a_valid=auto_in_a_valid&requestAIO_0_3; 
  assign auto_out_3_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_3_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_3_a_bits_size=auto_in_a_bits_size[2:0]; 
  assign auto_out_3_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_3_a_bits_address=auto_in_a_bits_address[11:0]; 
  assign auto_out_3_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_3_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_3_a_bits_corrupt=auto_in_a_bits_corrupt; 
  assign auto_out_3_d_ready=auto_in_d_ready&(idle ? readys_readys[3]:state_3); 
  assign auto_out_2_a_valid=auto_in_a_valid&requestAIO_0_2; 
  assign auto_out_2_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_2_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_2_a_bits_size=auto_in_a_bits_size[2:0]; 
  assign auto_out_2_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_2_a_bits_address=auto_in_a_bits_address[25:0]; 
  assign auto_out_2_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_2_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_2_a_bits_corrupt=auto_in_a_bits_corrupt; 
  assign auto_out_2_d_ready=auto_in_d_ready&(idle ? readys_readys[2]:state_2); 
  assign auto_out_1_a_valid=auto_in_a_valid&auto_in_a_bits_address[27]; 
  assign auto_out_1_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_1_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_1_a_bits_size=auto_in_a_bits_size[2:0]; 
  assign auto_out_1_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_1_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_1_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_1_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_1_a_bits_corrupt=auto_in_a_bits_corrupt; 
  assign auto_out_1_d_ready=auto_in_d_ready&(idle ? readys_readys[1]:state_1); 
  assign auto_out_0_a_valid=auto_in_a_valid&requestAIO_0_0; 
  assign auto_out_0_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_0_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_0_a_bits_size=auto_in_a_bits_size; 
  assign auto_out_0_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_0_a_bits_address=auto_in_a_bits_address[13:0]; 
  assign auto_out_0_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_0_a_bits_corrupt=auto_in_a_bits_corrupt; 
  assign auto_out_0_d_ready=auto_in_d_ready&(idle ? readys_readys[0]:state_0); 
endmodule
 
module TLMonitor_10 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [27:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [4:0] source ;  
   reg [27:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg sink ;  
   reg denied ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [151:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>{69'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _GEN_0={27'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [31:0] _GEN_2={27'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [151:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_a_bits_address[27:12]==16'h0 ;  
   wire _GEN_7={io_in_a_bits_address[27:14],~(io_in_a_bits_address[13:12])}==16'h0 ;  
   wire _GEN_8={io_in_a_bits_address[27:17],~(io_in_a_bits_address[16])}==12'h0 ;  
   wire _GEN_9={io_in_a_bits_address[27:26],io_in_a_bits_address[25:16]^10'h200}==12'h0 ;  
   wire _GEN_10=_source_ok_T_12&io_in_a_bits_size==4'h6&_GEN_4&(_GEN_6|_GEN_7|_GEN_8|_GEN_9|(&(io_in_a_bits_address[27:26]))) ;  
   wire _GEN_11=io_in_a_bits_param>3'h2 ;  
   wire _GEN_12=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_13=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_14=_GEN_4&(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14) ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_16=_GEN_4&_GEN_7 ;  
   wire _GEN_17=io_in_a_bits_size<4'h7 ;  
   wire _GEN_18=io_in_a_bits_mask!=mask ;  
   wire _GEN_19=_GEN_14&(_GEN_16|_GEN_17&(_GEN_6|_GEN_9|(&(io_in_a_bits_address[27:26])))) ;  
   wire _GEN_20=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_22=_GEN_14&io_in_a_bits_size<4'h4&_GEN_7 ;  
   wire _GEN_23=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_26=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_27=io_in_d_bits_size<4'h3 ;  
   wire _GEN_28=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_29=io_in_d_bits_param==2'h2 ;  
   wire _GEN_30=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_31=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_32=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_33=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_35=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_36=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [151:0] _GEN_37={144'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [31:0] _a_set_wo_ready_T=32'h1<<_GEN_0 ;  
   wire [18:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_38=io_in_d_valid&d_first_1 ;  
   wire _GEN_39=_GEN_38&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_40={14'h0,io_in_d_bits_source} ;  
   wire _GEN_41=_GEN_39&same_cycle_resp&~reset ;  
   wire _GEN_42=_GEN_39&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_43={4'h0,io_in_d_bits_size} ;  
   wire _GEN_44=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_45=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_46=inflight>>_GEN_40 ;  
   wire [151:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_37 ;  
   wire [31:0] _d_clr_wo_ready_T=32'h1<<_GEN_2 ;  
   wire [18:0] _GEN_47=inflight_1>>_GEN_40 ;  
   wire [151:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_37 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~(_GEN_16|_GEN_17&(_GEN_6|_GEN_8|_GEN_9|(&(io_in_a_bits_address[27:26])))))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~(_GEN_14&_GEN_16))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_45[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&~reset&~(_GEN_46[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_43!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_39 ? _d_clr_wo_ready_T[18:0]:19'h0)|a_set_wo_ready==19'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 2 (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~(_GEN_47[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&_GEN_43!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:55:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_48={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_48 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_48 ;  
   wire [270:0] _GEN_49={263'h0,io_in_d_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_2 ;  
   wire [31:0] _a_set_T=32'h1<<_GEN_0 ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<{264'h0,io_in_d_bits_source,2'h0} ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _d_sizes_clr_T_5=271'hFF<<_GEN_49 ;  
   wire [259:0] _a_sizes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{252'h0,io_in_a_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_2 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hFF<<_GEN_49 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_50=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_51=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=152'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=152'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[18:0]:19'h0))&~(_GEN_50 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_50 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[151:0]:152'h0))&~(_GEN_50 ? _d_sizes_clr_T_5[151:0]:152'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_51 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_51 ? _d_sizes_clr_T_11[151:0]:152'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module ram_source_2x5 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [4:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [4:0] W0_data) ; 
   reg [4:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:5'bx; 
endmodule
 
module ram_address_2x28 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [27:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [27:0] W0_data) ; 
   reg [27:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:28'bx; 
endmodule
 
module Queue_35 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input [27:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input [63:0] io_enq_bits_data,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source,
  output [27:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x3 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_source_2x5 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_address_2x28 ram_address_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_address),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_address)); 
  ram_2x8 ram_mask_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_mask),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_mask)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_corrupt)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_36 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [1:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input io_enq_bits_sink,
  input io_enq_bits_denied,
  input [63:0] io_enq_bits_data,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [1:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source,
  output io_deq_bits_sink,
  output io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x2 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_source_2x5 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_2x1 ram_sink_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_sink),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_sink)); 
  ram_2x1 ram_denied_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_denied),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_denied)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_corrupt)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module TLBuffer_4 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [27:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [4:0] auto_out_a_bits_source,
  output [27:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [4:0] auto_out_d_bits_source,
  input auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   wire _nodeIn_d_q_io_deq_valid ;  
   wire [2:0] _nodeIn_d_q_io_deq_bits_opcode ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_param ;  
   wire [3:0] _nodeIn_d_q_io_deq_bits_size ;  
   wire [4:0] _nodeIn_d_q_io_deq_bits_source ;  
   wire _nodeIn_d_q_io_deq_bits_sink ;  
   wire _nodeIn_d_q_io_deq_bits_denied ;  
   wire _nodeIn_d_q_io_deq_bits_corrupt ;  
   wire _nodeOut_a_q_io_enq_ready ;  
  TLMonitor_10 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_nodeOut_a_q_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(_nodeIn_d_q_io_deq_valid),.io_in_d_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_in_d_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_in_d_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_in_d_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_in_d_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_in_d_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_in_d_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  Queue_35 nodeOut_a_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_a_q_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_data(auto_in_a_bits_data),.io_enq_bits_corrupt(auto_in_a_bits_corrupt),.io_deq_ready(auto_out_a_ready),.io_deq_valid(auto_out_a_valid),.io_deq_bits_opcode(auto_out_a_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(auto_out_a_bits_size),.io_deq_bits_source(auto_out_a_bits_source),.io_deq_bits_address(auto_out_a_bits_address),.io_deq_bits_mask(auto_out_a_bits_mask),.io_deq_bits_data(auto_out_a_bits_data),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  Queue_36 nodeIn_d_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_d_ready),.io_enq_valid(auto_out_d_valid),.io_enq_bits_opcode(auto_out_d_bits_opcode),.io_enq_bits_param(auto_out_d_bits_param),.io_enq_bits_size(auto_out_d_bits_size),.io_enq_bits_source(auto_out_d_bits_source),.io_enq_bits_sink(auto_out_d_bits_sink),.io_enq_bits_denied(auto_out_d_bits_denied),.io_enq_bits_data(auto_out_d_bits_data),.io_enq_bits_corrupt(auto_out_d_bits_corrupt),.io_deq_ready(auto_in_d_ready),.io_deq_valid(_nodeIn_d_q_io_deq_valid),.io_deq_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_deq_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_deq_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_deq_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_deq_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_deq_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_deq_bits_data(auto_in_d_bits_data),.io_deq_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  assign auto_in_a_ready=_nodeOut_a_q_io_enq_ready; 
  assign auto_in_d_valid=_nodeIn_d_q_io_deq_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_q_io_deq_bits_opcode; 
  assign auto_in_d_bits_param=_nodeIn_d_q_io_deq_bits_param; 
  assign auto_in_d_bits_size=_nodeIn_d_q_io_deq_bits_size; 
  assign auto_in_d_bits_source=_nodeIn_d_q_io_deq_bits_source; 
  assign auto_in_d_bits_sink=_nodeIn_d_q_io_deq_bits_sink; 
  assign auto_in_d_bits_denied=_nodeIn_d_q_io_deq_bits_denied; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_q_io_deq_bits_corrupt; 
endmodule
 
module TLMonitor_11 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [27:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [4:0] source ;  
   reg [27:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg sink ;  
   reg denied ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [151:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>{69'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _GEN_0={27'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [31:0] _GEN_2={27'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [151:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_a_bits_address[27:12]==16'h0 ;  
   wire _GEN_7={io_in_a_bits_address[27:14],~(io_in_a_bits_address[13:12])}==16'h0 ;  
   wire _GEN_8={io_in_a_bits_address[27:17],~(io_in_a_bits_address[16])}==12'h0 ;  
   wire _GEN_9={io_in_a_bits_address[27:26],io_in_a_bits_address[25:16]^10'h200}==12'h0 ;  
   wire _GEN_10=_GEN_6|_GEN_7 ;  
   wire _GEN_11=_source_ok_T_12&io_in_a_bits_size==4'h6&_GEN_4&(_GEN_10|_GEN_8|_GEN_9|(&(io_in_a_bits_address[27:26]))) ;  
   wire _GEN_12=io_in_a_bits_param>3'h2 ;  
   wire _GEN_13=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_14=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_15=_GEN_4&(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14) ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_17=_GEN_4&_GEN_7 ;  
   wire _GEN_18=io_in_a_bits_size<4'h7 ;  
   wire _GEN_19=io_in_a_bits_mask!=mask ;  
   wire _GEN_20=_GEN_15&(_GEN_17|_GEN_18&(_GEN_6|_GEN_9|(&(io_in_a_bits_address[27:26])))) ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_22=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_23=_GEN_15&io_in_a_bits_size<4'h4&(_GEN_10|_GEN_9|(&(io_in_a_bits_address[27:26]))) ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_26=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_27=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_28=io_in_d_bits_size<4'h3 ;  
   wire _GEN_29=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_30=io_in_d_bits_param==2'h2 ;  
   wire _GEN_31=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_32=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_33=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_35=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_36=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_37=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [151:0] _GEN_38={144'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [31:0] _a_set_wo_ready_T=32'h1<<_GEN_0 ;  
   wire [18:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_39=io_in_d_valid&d_first_1 ;  
   wire _GEN_40=_GEN_39&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_41={14'h0,io_in_d_bits_source} ;  
   wire _GEN_42=_GEN_40&same_cycle_resp&~reset ;  
   wire _GEN_43=_GEN_40&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_44={4'h0,io_in_d_bits_size} ;  
   wire _GEN_45=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_46=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_47=inflight>>_GEN_41 ;  
   wire [151:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_38 ;  
   wire [31:0] _d_clr_wo_ready_T=32'h1<<_GEN_2 ;  
   wire [18:0] _GEN_48=inflight_1>>_GEN_41 ;  
   wire [151:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_38 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~(_GEN_17|_GEN_18&(_GEN_6|_GEN_8|_GEN_9|(&(io_in_a_bits_address[27:26])))))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(_GEN_15&_GEN_17))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_28)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_46[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~reset&~(_GEN_47[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&_GEN_44!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_40 ? _d_clr_wo_ready_T[18:0]:19'h0)|a_set_wo_ready==19'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 2 (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&~(_GEN_48[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&_GEN_44!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/PeripheryBus.scala:58:7)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_49={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_49 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_49 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_49 ;  
   wire [270:0] _GEN_50={263'h0,io_in_d_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_2 ;  
   wire [31:0] _a_set_T=32'h1<<_GEN_0 ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<{264'h0,io_in_d_bits_source,2'h0} ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _d_sizes_clr_T_5=271'hFF<<_GEN_50 ;  
   wire [259:0] _a_sizes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{252'h0,io_in_a_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_2 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hFF<<_GEN_50 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_51=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_52=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=152'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=152'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[18:0]:19'h0))&~(_GEN_51 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_51 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[151:0]:152'h0))&~(_GEN_51 ? _d_sizes_clr_T_5[151:0]:152'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_52 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_52 ? _d_sizes_clr_T_11[151:0]:152'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLAtomicAutomata_1 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [27:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [4:0] auto_out_a_bits_source,
  output [27:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [4:0] auto_out_d_bits_source,
  input auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   wire source_i_ready ;  
   reg [1:0] cam_s_state_0 ;  
   reg [2:0] cam_a_0_bits_opcode ;  
   reg [2:0] cam_a_0_bits_param ;  
   reg [3:0] cam_a_0_bits_size ;  
   reg [4:0] cam_a_0_bits_source ;  
   reg [27:0] cam_a_0_bits_address ;  
   reg [7:0] cam_a_0_bits_mask ;  
   reg [63:0] cam_a_0_bits_data ;  
   reg cam_a_0_bits_corrupt ;  
   reg [3:0] cam_a_0_lut ;  
   reg [63:0] cam_d_data_0 ;  
   reg cam_d_denied_0 ;  
   reg cam_d_corrupt_0 ;  
   wire cam_free_0=cam_s_state_0==2'h0 ;  
   wire winner_0=cam_s_state_0==2'h2 ;  
   wire _a_canArithmetic_T_3=auto_in_a_bits_size<4'h4 ;  
   wire [3:0] _GEN={auto_in_a_bits_address[27],auto_in_a_bits_address[25],auto_in_a_bits_address[16],~(auto_in_a_bits_address[13])} ;  
   wire a_isSupported=auto_in_a_bits_opcode==3'h3 ? _a_canArithmetic_T_3&~(|_GEN):auto_in_a_bits_opcode!=3'h2|_a_canArithmetic_T_3&~(|_GEN) ;  
   wire [3:0] _logic_out_T=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[0],cam_d_data_0[0]} ;  
   wire [3:0] _logic_out_T_2=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[1],cam_d_data_0[1]} ;  
   wire [3:0] _logic_out_T_4=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[2],cam_d_data_0[2]} ;  
   wire [3:0] _logic_out_T_6=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[3],cam_d_data_0[3]} ;  
   wire [3:0] _logic_out_T_8=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[4],cam_d_data_0[4]} ;  
   wire [3:0] _logic_out_T_10=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[5],cam_d_data_0[5]} ;  
   wire [3:0] _logic_out_T_12=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[6],cam_d_data_0[6]} ;  
   wire [3:0] _logic_out_T_14=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[7],cam_d_data_0[7]} ;  
   wire [3:0] _logic_out_T_16=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[8],cam_d_data_0[8]} ;  
   wire [3:0] _logic_out_T_18=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[9],cam_d_data_0[9]} ;  
   wire [3:0] _logic_out_T_20=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[10],cam_d_data_0[10]} ;  
   wire [3:0] _logic_out_T_22=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[11],cam_d_data_0[11]} ;  
   wire [3:0] _logic_out_T_24=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[12],cam_d_data_0[12]} ;  
   wire [3:0] _logic_out_T_26=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[13],cam_d_data_0[13]} ;  
   wire [3:0] _logic_out_T_28=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[14],cam_d_data_0[14]} ;  
   wire [3:0] _logic_out_T_30=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[15],cam_d_data_0[15]} ;  
   wire [3:0] _logic_out_T_32=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[16],cam_d_data_0[16]} ;  
   wire [3:0] _logic_out_T_34=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[17],cam_d_data_0[17]} ;  
   wire [3:0] _logic_out_T_36=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[18],cam_d_data_0[18]} ;  
   wire [3:0] _logic_out_T_38=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[19],cam_d_data_0[19]} ;  
   wire [3:0] _logic_out_T_40=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[20],cam_d_data_0[20]} ;  
   wire [3:0] _logic_out_T_42=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[21],cam_d_data_0[21]} ;  
   wire [3:0] _logic_out_T_44=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[22],cam_d_data_0[22]} ;  
   wire [3:0] _logic_out_T_46=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[23],cam_d_data_0[23]} ;  
   wire [3:0] _logic_out_T_48=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[24],cam_d_data_0[24]} ;  
   wire [3:0] _logic_out_T_50=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[25],cam_d_data_0[25]} ;  
   wire [3:0] _logic_out_T_52=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[26],cam_d_data_0[26]} ;  
   wire [3:0] _logic_out_T_54=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[27],cam_d_data_0[27]} ;  
   wire [3:0] _logic_out_T_56=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[28],cam_d_data_0[28]} ;  
   wire [3:0] _logic_out_T_58=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[29],cam_d_data_0[29]} ;  
   wire [3:0] _logic_out_T_60=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[30],cam_d_data_0[30]} ;  
   wire [3:0] _logic_out_T_62=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[31],cam_d_data_0[31]} ;  
   wire [3:0] _logic_out_T_64=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[32],cam_d_data_0[32]} ;  
   wire [3:0] _logic_out_T_66=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[33],cam_d_data_0[33]} ;  
   wire [3:0] _logic_out_T_68=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[34],cam_d_data_0[34]} ;  
   wire [3:0] _logic_out_T_70=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[35],cam_d_data_0[35]} ;  
   wire [3:0] _logic_out_T_72=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[36],cam_d_data_0[36]} ;  
   wire [3:0] _logic_out_T_74=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[37],cam_d_data_0[37]} ;  
   wire [3:0] _logic_out_T_76=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[38],cam_d_data_0[38]} ;  
   wire [3:0] _logic_out_T_78=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[39],cam_d_data_0[39]} ;  
   wire [3:0] _logic_out_T_80=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[40],cam_d_data_0[40]} ;  
   wire [3:0] _logic_out_T_82=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[41],cam_d_data_0[41]} ;  
   wire [3:0] _logic_out_T_84=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[42],cam_d_data_0[42]} ;  
   wire [3:0] _logic_out_T_86=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[43],cam_d_data_0[43]} ;  
   wire [3:0] _logic_out_T_88=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[44],cam_d_data_0[44]} ;  
   wire [3:0] _logic_out_T_90=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[45],cam_d_data_0[45]} ;  
   wire [3:0] _logic_out_T_92=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[46],cam_d_data_0[46]} ;  
   wire [3:0] _logic_out_T_94=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[47],cam_d_data_0[47]} ;  
   wire [3:0] _logic_out_T_96=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[48],cam_d_data_0[48]} ;  
   wire [3:0] _logic_out_T_98=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[49],cam_d_data_0[49]} ;  
   wire [3:0] _logic_out_T_100=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[50],cam_d_data_0[50]} ;  
   wire [3:0] _logic_out_T_102=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[51],cam_d_data_0[51]} ;  
   wire [3:0] _logic_out_T_104=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[52],cam_d_data_0[52]} ;  
   wire [3:0] _logic_out_T_106=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[53],cam_d_data_0[53]} ;  
   wire [3:0] _logic_out_T_108=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[54],cam_d_data_0[54]} ;  
   wire [3:0] _logic_out_T_110=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[55],cam_d_data_0[55]} ;  
   wire [3:0] _logic_out_T_112=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[56],cam_d_data_0[56]} ;  
   wire [3:0] _logic_out_T_114=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[57],cam_d_data_0[57]} ;  
   wire [3:0] _logic_out_T_116=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[58],cam_d_data_0[58]} ;  
   wire [3:0] _logic_out_T_118=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[59],cam_d_data_0[59]} ;  
   wire [3:0] _logic_out_T_120=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[60],cam_d_data_0[60]} ;  
   wire [3:0] _logic_out_T_122=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[61],cam_d_data_0[61]} ;  
   wire [3:0] _logic_out_T_124=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[62],cam_d_data_0[62]} ;  
   wire [3:0] _logic_out_T_126=cam_a_0_lut>>{2'h0,cam_a_0_bits_data[63],cam_d_data_0[63]} ;  
   wire [6:0] _GEN_0=~(cam_a_0_bits_mask[6:0])|cam_a_0_bits_mask[7:1] ;  
   wire [6:0] _signbit_a_T={cam_a_0_bits_data[55],cam_a_0_bits_data[47],cam_a_0_bits_data[39],cam_a_0_bits_data[31],cam_a_0_bits_data[23],cam_a_0_bits_data[15],cam_a_0_bits_data[7]}&~_GEN_0 ;  
   wire [6:0] _signbit_d_T={cam_d_data_0[55],cam_d_data_0[47],cam_d_data_0[39],cam_d_data_0[31],cam_d_data_0[23],cam_d_data_0[15],cam_d_data_0[7]}&~_GEN_0 ;  
   wire [5:0] _GEN_1=_signbit_a_T[6:1]|_signbit_a_T[5:0] ;  
   wire [3:0] _GEN_2=_GEN_1[5:2]|_GEN_1[3:0] ;  
   wire _signext_a_T_24=_GEN_1[1]|_signbit_a_T[0] ;  
   wire [5:0] _GEN_3=_signbit_d_T[6:1]|_signbit_d_T[5:0] ;  
   wire [3:0] _GEN_4=_GEN_3[5:2]|_GEN_3[3:0] ;  
   wire _signext_d_T_24=_GEN_3[1]|_signbit_d_T[0] ;  
   wire [63:0] wide_mask={{8{cam_a_0_bits_mask[7]}},{8{cam_a_0_bits_mask[6]}},{8{cam_a_0_bits_mask[5]}},{8{cam_a_0_bits_mask[4]}},{8{cam_a_0_bits_mask[3]}},{8{cam_a_0_bits_mask[2]}},{8{cam_a_0_bits_mask[1]}},{8{cam_a_0_bits_mask[0]}}} ;  
   wire [63:0] a_a_ext=cam_a_0_bits_data&wide_mask|{{8{_GEN_2[3]|_signext_a_T_24}},{8{_GEN_2[2]|_GEN_1[0]}},{8{_GEN_2[1]|_signbit_a_T[0]}},{8{_GEN_2[0]}},{8{_signext_a_T_24}},{8{_GEN_1[0]}},{8{_signbit_a_T[0]}},8'h0} ;  
   wire [63:0] a_d_ext=cam_d_data_0&wide_mask|{{8{_GEN_4[3]|_signext_d_T_24}},{8{_GEN_4[2]|_GEN_3[0]}},{8{_GEN_4[1]|_signbit_d_T[0]}},{8{_GEN_4[0]}},{8{_signext_d_T_24}},{8{_GEN_3[0]}},{8{_signbit_d_T[0]}},8'h0} ;  
   wire [63:0] _adder_out_T=a_a_ext+({64{~(cam_a_0_bits_param[2])}}^a_d_ext) ;  
   wire a_allow=~((&cam_s_state_0)|winner_0)&(a_isSupported|cam_free_0) ;  
   wire nodeIn_a_ready=source_i_ready&a_allow ;  
   wire source_i_valid=auto_in_a_valid&a_allow ;  
   wire _source_c_bits_a_mask_T=cam_a_0_bits_size>4'h2 ;  
   wire source_c_bits_a_mask_size=cam_a_0_bits_size[1:0]==2'h2 ;  
   wire source_c_bits_a_mask_acc=_source_c_bits_a_mask_T|source_c_bits_a_mask_size&~(cam_a_0_bits_address[2]) ;  
   wire source_c_bits_a_mask_acc_1=_source_c_bits_a_mask_T|source_c_bits_a_mask_size&cam_a_0_bits_address[2] ;  
   wire source_c_bits_a_mask_size_1=cam_a_0_bits_size[1:0]==2'h1 ;  
   wire source_c_bits_a_mask_eq_2=~(cam_a_0_bits_address[2])&~(cam_a_0_bits_address[1]) ;  
   wire source_c_bits_a_mask_acc_2=source_c_bits_a_mask_acc|source_c_bits_a_mask_size_1&source_c_bits_a_mask_eq_2 ;  
   wire source_c_bits_a_mask_eq_3=~(cam_a_0_bits_address[2])&cam_a_0_bits_address[1] ;  
   wire source_c_bits_a_mask_acc_3=source_c_bits_a_mask_acc|source_c_bits_a_mask_size_1&source_c_bits_a_mask_eq_3 ;  
   wire source_c_bits_a_mask_eq_4=cam_a_0_bits_address[2]&~(cam_a_0_bits_address[1]) ;  
   wire source_c_bits_a_mask_acc_4=source_c_bits_a_mask_acc_1|source_c_bits_a_mask_size_1&source_c_bits_a_mask_eq_4 ;  
   wire source_c_bits_a_mask_eq_5=cam_a_0_bits_address[2]&cam_a_0_bits_address[1] ;  
   wire source_c_bits_a_mask_acc_5=source_c_bits_a_mask_acc_1|source_c_bits_a_mask_size_1&source_c_bits_a_mask_eq_5 ;  
   reg [8:0] beatsLeft ;  
   wire idle=beatsLeft==9'h0 ;  
   wire winner_1=~winner_0&source_i_valid ;  
   wire _nodeOut_a_valid_T=winner_0|source_i_valid ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~winner_0|~winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_nodeOut_a_valid_T|winner_0|winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg state_0 ;  
   reg state_1 ;  
   wire muxState_0=idle ? winner_0:state_0 ;  
   wire muxState_1=idle ? winner_1:state_1 ;  
  assign source_i_ready=auto_out_a_ready&(idle ? ~winner_0:state_1); 
   wire nodeOut_a_valid=idle ? _nodeOut_a_valid_T:state_0&winner_0|state_1&source_i_valid ;  
   reg [3:0] casez_tmp ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_param[1:0])
          2 'b00:
             casez_tmp =4'h6;
          2 'b01:
             casez_tmp =4'hE;
          2 'b10:
             casez_tmp =4'h8;
          default :
             casez_tmp =4'hC;
         endcase 
       end
  
   reg [8:0] d_first_counter ;  
   wire d_first=d_first_counter==9'h0 ;  
   wire d_cam_sel_0=cam_a_0_bits_source==auto_out_d_bits_source&(|cam_s_state_0) ;  
   wire d_ackd=auto_out_d_bits_opcode==3'h1 ;  
   wire d_drop=d_first&d_ackd&d_cam_sel_0 ;  
   wire d_replace=d_first&auto_out_d_bits_opcode==3'h0&d_cam_sel_0 ;  
   wire nodeIn_d_valid=auto_out_d_valid&~d_drop ;  
   wire nodeOut_d_ready=auto_in_d_ready|d_drop ;  
   wire [2:0] nodeIn_d_bits_opcode=d_replace ? 3'h1:auto_out_d_bits_opcode ;  
   wire nodeIn_d_bits_corrupt=d_replace ? cam_d_corrupt_0|auto_out_d_bits_denied:auto_out_d_bits_corrupt ;  
   wire nodeIn_d_bits_denied=d_replace&cam_d_denied_0|auto_out_d_bits_denied ;  
   wire [26:0] _decode_T_1=27'hFFF<<auto_in_a_bits_size ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<auto_out_d_bits_size ;  
   wire _GEN_5=source_i_ready&source_i_valid&~a_isSupported&cam_free_0 ;  
   wire _d_first_T=nodeOut_d_ready&auto_out_d_valid ;  
   wire _GEN_6=_d_first_T&d_first ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              cam_s_state_0 <=2'h0;
              beatsLeft <=9'h0;
              state_0 <=1'h0;
              state_1 <=1'h0;
              d_first_counter <=9'h0;
            end 
          else 
            begin 
              if (_GEN_6&d_cam_sel_0)
                 cam_s_state_0 <={d_ackd,1'h0};
               else 
                 if (auto_out_a_ready&(idle|state_0)&winner_0)
                    cam_s_state_0 <=2'h1;
                  else 
                    if (_GEN_5)
                       cam_s_state_0 <=2'h3;
              if (idle&auto_out_a_ready)
                 beatsLeft <=winner_1&~(auto_in_a_bits_opcode[2]) ? ~(_decode_T_1[11:3]):9'h0;
               else 
                 beatsLeft <=beatsLeft-{8'h0,auto_out_a_ready&nodeOut_a_valid};
              if (idle)
                 begin 
                   state_0 <=winner_0;
                   state_1 <=winner_1;
                 end 
              if (_d_first_T)
                 begin 
                   if (d_first)
                      d_first_counter <=auto_out_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                    else 
                      d_first_counter <=d_first_counter-9'h1;
                 end 
            end 
         if (_GEN_5)
            begin 
              cam_a_0_bits_opcode <=auto_in_a_bits_opcode;
              cam_a_0_bits_param <=auto_in_a_bits_param;
              cam_a_0_bits_size <=auto_in_a_bits_size;
              cam_a_0_bits_source <=auto_in_a_bits_source;
              cam_a_0_bits_address <=auto_in_a_bits_address;
              cam_a_0_bits_mask <=auto_in_a_bits_mask;
              cam_a_0_bits_data <=auto_in_a_bits_data;
              cam_a_0_bits_corrupt <=auto_in_a_bits_corrupt;
              cam_a_0_lut <=casez_tmp;
            end 
         if (_GEN_6&d_cam_sel_0&d_ackd)
            begin 
              cam_d_data_0 <=auto_out_d_bits_data;
              cam_d_denied_0 <=auto_out_d_bits_denied;
              cam_d_corrupt_0 <=auto_out_d_bits_corrupt;
            end 
       end
  
  TLMonitor_11 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(nodeIn_d_bits_opcode),.io_in_d_bits_param(auto_out_d_bits_param),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source),.io_in_d_bits_sink(auto_out_d_bits_sink),.io_in_d_bits_denied(nodeIn_d_bits_denied),.io_in_d_bits_corrupt(nodeIn_d_bits_corrupt)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=nodeIn_d_bits_opcode; 
  assign auto_in_d_bits_param=auto_out_d_bits_param; 
  assign auto_in_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source; 
  assign auto_in_d_bits_sink=auto_out_d_bits_sink; 
  assign auto_in_d_bits_denied=nodeIn_d_bits_denied; 
  assign auto_in_d_bits_data=d_replace ? cam_d_data_0:auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt=nodeIn_d_bits_corrupt; 
  assign auto_out_a_valid=nodeOut_a_valid; 
  assign auto_out_a_bits_opcode=muxState_1 ? (a_isSupported ? auto_in_a_bits_opcode:3'h4):3'h0; 
  assign auto_out_a_bits_param=muxState_1&a_isSupported ? auto_in_a_bits_param:3'h0; 
  assign auto_out_a_bits_size=(muxState_0 ? cam_a_0_bits_size:4'h0)|(muxState_1 ? auto_in_a_bits_size:4'h0); 
  assign auto_out_a_bits_source=(muxState_0 ? cam_a_0_bits_source:5'h0)|(muxState_1 ? auto_in_a_bits_source:5'h0); 
  assign auto_out_a_bits_address=(muxState_0 ? cam_a_0_bits_address:28'h0)|(muxState_1 ? auto_in_a_bits_address:28'h0); 
  assign auto_out_a_bits_mask=(muxState_0 ? {source_c_bits_a_mask_acc_5|source_c_bits_a_mask_eq_5&cam_a_0_bits_address[0],source_c_bits_a_mask_acc_5|source_c_bits_a_mask_eq_5&~(cam_a_0_bits_address[0]),source_c_bits_a_mask_acc_4|source_c_bits_a_mask_eq_4&cam_a_0_bits_address[0],source_c_bits_a_mask_acc_4|source_c_bits_a_mask_eq_4&~(cam_a_0_bits_address[0]),source_c_bits_a_mask_acc_3|source_c_bits_a_mask_eq_3&cam_a_0_bits_address[0],source_c_bits_a_mask_acc_3|source_c_bits_a_mask_eq_3&~(cam_a_0_bits_address[0]),source_c_bits_a_mask_acc_2|source_c_bits_a_mask_eq_2&cam_a_0_bits_address[0],source_c_bits_a_mask_acc_2|source_c_bits_a_mask_eq_2&~(cam_a_0_bits_address[0])}:8'h0)|(muxState_1 ? auto_in_a_bits_mask:8'h0); 
  assign auto_out_a_bits_data=(muxState_0 ? (cam_a_0_bits_opcode[0] ? {_logic_out_T_126[0],_logic_out_T_124[0],_logic_out_T_122[0],_logic_out_T_120[0],_logic_out_T_118[0],_logic_out_T_116[0],_logic_out_T_114[0],_logic_out_T_112[0],_logic_out_T_110[0],_logic_out_T_108[0],_logic_out_T_106[0],_logic_out_T_104[0],_logic_out_T_102[0],_logic_out_T_100[0],_logic_out_T_98[0],_logic_out_T_96[0],_logic_out_T_94[0],_logic_out_T_92[0],_logic_out_T_90[0],_logic_out_T_88[0],_logic_out_T_86[0],_logic_out_T_84[0],_logic_out_T_82[0],_logic_out_T_80[0],_logic_out_T_78[0],_logic_out_T_76[0],_logic_out_T_74[0],_logic_out_T_72[0],_logic_out_T_70[0],_logic_out_T_68[0],_logic_out_T_66[0],_logic_out_T_64[0],_logic_out_T_62[0],_logic_out_T_60[0],_logic_out_T_58[0],_logic_out_T_56[0],_logic_out_T_54[0],_logic_out_T_52[0],_logic_out_T_50[0],_logic_out_T_48[0],_logic_out_T_46[0],_logic_out_T_44[0],_logic_out_T_42[0],_logic_out_T_40[0],_logic_out_T_38[0],_logic_out_T_36[0],_logic_out_T_34[0],_logic_out_T_32[0],_logic_out_T_30[0],_logic_out_T_28[0],_logic_out_T_26[0],_logic_out_T_24[0],_logic_out_T_22[0],_logic_out_T_20[0],_logic_out_T_18[0],_logic_out_T_16[0],_logic_out_T_14[0],_logic_out_T_12[0],_logic_out_T_10[0],_logic_out_T_8[0],_logic_out_T_6[0],_logic_out_T_4[0],_logic_out_T_2[0],_logic_out_T[0]}:cam_a_0_bits_param[2] ? _adder_out_T:cam_a_0_bits_param[0]==(a_a_ext[63]==a_d_ext[63] ? ~(_adder_out_T[63]):cam_a_0_bits_param[1]==a_a_ext[63]) ? cam_a_0_bits_data:cam_d_data_0):64'h0)|(muxState_1 ? auto_in_a_bits_data:64'h0); 
  assign auto_out_a_bits_corrupt=muxState_0&(cam_a_0_bits_corrupt|cam_d_corrupt_0)|muxState_1&auto_in_a_bits_corrupt; 
  assign auto_out_d_ready=nodeOut_d_ready; 
endmodule
 
module TLMonitor_12 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [13:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [3:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [4:0] source ;  
   reg [13:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [3:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [151:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>{69'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _GEN_0={27'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [31:0] _GEN_2={27'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [151:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=_GEN_4&(&(io_in_a_bits_address[13:12])) ;  
   wire _GEN_7=_source_ok_T_12&io_in_a_bits_size==4'h6&_GEN_6 ;  
   wire _GEN_8=io_in_a_bits_param>3'h2 ;  
   wire _GEN_9=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_10=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_11=_GEN_4&(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14) ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_13=io_in_a_bits_mask!=mask ;  
   wire _GEN_14=_GEN_11&_GEN_6 ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_17=_GEN_11&io_in_a_bits_size<4'h4&(&(io_in_a_bits_address[13:12])) ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_19=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_20=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_21=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_22=io_in_d_bits_size<4'h3 ;  
   wire _GEN_23=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_24=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_25=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_26=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_27=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_28=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_29=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [151:0] _GEN_30={144'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [31:0] _a_set_wo_ready_T=32'h1<<_GEN_0 ;  
   wire [18:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_31=io_in_d_valid&d_first_1 ;  
   wire _GEN_32=_GEN_31&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_33={14'h0,io_in_d_bits_source} ;  
   wire _GEN_34=_GEN_32&same_cycle_resp&~reset ;  
   wire _GEN_35=_GEN_32&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_36={4'h0,io_in_d_bits_size} ;  
   wire _GEN_37=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_38=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_39=inflight>>_GEN_33 ;  
   wire [151:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_30 ;  
   wire [31:0] _d_clr_wo_ready_T=32'h1<<_GEN_2 ;  
   wire [18:0] _GEN_40=inflight_1>>_GEN_33 ;  
   wire [151:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_30 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_38[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~reset&~(_GEN_39[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&_GEN_36!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_32 ? _d_clr_wo_ready_T[18:0]:19'h0)|a_set_wo_ready==19'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~(_GEN_40[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&_GEN_36!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:43:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_41={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_41 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_41 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_41 ;  
   wire [270:0] _GEN_42={263'h0,io_in_d_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_2 ;  
   wire [31:0] _a_set_T=32'h1<<_GEN_0 ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<{264'h0,io_in_d_bits_source,2'h0} ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _d_sizes_clr_T_5=271'hFF<<_GEN_42 ;  
   wire [259:0] _a_sizes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{252'h0,io_in_a_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_2 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hFF<<_GEN_42 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_43=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_44=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=152'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=152'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[18:0]:19'h0))&~(_GEN_43 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_43 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[151:0]:152'h0))&~(_GEN_43 ? _d_sizes_clr_T_5[151:0]:152'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_44 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_44 ? _d_sizes_clr_T_11[151:0]:152'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module Queue_37 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [3:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source) ; 
   reg [4:0] ram_source ;  
   reg [3:0] ram_size ;  
   reg [2:0] ram_opcode ;  
   reg full ;  
   wire do_enq=~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_source <=io_enq_bits_source;
              ram_size <=io_enq_bits_size;
              ram_opcode <=io_enq_bits_opcode;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(io_deq_ready&full)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=full; 
  assign io_deq_bits_opcode=ram_opcode; 
  assign io_deq_bits_size=ram_size; 
  assign io_deq_bits_source=ram_source; 
endmodule
 
module TLError (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [13:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [3:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output auto_in_d_bits_corrupt) ; 
   reg [2:0] casez_tmp ;  
   wire _a_q_io_enq_ready ;  
   wire _a_q_io_deq_valid ;  
   wire [2:0] _a_q_io_deq_bits_opcode ;  
   wire [3:0] _a_q_io_deq_bits_size ;  
   wire [4:0] _a_q_io_deq_bits_source ;  
   wire [26:0] _GEN={23'h0,_a_q_io_deq_bits_size} ;  
   wire [26:0] _a_last_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [8:0] a_last_beats1=_a_q_io_deq_bits_opcode[2] ? 9'h0:~(_a_last_beats1_decode_T_1[11:3]) ;  
   reg [8:0] a_last_counter ;  
   wire a_last=a_last_counter==9'h1|a_last_beats1==9'h0 ;  
   wire [26:0] _beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [8:0] beats1=casez_tmp[0] ? ~(_beats1_decode_T_1[11:3]):9'h0 ;  
   reg [8:0] counter ;  
   wire a_q_io_deq_ready=auto_in_d_ready&(counter==9'h1|beats1==9'h0)|~a_last ;  
   wire da_valid=_a_q_io_deq_valid&a_last ;  
  always @(*)
       begin 
         casez (_a_q_io_deq_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_last_counter <=9'h0;
              counter <=9'h0;
            end 
          else 
            begin 
              if (a_q_io_deq_ready&_a_q_io_deq_valid)
                 begin 
                   if (a_last_counter==9'h0)
                      a_last_counter <=a_last_beats1;
                    else 
                      a_last_counter <=a_last_counter-9'h1;
                 end 
              if (auto_in_d_ready&da_valid)
                 begin 
                   if (counter==9'h0)
                      counter <=beats1;
                    else 
                      counter <=counter-9'h1;
                 end 
            end 
       end
  
  TLMonitor_12 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_a_q_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(da_valid),.io_in_d_bits_opcode(casez_tmp),.io_in_d_bits_size(_a_q_io_deq_bits_size),.io_in_d_bits_source(_a_q_io_deq_bits_source),.io_in_d_bits_corrupt(casez_tmp[0])); 
  Queue_37 a_q(.clock(clock),.reset(reset),.io_enq_ready(_a_q_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_deq_ready(a_q_io_deq_ready),.io_deq_valid(_a_q_io_deq_valid),.io_deq_bits_opcode(_a_q_io_deq_bits_opcode),.io_deq_bits_size(_a_q_io_deq_bits_size),.io_deq_bits_source(_a_q_io_deq_bits_source)); 
  assign auto_in_a_ready=_a_q_io_enq_ready; 
  assign auto_in_d_valid=da_valid; 
  assign auto_in_d_bits_opcode=casez_tmp; 
  assign auto_in_d_bits_size=_a_q_io_deq_bits_size; 
  assign auto_in_d_bits_source=_a_q_io_deq_bits_source; 
  assign auto_in_d_bits_corrupt=casez_tmp[0]; 
endmodule
 
module TLMonitor_13 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [13:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [4:0] source ;  
   reg [13:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg sink ;  
   reg denied ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [151:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>{69'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _GEN_0={27'h0,io_in_a_bits_source} ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [31:0] _GEN_2={27'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [151:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_3=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_bits_size<4'hD ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=_GEN_4&(&(io_in_a_bits_address[13:12])) ;  
   wire _GEN_7=_source_ok_T_12&io_in_a_bits_size==4'h6&_GEN_6 ;  
   wire _GEN_8=io_in_a_bits_param>3'h2 ;  
   wire _GEN_9=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_10=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_11=_GEN_4&(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14) ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_13=io_in_a_bits_mask!=mask ;  
   wire _GEN_14=_GEN_11&_GEN_6 ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_17=_GEN_11&io_in_a_bits_size<4'h4&(&(io_in_a_bits_address[13:12])) ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_19=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_20=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_21=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_22=io_in_d_bits_size<4'h3 ;  
   wire _GEN_23=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_24=io_in_d_bits_param==2'h2 ;  
   wire _GEN_25=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_26=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_27=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_28=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_29=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_30=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_31=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire [151:0] _GEN_32={144'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [31:0] _a_set_wo_ready_T=32'h1<<_GEN_0 ;  
   wire [18:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_33=io_in_d_valid&d_first_1 ;  
   wire _GEN_34=_GEN_33&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_35={14'h0,io_in_d_bits_source} ;  
   wire _GEN_36=_GEN_34&same_cycle_resp&~reset ;  
   wire _GEN_37=_GEN_34&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_38={4'h0,io_in_d_bits_size} ;  
   wire _GEN_39=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_40=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_41=inflight>>_GEN_35 ;  
   wire [151:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_32 ;  
   wire [31:0] _d_clr_wo_ready_T=32'h1<<_GEN_2 ;  
   wire [18:0] _GEN_42=inflight_1>>_GEN_35 ;  
   wire [151:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_32 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_40[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~reset&~(_GEN_41[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&_GEN_38!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_34 ? _d_clr_wo_ready_T[18:0]:19'h0)|a_set_wo_ready==19'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&~(_GEN_42[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&_GEN_38!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CanHaveBuiltInDevices.scala:44:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_43={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_43 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_43 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_43 ;  
   wire [270:0] _GEN_44={263'h0,io_in_d_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_2 ;  
   wire [31:0] _a_set_T=32'h1<<_GEN_0 ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<{264'h0,io_in_d_bits_source,2'h0} ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _d_sizes_clr_T_5=271'hFF<<_GEN_44 ;  
   wire [259:0] _a_sizes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:5'h0}<<{252'h0,io_in_a_bits_source,3'h0} ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_2 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hFF<<_GEN_44 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_45=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_46=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=152'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=152'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[18:0]:19'h0))&~(_GEN_45 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_45 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[151:0]:152'h0))&~(_GEN_45 ? _d_sizes_clr_T_5[151:0]:152'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_46 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_46 ? _d_sizes_clr_T_11[151:0]:152'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module ram_address_2x14 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [13:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [13:0] W0_data) ; 
   reg [13:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:14'bx; 
endmodule
 
module Queue_38 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input [13:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source,
  output [13:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x3 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_source_2x5 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_address_2x14 ram_address_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_address),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_address)); 
  ram_2x8 ram_mask_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_mask),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_mask)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_corrupt)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module TLBuffer_5 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [13:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [4:0] auto_out_a_bits_source,
  output [13:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [3:0] auto_out_d_bits_size,
  input [4:0] auto_out_d_bits_source,
  input auto_out_d_bits_corrupt) ; 
   wire _nodeIn_d_q_io_deq_valid ;  
   wire [2:0] _nodeIn_d_q_io_deq_bits_opcode ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_param ;  
   wire [3:0] _nodeIn_d_q_io_deq_bits_size ;  
   wire [4:0] _nodeIn_d_q_io_deq_bits_source ;  
   wire _nodeIn_d_q_io_deq_bits_sink ;  
   wire _nodeIn_d_q_io_deq_bits_denied ;  
   wire _nodeIn_d_q_io_deq_bits_corrupt ;  
   wire _nodeOut_a_q_io_enq_ready ;  
  TLMonitor_13 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_nodeOut_a_q_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(_nodeIn_d_q_io_deq_valid),.io_in_d_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_in_d_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_in_d_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_in_d_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_in_d_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_in_d_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_in_d_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  Queue_38 nodeOut_a_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_a_q_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_corrupt(auto_in_a_bits_corrupt),.io_deq_ready(auto_out_a_ready),.io_deq_valid(auto_out_a_valid),.io_deq_bits_opcode(auto_out_a_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(auto_out_a_bits_size),.io_deq_bits_source(auto_out_a_bits_source),.io_deq_bits_address(auto_out_a_bits_address),.io_deq_bits_mask(auto_out_a_bits_mask),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  Queue_36 nodeIn_d_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_d_ready),.io_enq_valid(auto_out_d_valid),.io_enq_bits_opcode(auto_out_d_bits_opcode),.io_enq_bits_param(2'h0),.io_enq_bits_size(auto_out_d_bits_size),.io_enq_bits_source(auto_out_d_bits_source),.io_enq_bits_sink(1'h0),.io_enq_bits_denied(1'h1),.io_enq_bits_data(64'h0),.io_enq_bits_corrupt(auto_out_d_bits_corrupt),.io_deq_ready(auto_in_d_ready),.io_deq_valid(_nodeIn_d_q_io_deq_valid),.io_deq_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_deq_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_deq_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_deq_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_deq_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_deq_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_deq_bits_data(auto_in_d_bits_data),.io_deq_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  assign auto_in_a_ready=_nodeOut_a_q_io_enq_ready; 
  assign auto_in_d_valid=_nodeIn_d_q_io_deq_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_q_io_deq_bits_opcode; 
  assign auto_in_d_bits_param=_nodeIn_d_q_io_deq_bits_param; 
  assign auto_in_d_bits_size=_nodeIn_d_q_io_deq_bits_size; 
  assign auto_in_d_bits_source=_nodeIn_d_q_io_deq_bits_source; 
  assign auto_in_d_bits_sink=_nodeIn_d_q_io_deq_bits_sink; 
  assign auto_in_d_bits_denied=_nodeIn_d_q_io_deq_bits_denied; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_q_io_deq_bits_corrupt; 
endmodule
 
module ErrorDeviceWrapper (
  input clock,
  input reset,
  output auto_buffer_in_a_ready,
  input auto_buffer_in_a_valid,
  input [2:0] auto_buffer_in_a_bits_opcode,
  input [2:0] auto_buffer_in_a_bits_param,
  input [3:0] auto_buffer_in_a_bits_size,
  input [4:0] auto_buffer_in_a_bits_source,
  input [13:0] auto_buffer_in_a_bits_address,
  input [7:0] auto_buffer_in_a_bits_mask,
  input auto_buffer_in_a_bits_corrupt,
  input auto_buffer_in_d_ready,
  output auto_buffer_in_d_valid,
  output [2:0] auto_buffer_in_d_bits_opcode,
  output [1:0] auto_buffer_in_d_bits_param,
  output [3:0] auto_buffer_in_d_bits_size,
  output [4:0] auto_buffer_in_d_bits_source,
  output auto_buffer_in_d_bits_sink,
  output auto_buffer_in_d_bits_denied,
  output [63:0] auto_buffer_in_d_bits_data,
  output auto_buffer_in_d_bits_corrupt) ; 
   wire _buffer_auto_out_a_valid ;  
   wire [2:0] _buffer_auto_out_a_bits_opcode ;  
   wire [2:0] _buffer_auto_out_a_bits_param ;  
   wire [3:0] _buffer_auto_out_a_bits_size ;  
   wire [4:0] _buffer_auto_out_a_bits_source ;  
   wire [13:0] _buffer_auto_out_a_bits_address ;  
   wire [7:0] _buffer_auto_out_a_bits_mask ;  
   wire _buffer_auto_out_a_bits_corrupt ;  
   wire _buffer_auto_out_d_ready ;  
   wire _error_auto_in_a_ready ;  
   wire _error_auto_in_d_valid ;  
   wire [2:0] _error_auto_in_d_bits_opcode ;  
   wire [3:0] _error_auto_in_d_bits_size ;  
   wire [4:0] _error_auto_in_d_bits_source ;  
   wire _error_auto_in_d_bits_corrupt ;  
  TLError error(.clock(clock),.reset(reset),.auto_in_a_ready(_error_auto_in_a_ready),.auto_in_a_valid(_buffer_auto_out_a_valid),.auto_in_a_bits_opcode(_buffer_auto_out_a_bits_opcode),.auto_in_a_bits_param(_buffer_auto_out_a_bits_param),.auto_in_a_bits_size(_buffer_auto_out_a_bits_size),.auto_in_a_bits_source(_buffer_auto_out_a_bits_source),.auto_in_a_bits_address(_buffer_auto_out_a_bits_address),.auto_in_a_bits_mask(_buffer_auto_out_a_bits_mask),.auto_in_a_bits_corrupt(_buffer_auto_out_a_bits_corrupt),.auto_in_d_ready(_buffer_auto_out_d_ready),.auto_in_d_valid(_error_auto_in_d_valid),.auto_in_d_bits_opcode(_error_auto_in_d_bits_opcode),.auto_in_d_bits_size(_error_auto_in_d_bits_size),.auto_in_d_bits_source(_error_auto_in_d_bits_source),.auto_in_d_bits_corrupt(_error_auto_in_d_bits_corrupt)); 
  TLBuffer_5 buffer(.clock(clock),.reset(reset),.auto_in_a_ready(auto_buffer_in_a_ready),.auto_in_a_valid(auto_buffer_in_a_valid),.auto_in_a_bits_opcode(auto_buffer_in_a_bits_opcode),.auto_in_a_bits_param(auto_buffer_in_a_bits_param),.auto_in_a_bits_size(auto_buffer_in_a_bits_size),.auto_in_a_bits_source(auto_buffer_in_a_bits_source),.auto_in_a_bits_address(auto_buffer_in_a_bits_address),.auto_in_a_bits_mask(auto_buffer_in_a_bits_mask),.auto_in_a_bits_corrupt(auto_buffer_in_a_bits_corrupt),.auto_in_d_ready(auto_buffer_in_d_ready),.auto_in_d_valid(auto_buffer_in_d_valid),.auto_in_d_bits_opcode(auto_buffer_in_d_bits_opcode),.auto_in_d_bits_param(auto_buffer_in_d_bits_param),.auto_in_d_bits_size(auto_buffer_in_d_bits_size),.auto_in_d_bits_source(auto_buffer_in_d_bits_source),.auto_in_d_bits_sink(auto_buffer_in_d_bits_sink),.auto_in_d_bits_denied(auto_buffer_in_d_bits_denied),.auto_in_d_bits_data(auto_buffer_in_d_bits_data),.auto_in_d_bits_corrupt(auto_buffer_in_d_bits_corrupt),.auto_out_a_ready(_error_auto_in_a_ready),.auto_out_a_valid(_buffer_auto_out_a_valid),.auto_out_a_bits_opcode(_buffer_auto_out_a_bits_opcode),.auto_out_a_bits_param(_buffer_auto_out_a_bits_param),.auto_out_a_bits_size(_buffer_auto_out_a_bits_size),.auto_out_a_bits_source(_buffer_auto_out_a_bits_source),.auto_out_a_bits_address(_buffer_auto_out_a_bits_address),.auto_out_a_bits_mask(_buffer_auto_out_a_bits_mask),.auto_out_a_bits_corrupt(_buffer_auto_out_a_bits_corrupt),.auto_out_d_ready(_buffer_auto_out_d_ready),.auto_out_d_valid(_error_auto_in_d_valid),.auto_out_d_bits_opcode(_error_auto_in_d_bits_opcode),.auto_out_d_bits_size(_error_auto_in_d_bits_size),.auto_out_d_bits_source(_error_auto_in_d_bits_source),.auto_out_d_bits_corrupt(_error_auto_in_d_bits_corrupt)); 
endmodule
 
module TLMonitor_14 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [27:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [2:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [27:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [2:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [75:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [75:0] _GEN_0={69'h0,io_in_d_bits_source,2'h0} ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_0 ;  
   wire [31:0] _GEN_1={27'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [31:0] _GEN_3={27'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [75:0] inflight_sizes_1 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_4=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=_source_ok_T_12&io_in_a_bits_size==3'h6&(&(io_in_a_bits_address[27:26])) ;  
   wire _GEN_7=io_in_a_bits_param>3'h2 ;  
   wire _GEN_8=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_9=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_10=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_12=io_in_a_bits_size!=3'h7&(&(io_in_a_bits_address[27:26])) ;  
   wire _GEN_13=io_in_a_bits_mask!=mask ;  
   wire _GEN_14=_GEN_10&_GEN_12 ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_17=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_19=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_20=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_21=io_in_d_bits_size<3'h3 ;  
   wire _GEN_22=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_23=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_24=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_25=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [31:0] _a_set_wo_ready_T=32'h1<<_GEN_1 ;  
   wire [18:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_26=io_in_d_valid&d_first_1 ;  
   wire _GEN_27=_GEN_26&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_28={14'h0,io_in_d_bits_source} ;  
   wire _GEN_29=_GEN_27&same_cycle_resp&~reset ;  
   wire _GEN_30=_GEN_27&~same_cycle_resp&~reset ;  
   wire _GEN_31=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_32=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_33=inflight>>_GEN_28 ;  
   wire [75:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_0 ;  
   wire [31:0] _d_clr_wo_ready_T=32'h1<<_GEN_3 ;  
   wire [18:0] _GEN_34=inflight_1>>_GEN_28 ;  
   wire [75:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_0 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_32[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~reset&~(_GEN_33[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_27 ? _d_clr_wo_ready_T[18:0]:19'h0)|a_set_wo_ready==19'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&~(_GEN_34[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_31&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/Plic.scala:364:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_35={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_35 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_35 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_35 ;  
   wire [258:0] _GEN_36={252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _GEN_37={264'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_3 ;  
   wire [31:0] _a_set_T=32'h1<<_GEN_1 ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<_GEN_37 ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_36 ;  
   wire [270:0] _d_sizes_clr_T_5=271'hF<<_GEN_37 ;  
   wire [258:0] _a_sizes_set_T_1={255'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_36 ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_3 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hF<<_GEN_37 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_38=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_39=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=76'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=76'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_2 ? _a_set_T[18:0]:19'h0))&~(_GEN_38 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_38 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[75:0]:76'h0))&~(_GEN_38 ? _d_sizes_clr_T_5[75:0]:76'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_39 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_39 ? _d_sizes_clr_T_11[75:0]:76'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module Repeater (
  input clock,
  input reset,
  input io_repeat,
  output io_full,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [2:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input [27:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [2:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source,
  output [27:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output io_deq_bits_corrupt) ; 
   reg full ;  
   reg [2:0] saved_opcode ;  
   reg [2:0] saved_param ;  
   reg [2:0] saved_size ;  
   reg [4:0] saved_source ;  
   reg [27:0] saved_address ;  
   reg [7:0] saved_mask ;  
   reg saved_corrupt ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire io_enq_ready_0=io_deq_ready&~full ;  
   wire _GEN=io_enq_ready_0&io_enq_valid&io_repeat ;  
  always @( posedge clock)
       begin 
         if (reset)
            full <=1'h0;
          else 
            full <=~(io_deq_ready&io_deq_valid_0&~io_repeat)&(_GEN|full);
         if (_GEN)
            begin 
              saved_opcode <=io_enq_bits_opcode;
              saved_param <=io_enq_bits_param;
              saved_size <=io_enq_bits_size;
              saved_source <=io_enq_bits_source;
              saved_address <=io_enq_bits_address;
              saved_mask <=io_enq_bits_mask;
              saved_corrupt <=io_enq_bits_corrupt;
            end 
       end
  
  assign io_full=full; 
  assign io_enq_ready=io_enq_ready_0; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_opcode=full ? saved_opcode:io_enq_bits_opcode; 
  assign io_deq_bits_param=full ? saved_param:io_enq_bits_param; 
  assign io_deq_bits_size=full ? saved_size:io_enq_bits_size; 
  assign io_deq_bits_source=full ? saved_source:io_enq_bits_source; 
  assign io_deq_bits_address=full ? saved_address:io_enq_bits_address; 
  assign io_deq_bits_mask=full ? saved_mask:io_enq_bits_mask; 
  assign io_deq_bits_corrupt=full ? saved_corrupt:io_enq_bits_corrupt; 
endmodule
 
module TLFragmenter (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [27:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [2:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [1:0] auto_out_a_bits_size,
  output [8:0] auto_out_a_bits_source,
  output [27:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_size,
  input [8:0] auto_out_d_bits_source,
  input [63:0] auto_out_d_bits_data) ; 
   wire _repeater_io_full ;  
   wire _repeater_io_enq_ready ;  
   wire _repeater_io_deq_valid ;  
   wire [2:0] _repeater_io_deq_bits_opcode ;  
   wire [2:0] _repeater_io_deq_bits_size ;  
   wire [4:0] _repeater_io_deq_bits_source ;  
   wire [27:0] _repeater_io_deq_bits_address ;  
   wire [7:0] _repeater_io_deq_bits_mask ;  
   reg [2:0] acknum ;  
   reg [2:0] dOrig ;  
   reg dToggle ;  
   wire dFirst=acknum==3'h0 ;  
   wire [5:0] _dsizeOH1_T_1=6'h7<<auto_out_d_bits_size ;  
   wire [2:0] _GEN=~(auto_out_d_bits_source[2:0]) ;  
   wire [2:0] dFirst_size_hi=auto_out_d_bits_source[2:0]&{1'h1,_GEN[2:1]} ;  
   wire [2:0] _dFirst_size_T_8={1'h0,dFirst_size_hi[2:1]}|~(_dsizeOH1_T_1[2:0])&{_GEN[0],_dsizeOH1_T_1[2:1]} ;  
   wire [2:0] dFirst_size={|dFirst_size_hi,|(_dFirst_size_T_8[2:1]),_dFirst_size_T_8[2]|_dFirst_size_T_8[0]} ;  
   wire drop=~(auto_out_d_bits_opcode[0])&(|(auto_out_d_bits_source[2:0])) ;  
   wire nodeOut_d_ready=auto_in_d_ready|drop ;  
   wire nodeIn_d_valid=auto_out_d_valid&~drop ;  
   wire [2:0] nodeIn_d_bits_size=dFirst ? dFirst_size:dOrig ;  
   wire [12:0] _aOrigOH1_T_1=13'h3F<<_repeater_io_deq_bits_size ;  
   reg [2:0] gennum ;  
   wire aFirst=gennum==3'h0 ;  
   wire [2:0] _old_gennum1_T_1=gennum-3'h1 ;  
   wire [2:0] aFragnum=aFirst ? ~(_aOrigOH1_T_1[5:3]):_old_gennum1_T_1 ;  
   reg aToggle_r ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~_repeater_io_full|_repeater_io_deq_bits_opcode[2]))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:311 assert (!repeater.io.full || !aHasData)\n");
              if (1)$display("");
            end 
         if (~reset&~(~_repeater_io_full|(&_repeater_io_deq_bits_mask)))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:314 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
              if (1)$display("");
            end 
       end
  
   wire _GEN_0=nodeOut_d_ready&auto_out_d_valid ;  
   wire _GEN_1=_GEN_0&dFirst ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              acknum <=3'h0;
              dToggle <=1'h0;
              gennum <=3'h0;
            end 
          else 
            begin 
              if (_GEN_0)
                 begin 
                   if (dFirst)
                      acknum <=auto_out_d_bits_source[2:0];
                    else 
                      acknum <=acknum-{2'h0,auto_out_d_bits_opcode[0]|(&auto_out_d_bits_size)};
                 end 
              if (_GEN_1)
                 dToggle <=auto_out_d_bits_source[3];
              if (auto_out_a_ready&_repeater_io_deq_valid)
                 begin 
                   if (aFirst)
                      gennum <=~(_aOrigOH1_T_1[5:3]);
                    else 
                      gennum <=_old_gennum1_T_1;
                 end 
            end 
         if (_GEN_1)
            dOrig <=dFirst_size;
         if (aFirst)
            aToggle_r <=dToggle;
       end
  
  TLMonitor_14 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_repeater_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_size(nodeIn_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source[8:4])); 
  Repeater repeater(.clock(clock),.reset(reset),.io_repeat(_repeater_io_deq_bits_opcode[2]&(|aFragnum)),.io_full(_repeater_io_full),.io_enq_ready(_repeater_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_corrupt(auto_in_a_bits_corrupt),.io_deq_ready(auto_out_a_ready),.io_deq_valid(_repeater_io_deq_valid),.io_deq_bits_opcode(_repeater_io_deq_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(_repeater_io_deq_bits_size),.io_deq_bits_source(_repeater_io_deq_bits_source),.io_deq_bits_address(_repeater_io_deq_bits_address),.io_deq_bits_mask(_repeater_io_deq_bits_mask),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  assign auto_in_a_ready=_repeater_io_enq_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size=nodeIn_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source[8:4]; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_out_a_valid=_repeater_io_deq_valid; 
  assign auto_out_a_bits_opcode=_repeater_io_deq_bits_opcode; 
  assign auto_out_a_bits_size=_repeater_io_deq_bits_size[2] ? 2'h3:_repeater_io_deq_bits_size[1:0]; 
  assign auto_out_a_bits_source={_repeater_io_deq_bits_source,~(aFirst ? dToggle:aToggle_r),aFragnum}; 
  assign auto_out_a_bits_address={_repeater_io_deq_bits_address[27:6],_repeater_io_deq_bits_address[5:0]|{~(aFragnum|_aOrigOH1_T_1[5:3]),3'h0}}; 
  assign auto_out_a_bits_mask=_repeater_io_full ? 8'hFF:auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_d_ready=nodeOut_d_ready; 
endmodule
 
module TLInterconnectCoupler_7 (
  input clock,
  input reset,
  input auto_fragmenter_out_a_ready,
  output auto_fragmenter_out_a_valid,
  output [2:0] auto_fragmenter_out_a_bits_opcode,
  output [2:0] auto_fragmenter_out_a_bits_param,
  output [1:0] auto_fragmenter_out_a_bits_size,
  output [8:0] auto_fragmenter_out_a_bits_source,
  output [27:0] auto_fragmenter_out_a_bits_address,
  output [7:0] auto_fragmenter_out_a_bits_mask,
  output [63:0] auto_fragmenter_out_a_bits_data,
  output auto_fragmenter_out_a_bits_corrupt,
  output auto_fragmenter_out_d_ready,
  input auto_fragmenter_out_d_valid,
  input [2:0] auto_fragmenter_out_d_bits_opcode,
  input [1:0] auto_fragmenter_out_d_bits_size,
  input [8:0] auto_fragmenter_out_d_bits_source,
  input [63:0] auto_fragmenter_out_d_bits_data,
  output auto_tl_in_a_ready,
  input auto_tl_in_a_valid,
  input [2:0] auto_tl_in_a_bits_opcode,
  input [2:0] auto_tl_in_a_bits_param,
  input [2:0] auto_tl_in_a_bits_size,
  input [4:0] auto_tl_in_a_bits_source,
  input [27:0] auto_tl_in_a_bits_address,
  input [7:0] auto_tl_in_a_bits_mask,
  input [63:0] auto_tl_in_a_bits_data,
  input auto_tl_in_a_bits_corrupt,
  input auto_tl_in_d_ready,
  output auto_tl_in_d_valid,
  output [2:0] auto_tl_in_d_bits_opcode,
  output [2:0] auto_tl_in_d_bits_size,
  output [4:0] auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data) ; 
  TLFragmenter fragmenter(.clock(clock),.reset(reset),.auto_in_a_ready(auto_tl_in_a_ready),.auto_in_a_valid(auto_tl_in_a_valid),.auto_in_a_bits_opcode(auto_tl_in_a_bits_opcode),.auto_in_a_bits_param(auto_tl_in_a_bits_param),.auto_in_a_bits_size(auto_tl_in_a_bits_size),.auto_in_a_bits_source(auto_tl_in_a_bits_source),.auto_in_a_bits_address(auto_tl_in_a_bits_address),.auto_in_a_bits_mask(auto_tl_in_a_bits_mask),.auto_in_a_bits_data(auto_tl_in_a_bits_data),.auto_in_a_bits_corrupt(auto_tl_in_a_bits_corrupt),.auto_in_d_ready(auto_tl_in_d_ready),.auto_in_d_valid(auto_tl_in_d_valid),.auto_in_d_bits_opcode(auto_tl_in_d_bits_opcode),.auto_in_d_bits_size(auto_tl_in_d_bits_size),.auto_in_d_bits_source(auto_tl_in_d_bits_source),.auto_in_d_bits_data(auto_tl_in_d_bits_data),.auto_out_a_ready(auto_fragmenter_out_a_ready),.auto_out_a_valid(auto_fragmenter_out_a_valid),.auto_out_a_bits_opcode(auto_fragmenter_out_a_bits_opcode),.auto_out_a_bits_param(auto_fragmenter_out_a_bits_param),.auto_out_a_bits_size(auto_fragmenter_out_a_bits_size),.auto_out_a_bits_source(auto_fragmenter_out_a_bits_source),.auto_out_a_bits_address(auto_fragmenter_out_a_bits_address),.auto_out_a_bits_mask(auto_fragmenter_out_a_bits_mask),.auto_out_a_bits_data(auto_fragmenter_out_a_bits_data),.auto_out_a_bits_corrupt(auto_fragmenter_out_a_bits_corrupt),.auto_out_d_ready(auto_fragmenter_out_d_ready),.auto_out_d_valid(auto_fragmenter_out_d_valid),.auto_out_d_bits_opcode(auto_fragmenter_out_d_bits_opcode),.auto_out_d_bits_size(auto_fragmenter_out_d_bits_size),.auto_out_d_bits_source(auto_fragmenter_out_d_bits_source),.auto_out_d_bits_data(auto_fragmenter_out_d_bits_data)); 
endmodule
 
module TLMonitor_15 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [25:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [2:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [25:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [2:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [75:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [75:0] _GEN_0={69'h0,io_in_d_bits_source,2'h0} ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_0 ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [75:0] inflight_sizes_1 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_2=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_3=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_4=io_in_a_bits_address[25:16]==10'h200 ;  
   wire _GEN_5=_source_ok_T_12&io_in_a_bits_size==3'h6&_GEN_4 ;  
   wire _GEN_6=io_in_a_bits_param>3'h2 ;  
   wire _GEN_7=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_8=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_9=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_11=io_in_a_bits_size!=3'h7&_GEN_4 ;  
   wire _GEN_12=io_in_a_bits_mask!=mask ;  
   wire _GEN_13=_GEN_9&_GEN_11 ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_17=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_19=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_20=io_in_d_bits_size<3'h3 ;  
   wire _GEN_21=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_22=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_23=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_24=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_25=io_in_d_valid&d_first_1 ;  
   wire _GEN_26=_GEN_25&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&a_first_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_27={14'h0,io_in_d_bits_source} ;  
   wire _GEN_28=_GEN_26&same_cycle_resp&~reset ;  
   wire _GEN_29=_GEN_26&~same_cycle_resp&~reset ;  
   wire _GEN_30=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_31=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_32=inflight>>_GEN_27 ;  
   wire [75:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_0 ;  
   wire [18:0] _GEN_33=inflight_1>>_GEN_27 ;  
   wire [75:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_0 ;  
  always @( posedge clock)
       begin 
         if (_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_31[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~reset&~(_GEN_32[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~(_GEN_33[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CLINT.scala:108:65)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_34={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_34 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_34 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_34 ;  
   wire [258:0] _GEN_35={252'h0,io_in_a_bits_source,2'h0} ;  
   wire [31:0] _GEN_36={27'h0,io_in_d_bits_source} ;  
   wire [270:0] _GEN_37={264'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_36 ;  
   wire [31:0] _a_set_T=32'h1<<io_in_a_bits_source ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<_GEN_37 ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_35 ;  
   wire [270:0] _d_sizes_clr_T_5=271'hF<<_GEN_37 ;  
   wire [258:0] _a_sizes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_35 ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_36 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hF<<_GEN_37 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_38=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_39=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=76'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=76'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[18:0]:19'h0))&~(_GEN_38 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_38 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[75:0]:76'h0))&~(_GEN_38 ? _d_sizes_clr_T_5[75:0]:76'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_39 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_39 ? _d_sizes_clr_T_11[75:0]:76'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module Repeater_1 (
  input clock,
  input reset,
  input io_repeat,
  output io_full,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [2:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input [25:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [2:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source,
  output [25:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output io_deq_bits_corrupt) ; 
   reg full ;  
   reg [2:0] saved_opcode ;  
   reg [2:0] saved_param ;  
   reg [2:0] saved_size ;  
   reg [4:0] saved_source ;  
   reg [25:0] saved_address ;  
   reg [7:0] saved_mask ;  
   reg saved_corrupt ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire io_enq_ready_0=io_deq_ready&~full ;  
   wire _GEN=io_enq_ready_0&io_enq_valid&io_repeat ;  
  always @( posedge clock)
       begin 
         if (reset)
            full <=1'h0;
          else 
            full <=~(io_deq_ready&io_deq_valid_0&~io_repeat)&(_GEN|full);
         if (_GEN)
            begin 
              saved_opcode <=io_enq_bits_opcode;
              saved_param <=io_enq_bits_param;
              saved_size <=io_enq_bits_size;
              saved_source <=io_enq_bits_source;
              saved_address <=io_enq_bits_address;
              saved_mask <=io_enq_bits_mask;
              saved_corrupt <=io_enq_bits_corrupt;
            end 
       end
  
  assign io_full=full; 
  assign io_enq_ready=io_enq_ready_0; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_opcode=full ? saved_opcode:io_enq_bits_opcode; 
  assign io_deq_bits_param=full ? saved_param:io_enq_bits_param; 
  assign io_deq_bits_size=full ? saved_size:io_enq_bits_size; 
  assign io_deq_bits_source=full ? saved_source:io_enq_bits_source; 
  assign io_deq_bits_address=full ? saved_address:io_enq_bits_address; 
  assign io_deq_bits_mask=full ? saved_mask:io_enq_bits_mask; 
  assign io_deq_bits_corrupt=full ? saved_corrupt:io_enq_bits_corrupt; 
endmodule
 
module TLFragmenter_1 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [25:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [2:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [1:0] auto_out_a_bits_size,
  output [8:0] auto_out_a_bits_source,
  output [25:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_size,
  input [8:0] auto_out_d_bits_source,
  input [63:0] auto_out_d_bits_data) ; 
   wire _repeater_io_full ;  
   wire _repeater_io_enq_ready ;  
   wire _repeater_io_deq_valid ;  
   wire [2:0] _repeater_io_deq_bits_opcode ;  
   wire [2:0] _repeater_io_deq_bits_size ;  
   wire [4:0] _repeater_io_deq_bits_source ;  
   wire [25:0] _repeater_io_deq_bits_address ;  
   wire [7:0] _repeater_io_deq_bits_mask ;  
   reg [2:0] acknum ;  
   reg [2:0] dOrig ;  
   reg dToggle ;  
   wire dFirst=acknum==3'h0 ;  
   wire [5:0] _dsizeOH1_T_1=6'h7<<auto_out_d_bits_size ;  
   wire [2:0] _GEN=~(auto_out_d_bits_source[2:0]) ;  
   wire [2:0] dFirst_size_hi=auto_out_d_bits_source[2:0]&{1'h1,_GEN[2:1]} ;  
   wire [2:0] _dFirst_size_T_8={1'h0,dFirst_size_hi[2:1]}|~(_dsizeOH1_T_1[2:0])&{_GEN[0],_dsizeOH1_T_1[2:1]} ;  
   wire [2:0] dFirst_size={|dFirst_size_hi,|(_dFirst_size_T_8[2:1]),_dFirst_size_T_8[2]|_dFirst_size_T_8[0]} ;  
   wire drop=~(auto_out_d_bits_opcode[0])&(|(auto_out_d_bits_source[2:0])) ;  
   wire nodeOut_d_ready=auto_in_d_ready|drop ;  
   wire nodeIn_d_valid=auto_out_d_valid&~drop ;  
   wire [2:0] nodeIn_d_bits_size=dFirst ? dFirst_size:dOrig ;  
   wire [12:0] _aOrigOH1_T_1=13'h3F<<_repeater_io_deq_bits_size ;  
   reg [2:0] gennum ;  
   wire aFirst=gennum==3'h0 ;  
   wire [2:0] _old_gennum1_T_1=gennum-3'h1 ;  
   wire [2:0] aFragnum=aFirst ? ~(_aOrigOH1_T_1[5:3]):_old_gennum1_T_1 ;  
   reg aToggle_r ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~_repeater_io_full|_repeater_io_deq_bits_opcode[2]))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:311 assert (!repeater.io.full || !aHasData)\n");
              if (1)$display("");
            end 
         if (~reset&~(~_repeater_io_full|(&_repeater_io_deq_bits_mask)))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:314 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
              if (1)$display("");
            end 
       end
  
   wire _GEN_0=nodeOut_d_ready&auto_out_d_valid ;  
   wire _GEN_1=_GEN_0&dFirst ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              acknum <=3'h0;
              dToggle <=1'h0;
              gennum <=3'h0;
            end 
          else 
            begin 
              if (_GEN_0)
                 begin 
                   if (dFirst)
                      acknum <=auto_out_d_bits_source[2:0];
                    else 
                      acknum <=acknum-{2'h0,auto_out_d_bits_opcode[0]|(&auto_out_d_bits_size)};
                 end 
              if (_GEN_1)
                 dToggle <=auto_out_d_bits_source[3];
              if (auto_out_a_ready&_repeater_io_deq_valid)
                 begin 
                   if (aFirst)
                      gennum <=~(_aOrigOH1_T_1[5:3]);
                    else 
                      gennum <=_old_gennum1_T_1;
                 end 
            end 
         if (_GEN_1)
            dOrig <=dFirst_size;
         if (aFirst)
            aToggle_r <=dToggle;
       end
  
  TLMonitor_15 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_repeater_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_size(nodeIn_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source[8:4])); 
  Repeater_1 repeater(.clock(clock),.reset(reset),.io_repeat(_repeater_io_deq_bits_opcode[2]&(|aFragnum)),.io_full(_repeater_io_full),.io_enq_ready(_repeater_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_corrupt(auto_in_a_bits_corrupt),.io_deq_ready(auto_out_a_ready),.io_deq_valid(_repeater_io_deq_valid),.io_deq_bits_opcode(_repeater_io_deq_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(_repeater_io_deq_bits_size),.io_deq_bits_source(_repeater_io_deq_bits_source),.io_deq_bits_address(_repeater_io_deq_bits_address),.io_deq_bits_mask(_repeater_io_deq_bits_mask),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  assign auto_in_a_ready=_repeater_io_enq_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size=nodeIn_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source[8:4]; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_out_a_valid=_repeater_io_deq_valid; 
  assign auto_out_a_bits_opcode=_repeater_io_deq_bits_opcode; 
  assign auto_out_a_bits_size=_repeater_io_deq_bits_size[2] ? 2'h3:_repeater_io_deq_bits_size[1:0]; 
  assign auto_out_a_bits_source={_repeater_io_deq_bits_source,~(aFirst ? dToggle:aToggle_r),aFragnum}; 
  assign auto_out_a_bits_address={_repeater_io_deq_bits_address[25:6],_repeater_io_deq_bits_address[5:0]|{~(aFragnum|_aOrigOH1_T_1[5:3]),3'h0}}; 
  assign auto_out_a_bits_mask=_repeater_io_full ? 8'hFF:auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_d_ready=nodeOut_d_ready; 
endmodule
 
module TLInterconnectCoupler_8 (
  input clock,
  input reset,
  input auto_fragmenter_out_a_ready,
  output auto_fragmenter_out_a_valid,
  output [2:0] auto_fragmenter_out_a_bits_opcode,
  output [2:0] auto_fragmenter_out_a_bits_param,
  output [1:0] auto_fragmenter_out_a_bits_size,
  output [8:0] auto_fragmenter_out_a_bits_source,
  output [25:0] auto_fragmenter_out_a_bits_address,
  output [7:0] auto_fragmenter_out_a_bits_mask,
  output [63:0] auto_fragmenter_out_a_bits_data,
  output auto_fragmenter_out_a_bits_corrupt,
  output auto_fragmenter_out_d_ready,
  input auto_fragmenter_out_d_valid,
  input [2:0] auto_fragmenter_out_d_bits_opcode,
  input [1:0] auto_fragmenter_out_d_bits_size,
  input [8:0] auto_fragmenter_out_d_bits_source,
  input [63:0] auto_fragmenter_out_d_bits_data,
  output auto_tl_in_a_ready,
  input auto_tl_in_a_valid,
  input [2:0] auto_tl_in_a_bits_opcode,
  input [2:0] auto_tl_in_a_bits_param,
  input [2:0] auto_tl_in_a_bits_size,
  input [4:0] auto_tl_in_a_bits_source,
  input [25:0] auto_tl_in_a_bits_address,
  input [7:0] auto_tl_in_a_bits_mask,
  input [63:0] auto_tl_in_a_bits_data,
  input auto_tl_in_a_bits_corrupt,
  input auto_tl_in_d_ready,
  output auto_tl_in_d_valid,
  output [2:0] auto_tl_in_d_bits_opcode,
  output [2:0] auto_tl_in_d_bits_size,
  output [4:0] auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data) ; 
  TLFragmenter_1 fragmenter(.clock(clock),.reset(reset),.auto_in_a_ready(auto_tl_in_a_ready),.auto_in_a_valid(auto_tl_in_a_valid),.auto_in_a_bits_opcode(auto_tl_in_a_bits_opcode),.auto_in_a_bits_param(auto_tl_in_a_bits_param),.auto_in_a_bits_size(auto_tl_in_a_bits_size),.auto_in_a_bits_source(auto_tl_in_a_bits_source),.auto_in_a_bits_address(auto_tl_in_a_bits_address),.auto_in_a_bits_mask(auto_tl_in_a_bits_mask),.auto_in_a_bits_data(auto_tl_in_a_bits_data),.auto_in_a_bits_corrupt(auto_tl_in_a_bits_corrupt),.auto_in_d_ready(auto_tl_in_d_ready),.auto_in_d_valid(auto_tl_in_d_valid),.auto_in_d_bits_opcode(auto_tl_in_d_bits_opcode),.auto_in_d_bits_size(auto_tl_in_d_bits_size),.auto_in_d_bits_source(auto_tl_in_d_bits_source),.auto_in_d_bits_data(auto_tl_in_d_bits_data),.auto_out_a_ready(auto_fragmenter_out_a_ready),.auto_out_a_valid(auto_fragmenter_out_a_valid),.auto_out_a_bits_opcode(auto_fragmenter_out_a_bits_opcode),.auto_out_a_bits_param(auto_fragmenter_out_a_bits_param),.auto_out_a_bits_size(auto_fragmenter_out_a_bits_size),.auto_out_a_bits_source(auto_fragmenter_out_a_bits_source),.auto_out_a_bits_address(auto_fragmenter_out_a_bits_address),.auto_out_a_bits_mask(auto_fragmenter_out_a_bits_mask),.auto_out_a_bits_data(auto_fragmenter_out_a_bits_data),.auto_out_a_bits_corrupt(auto_fragmenter_out_a_bits_corrupt),.auto_out_d_ready(auto_fragmenter_out_d_ready),.auto_out_d_valid(auto_fragmenter_out_d_valid),.auto_out_d_bits_opcode(auto_fragmenter_out_d_bits_opcode),.auto_out_d_bits_size(auto_fragmenter_out_d_bits_size),.auto_out_d_bits_source(auto_fragmenter_out_d_bits_source),.auto_out_d_bits_data(auto_fragmenter_out_d_bits_data)); 
endmodule
 
module TLMonitor_16 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [11:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [2:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [11:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [2:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [75:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [75:0] _GEN_0={69'h0,io_in_d_bits_source,2'h0} ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_0 ;  
   wire _GEN_1=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [75:0] inflight_sizes_1 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_2=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_3=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_4=_source_ok_T_12&io_in_a_bits_size==3'h6 ;  
   wire _GEN_5=io_in_a_bits_param>3'h2 ;  
   wire _GEN_6=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_7=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_8=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire _GEN_9=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_10=io_in_a_bits_size!=3'h7 ;  
   wire _GEN_11=io_in_a_bits_mask!=mask ;  
   wire _GEN_12=_GEN_8&_GEN_10 ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_17=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_18=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_19=io_in_d_bits_size<3'h3 ;  
   wire _GEN_20=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_21=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_22=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_23=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_24=io_in_d_valid&d_first_1 ;  
   wire _GEN_25=_GEN_24&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&a_first_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_26={14'h0,io_in_d_bits_source} ;  
   wire _GEN_27=_GEN_25&same_cycle_resp&~reset ;  
   wire _GEN_28=_GEN_25&~same_cycle_resp&~reset ;  
   wire _GEN_29=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [18:0] _GEN_30=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_31=inflight>>_GEN_26 ;  
   wire [75:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_0 ;  
   wire [18:0] _GEN_32=inflight_1>>_GEN_26 ;  
   wire [75:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_0 ;  
  always @( posedge clock)
       begin 
         if (_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|_GEN_2))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_30[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~reset&~(_GEN_31[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~(_GEN_32[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Periphery.scala:87:63)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_33={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_33 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_33 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_33 ;  
   wire [258:0] _GEN_34={252'h0,io_in_a_bits_source,2'h0} ;  
   wire [31:0] _GEN_35={27'h0,io_in_d_bits_source} ;  
   wire [270:0] _GEN_36={264'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_35 ;  
   wire [31:0] _a_set_T=32'h1<<io_in_a_bits_source ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<_GEN_36 ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_34 ;  
   wire [270:0] _d_sizes_clr_T_5=271'hF<<_GEN_36 ;  
   wire [258:0] _a_sizes_set_T_1={255'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_34 ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_35 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hF<<_GEN_36 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_37=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_38=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=76'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=76'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[18:0]:19'h0))&~(_GEN_37 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_37 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[75:0]:76'h0))&~(_GEN_37 ? _d_sizes_clr_T_5[75:0]:76'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_38 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_38 ? _d_sizes_clr_T_11[75:0]:76'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module Repeater_2 (
  input clock,
  input reset,
  input io_repeat,
  output io_full,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [2:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input [11:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [2:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source,
  output [11:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output io_deq_bits_corrupt) ; 
   reg full ;  
   reg [2:0] saved_opcode ;  
   reg [2:0] saved_param ;  
   reg [2:0] saved_size ;  
   reg [4:0] saved_source ;  
   reg [11:0] saved_address ;  
   reg [7:0] saved_mask ;  
   reg saved_corrupt ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire io_enq_ready_0=io_deq_ready&~full ;  
   wire _GEN=io_enq_ready_0&io_enq_valid&io_repeat ;  
  always @( posedge clock)
       begin 
         if (reset)
            full <=1'h0;
          else 
            full <=~(io_deq_ready&io_deq_valid_0&~io_repeat)&(_GEN|full);
         if (_GEN)
            begin 
              saved_opcode <=io_enq_bits_opcode;
              saved_param <=io_enq_bits_param;
              saved_size <=io_enq_bits_size;
              saved_source <=io_enq_bits_source;
              saved_address <=io_enq_bits_address;
              saved_mask <=io_enq_bits_mask;
              saved_corrupt <=io_enq_bits_corrupt;
            end 
       end
  
  assign io_full=full; 
  assign io_enq_ready=io_enq_ready_0; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_opcode=full ? saved_opcode:io_enq_bits_opcode; 
  assign io_deq_bits_param=full ? saved_param:io_enq_bits_param; 
  assign io_deq_bits_size=full ? saved_size:io_enq_bits_size; 
  assign io_deq_bits_source=full ? saved_source:io_enq_bits_source; 
  assign io_deq_bits_address=full ? saved_address:io_enq_bits_address; 
  assign io_deq_bits_mask=full ? saved_mask:io_enq_bits_mask; 
  assign io_deq_bits_corrupt=full ? saved_corrupt:io_enq_bits_corrupt; 
endmodule
 
module TLFragmenter_2 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [11:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [2:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [1:0] auto_out_a_bits_size,
  output [8:0] auto_out_a_bits_source,
  output [11:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_size,
  input [8:0] auto_out_d_bits_source,
  input [63:0] auto_out_d_bits_data) ; 
   wire _repeater_io_full ;  
   wire _repeater_io_enq_ready ;  
   wire _repeater_io_deq_valid ;  
   wire [2:0] _repeater_io_deq_bits_opcode ;  
   wire [2:0] _repeater_io_deq_bits_size ;  
   wire [4:0] _repeater_io_deq_bits_source ;  
   wire [11:0] _repeater_io_deq_bits_address ;  
   wire [7:0] _repeater_io_deq_bits_mask ;  
   reg [2:0] acknum ;  
   reg [2:0] dOrig ;  
   reg dToggle ;  
   wire dFirst=acknum==3'h0 ;  
   wire [5:0] _dsizeOH1_T_1=6'h7<<auto_out_d_bits_size ;  
   wire [2:0] _GEN=~(auto_out_d_bits_source[2:0]) ;  
   wire [2:0] dFirst_size_hi=auto_out_d_bits_source[2:0]&{1'h1,_GEN[2:1]} ;  
   wire [2:0] _dFirst_size_T_8={1'h0,dFirst_size_hi[2:1]}|~(_dsizeOH1_T_1[2:0])&{_GEN[0],_dsizeOH1_T_1[2:1]} ;  
   wire [2:0] dFirst_size={|dFirst_size_hi,|(_dFirst_size_T_8[2:1]),_dFirst_size_T_8[2]|_dFirst_size_T_8[0]} ;  
   wire drop=~(auto_out_d_bits_opcode[0])&(|(auto_out_d_bits_source[2:0])) ;  
   wire nodeOut_d_ready=auto_in_d_ready|drop ;  
   wire nodeIn_d_valid=auto_out_d_valid&~drop ;  
   wire [2:0] nodeIn_d_bits_size=dFirst ? dFirst_size:dOrig ;  
   wire [12:0] _aOrigOH1_T_1=13'h3F<<_repeater_io_deq_bits_size ;  
   reg [2:0] gennum ;  
   wire aFirst=gennum==3'h0 ;  
   wire [2:0] _old_gennum1_T_1=gennum-3'h1 ;  
   wire [2:0] aFragnum=aFirst ? ~(_aOrigOH1_T_1[5:3]):_old_gennum1_T_1 ;  
   reg aToggle_r ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~_repeater_io_full|_repeater_io_deq_bits_opcode[2]))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:311 assert (!repeater.io.full || !aHasData)\n");
              if (1)$display("");
            end 
         if (~reset&~(~_repeater_io_full|(&_repeater_io_deq_bits_mask)))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:314 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
              if (1)$display("");
            end 
       end
  
   wire _GEN_0=nodeOut_d_ready&auto_out_d_valid ;  
   wire _GEN_1=_GEN_0&dFirst ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              acknum <=3'h0;
              dToggle <=1'h0;
              gennum <=3'h0;
            end 
          else 
            begin 
              if (_GEN_0)
                 begin 
                   if (dFirst)
                      acknum <=auto_out_d_bits_source[2:0];
                    else 
                      acknum <=acknum-{2'h0,auto_out_d_bits_opcode[0]|(&auto_out_d_bits_size)};
                 end 
              if (_GEN_1)
                 dToggle <=auto_out_d_bits_source[3];
              if (auto_out_a_ready&_repeater_io_deq_valid)
                 begin 
                   if (aFirst)
                      gennum <=~(_aOrigOH1_T_1[5:3]);
                    else 
                      gennum <=_old_gennum1_T_1;
                 end 
            end 
         if (_GEN_1)
            dOrig <=dFirst_size;
         if (aFirst)
            aToggle_r <=dToggle;
       end
  
  TLMonitor_16 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_repeater_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_size(nodeIn_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source[8:4])); 
  Repeater_2 repeater(.clock(clock),.reset(reset),.io_repeat(_repeater_io_deq_bits_opcode[2]&(|aFragnum)),.io_full(_repeater_io_full),.io_enq_ready(_repeater_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_corrupt(auto_in_a_bits_corrupt),.io_deq_ready(auto_out_a_ready),.io_deq_valid(_repeater_io_deq_valid),.io_deq_bits_opcode(_repeater_io_deq_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(_repeater_io_deq_bits_size),.io_deq_bits_source(_repeater_io_deq_bits_source),.io_deq_bits_address(_repeater_io_deq_bits_address),.io_deq_bits_mask(_repeater_io_deq_bits_mask),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  assign auto_in_a_ready=_repeater_io_enq_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size=nodeIn_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source[8:4]; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_out_a_valid=_repeater_io_deq_valid; 
  assign auto_out_a_bits_opcode=_repeater_io_deq_bits_opcode; 
  assign auto_out_a_bits_size=_repeater_io_deq_bits_size[2] ? 2'h3:_repeater_io_deq_bits_size[1:0]; 
  assign auto_out_a_bits_source={_repeater_io_deq_bits_source,~(aFirst ? dToggle:aToggle_r),aFragnum}; 
  assign auto_out_a_bits_address={_repeater_io_deq_bits_address[11:6],_repeater_io_deq_bits_address[5:0]|{~(aFragnum|_aOrigOH1_T_1[5:3]),3'h0}}; 
  assign auto_out_a_bits_mask=_repeater_io_full ? 8'hFF:auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_d_ready=nodeOut_d_ready; 
endmodule
 
module TLInterconnectCoupler_10 (
  input clock,
  input reset,
  input auto_fragmenter_out_a_ready,
  output auto_fragmenter_out_a_valid,
  output [2:0] auto_fragmenter_out_a_bits_opcode,
  output [2:0] auto_fragmenter_out_a_bits_param,
  output [1:0] auto_fragmenter_out_a_bits_size,
  output [8:0] auto_fragmenter_out_a_bits_source,
  output [11:0] auto_fragmenter_out_a_bits_address,
  output [7:0] auto_fragmenter_out_a_bits_mask,
  output [63:0] auto_fragmenter_out_a_bits_data,
  output auto_fragmenter_out_a_bits_corrupt,
  output auto_fragmenter_out_d_ready,
  input auto_fragmenter_out_d_valid,
  input [2:0] auto_fragmenter_out_d_bits_opcode,
  input [1:0] auto_fragmenter_out_d_bits_size,
  input [8:0] auto_fragmenter_out_d_bits_source,
  input [63:0] auto_fragmenter_out_d_bits_data,
  output auto_tl_in_a_ready,
  input auto_tl_in_a_valid,
  input [2:0] auto_tl_in_a_bits_opcode,
  input [2:0] auto_tl_in_a_bits_param,
  input [2:0] auto_tl_in_a_bits_size,
  input [4:0] auto_tl_in_a_bits_source,
  input [11:0] auto_tl_in_a_bits_address,
  input [7:0] auto_tl_in_a_bits_mask,
  input [63:0] auto_tl_in_a_bits_data,
  input auto_tl_in_a_bits_corrupt,
  input auto_tl_in_d_ready,
  output auto_tl_in_d_valid,
  output [2:0] auto_tl_in_d_bits_opcode,
  output [2:0] auto_tl_in_d_bits_size,
  output [4:0] auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data) ; 
  TLFragmenter_2 fragmenter(.clock(clock),.reset(reset),.auto_in_a_ready(auto_tl_in_a_ready),.auto_in_a_valid(auto_tl_in_a_valid),.auto_in_a_bits_opcode(auto_tl_in_a_bits_opcode),.auto_in_a_bits_param(auto_tl_in_a_bits_param),.auto_in_a_bits_size(auto_tl_in_a_bits_size),.auto_in_a_bits_source(auto_tl_in_a_bits_source),.auto_in_a_bits_address(auto_tl_in_a_bits_address),.auto_in_a_bits_mask(auto_tl_in_a_bits_mask),.auto_in_a_bits_data(auto_tl_in_a_bits_data),.auto_in_a_bits_corrupt(auto_tl_in_a_bits_corrupt),.auto_in_d_ready(auto_tl_in_d_ready),.auto_in_d_valid(auto_tl_in_d_valid),.auto_in_d_bits_opcode(auto_tl_in_d_bits_opcode),.auto_in_d_bits_size(auto_tl_in_d_bits_size),.auto_in_d_bits_source(auto_tl_in_d_bits_source),.auto_in_d_bits_data(auto_tl_in_d_bits_data),.auto_out_a_ready(auto_fragmenter_out_a_ready),.auto_out_a_valid(auto_fragmenter_out_a_valid),.auto_out_a_bits_opcode(auto_fragmenter_out_a_bits_opcode),.auto_out_a_bits_param(auto_fragmenter_out_a_bits_param),.auto_out_a_bits_size(auto_fragmenter_out_a_bits_size),.auto_out_a_bits_source(auto_fragmenter_out_a_bits_source),.auto_out_a_bits_address(auto_fragmenter_out_a_bits_address),.auto_out_a_bits_mask(auto_fragmenter_out_a_bits_mask),.auto_out_a_bits_data(auto_fragmenter_out_a_bits_data),.auto_out_a_bits_corrupt(auto_fragmenter_out_a_bits_corrupt),.auto_out_d_ready(auto_fragmenter_out_d_ready),.auto_out_d_valid(auto_fragmenter_out_d_valid),.auto_out_d_bits_opcode(auto_fragmenter_out_d_bits_opcode),.auto_out_d_bits_size(auto_fragmenter_out_d_bits_size),.auto_out_d_bits_source(auto_fragmenter_out_d_bits_source),.auto_out_d_bits_data(auto_fragmenter_out_d_bits_data)); 
endmodule
 
module TLMonitor_17 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [16:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [16:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [75:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [75:0] _GEN={69'h0,io_in_d_bits_source,2'h0} ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire _GEN_0=a_first_done&a_first_1 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<io_in_a_bits_size ;  
   wire [5:0] _GEN_1=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_3=_source_ok_T_12&io_in_a_bits_size==3'h6&io_in_a_bits_address[16] ;  
   wire _GEN_4=io_in_a_bits_param>3'h2 ;  
   wire _GEN_5=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_6=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_7=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_8=io_in_a_bits_mask!=mask ;  
   wire _GEN_9=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_14=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_15=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_16=io_in_d_valid&d_first_1 ;  
   wire same_cycle_resp=io_in_a_valid&a_first_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_17=_GEN_16&same_cycle_resp&~reset ;  
   wire _GEN_18=_GEN_16&~same_cycle_resp&~reset ;  
   wire [18:0] _GEN_19=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_20=inflight>>io_in_d_bits_source ;  
   wire [75:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~(~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~(io_in_a_bits_size!=3'h7&io_in_a_bits_address[16]))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&~(io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&_GEN_19[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~reset&~(_GEN_20[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~(casez_tmp==3'h1|casez_tmp_0==3'h1))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~(casez_tmp_1==3'h1|casez_tmp_2==3'h1))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/BootROM.scala:86:68)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _GEN_21={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_21 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_21 ;  
   wire [258:0] _GEN_22={252'h0,io_in_a_bits_source,2'h0} ;  
   wire [270:0] _GEN_23={264'h0,io_in_d_bits_source,2'h0} ;  
   wire [31:0] _d_clr_T=32'h1<<io_in_d_bits_source ;  
   wire [31:0] _a_set_T=32'h1<<io_in_a_bits_source ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<_GEN_23 ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_0 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_22 ;  
   wire [270:0] _d_sizes_clr_T_5=271'hF<<_GEN_23 ;  
   wire [258:0] _a_sizes_set_T_1={255'h0,_GEN_0 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_22 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_24=_d_first_T_2&d_first_1 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=76'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
            end 
          else 
            begin 
              if (a_first_done)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=3'h0;
                   if (a_first_1)
                      a_first_counter_1 <=3'h0;
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=~(_d_first_beats1_decode_T_1[5:3]);
                   if (d_first_1)
                      d_first_counter_1 <=~(_d_first_beats1_decode_T_5[5:3]);
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                 end 
              inflight <=(inflight|(_GEN_0 ? _a_set_T[18:0]:19'h0))&~(_GEN_24 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_0 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_24 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_0 ? _a_sizes_set_T_1[75:0]:76'h0))&~(_GEN_24 ? _d_sizes_clr_T_5[75:0]:76'h0);
              if (a_first_done|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
            end 
         if (a_first_done&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module Repeater_3 (
  input clock,
  input reset,
  input io_repeat,
  output io_full,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [2:0] io_enq_bits_size,
  input [4:0] io_enq_bits_source,
  input [16:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [2:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source,
  output [16:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output io_deq_bits_corrupt) ; 
   reg full ;  
   reg [2:0] saved_opcode ;  
   reg [2:0] saved_param ;  
   reg [2:0] saved_size ;  
   reg [4:0] saved_source ;  
   reg [16:0] saved_address ;  
   reg [7:0] saved_mask ;  
   reg saved_corrupt ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire io_enq_ready_0=io_deq_ready&~full ;  
   wire _GEN=io_enq_ready_0&io_enq_valid&io_repeat ;  
  always @( posedge clock)
       begin 
         if (reset)
            full <=1'h0;
          else 
            full <=~(io_deq_ready&io_deq_valid_0&~io_repeat)&(_GEN|full);
         if (_GEN)
            begin 
              saved_opcode <=io_enq_bits_opcode;
              saved_param <=io_enq_bits_param;
              saved_size <=io_enq_bits_size;
              saved_source <=io_enq_bits_source;
              saved_address <=io_enq_bits_address;
              saved_mask <=io_enq_bits_mask;
              saved_corrupt <=io_enq_bits_corrupt;
            end 
       end
  
  assign io_full=full; 
  assign io_enq_ready=io_enq_ready_0; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_opcode=full ? saved_opcode:io_enq_bits_opcode; 
  assign io_deq_bits_param=full ? saved_param:io_enq_bits_param; 
  assign io_deq_bits_size=full ? saved_size:io_enq_bits_size; 
  assign io_deq_bits_source=full ? saved_source:io_enq_bits_source; 
  assign io_deq_bits_address=full ? saved_address:io_enq_bits_address; 
  assign io_deq_bits_mask=full ? saved_mask:io_enq_bits_mask; 
  assign io_deq_bits_corrupt=full ? saved_corrupt:io_enq_bits_corrupt; 
endmodule
 
module TLFragmenter_3 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [16:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [1:0] auto_out_a_bits_size,
  output [8:0] auto_out_a_bits_source,
  output [16:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [1:0] auto_out_d_bits_size,
  input [8:0] auto_out_d_bits_source,
  input [63:0] auto_out_d_bits_data) ; 
   wire _repeater_io_full ;  
   wire _repeater_io_enq_ready ;  
   wire _repeater_io_deq_valid ;  
   wire [2:0] _repeater_io_deq_bits_size ;  
   wire [4:0] _repeater_io_deq_bits_source ;  
   wire [16:0] _repeater_io_deq_bits_address ;  
   wire [7:0] _repeater_io_deq_bits_mask ;  
   reg [2:0] acknum ;  
   reg [2:0] dOrig ;  
   reg dToggle ;  
   wire dFirst=acknum==3'h0 ;  
   wire [5:0] _dsizeOH1_T_1=6'h7<<auto_out_d_bits_size ;  
   wire [2:0] _GEN=~(auto_out_d_bits_source[2:0]) ;  
   wire [2:0] dFirst_size_hi=auto_out_d_bits_source[2:0]&{1'h1,_GEN[2:1]} ;  
   wire [2:0] _dFirst_size_T_8={1'h0,dFirst_size_hi[2:1]}|~(_dsizeOH1_T_1[2:0])&{_GEN[0],_dsizeOH1_T_1[2:1]} ;  
   wire [2:0] dFirst_size={|dFirst_size_hi,|(_dFirst_size_T_8[2:1]),_dFirst_size_T_8[2]|_dFirst_size_T_8[0]} ;  
   wire [2:0] nodeIn_d_bits_size=dFirst ? dFirst_size:dOrig ;  
   wire [12:0] _aOrigOH1_T_1=13'h3F<<_repeater_io_deq_bits_size ;  
   reg [2:0] gennum ;  
   wire aFirst=gennum==3'h0 ;  
   wire [2:0] _old_gennum1_T_1=gennum-3'h1 ;  
   wire [2:0] aFragnum=aFirst ? ~(_aOrigOH1_T_1[5:3]):_old_gennum1_T_1 ;  
   reg aToggle_r ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~_repeater_io_full|(&_repeater_io_deq_bits_mask)))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:314 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
              if (1)$display("");
            end 
       end
  
   wire _GEN_0=auto_in_d_ready&auto_out_d_valid ;  
   wire _GEN_1=_GEN_0&dFirst ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              acknum <=3'h0;
              dToggle <=1'h0;
              gennum <=3'h0;
            end 
          else 
            begin 
              if (_GEN_0)
                 begin 
                   if (dFirst)
                      acknum <=auto_out_d_bits_source[2:0];
                    else 
                      acknum <=acknum-3'h1;
                 end 
              if (_GEN_1)
                 dToggle <=auto_out_d_bits_source[3];
              if (auto_out_a_ready&_repeater_io_deq_valid)
                 begin 
                   if (aFirst)
                      gennum <=~(_aOrigOH1_T_1[5:3]);
                    else 
                      gennum <=_old_gennum1_T_1;
                 end 
            end 
         if (_GEN_1)
            dOrig <=dFirst_size;
         if (aFirst)
            aToggle_r <=dToggle;
       end
  
  TLMonitor_17 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_repeater_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_out_d_valid),.io_in_d_bits_size(nodeIn_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source[8:4])); 
  Repeater_3 repeater(.clock(clock),.reset(reset),.io_repeat(|aFragnum),.io_full(_repeater_io_full),.io_enq_ready(_repeater_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_corrupt(auto_in_a_bits_corrupt),.io_deq_ready(auto_out_a_ready),.io_deq_valid(_repeater_io_deq_valid),.io_deq_bits_opcode(auto_out_a_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(_repeater_io_deq_bits_size),.io_deq_bits_source(_repeater_io_deq_bits_source),.io_deq_bits_address(_repeater_io_deq_bits_address),.io_deq_bits_mask(_repeater_io_deq_bits_mask),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  assign auto_in_a_ready=_repeater_io_enq_ready; 
  assign auto_in_d_valid=auto_out_d_valid; 
  assign auto_in_d_bits_size=nodeIn_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source[8:4]; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_out_a_valid=_repeater_io_deq_valid; 
  assign auto_out_a_bits_size=_repeater_io_deq_bits_size[2] ? 2'h3:_repeater_io_deq_bits_size[1:0]; 
  assign auto_out_a_bits_source={_repeater_io_deq_bits_source,~(aFirst ? dToggle:aToggle_r),aFragnum}; 
  assign auto_out_a_bits_address={_repeater_io_deq_bits_address[16:6],_repeater_io_deq_bits_address[5:0]|{~(aFragnum|_aOrigOH1_T_1[5:3]),3'h0}}; 
  assign auto_out_a_bits_mask=_repeater_io_full ? 8'hFF:auto_in_a_bits_mask; 
  assign auto_out_d_ready=auto_in_d_ready; 
endmodule
 
module TLInterconnectCoupler_11 (
  input clock,
  input reset,
  input auto_fragmenter_out_a_ready,
  output auto_fragmenter_out_a_valid,
  output [2:0] auto_fragmenter_out_a_bits_opcode,
  output [2:0] auto_fragmenter_out_a_bits_param,
  output [1:0] auto_fragmenter_out_a_bits_size,
  output [8:0] auto_fragmenter_out_a_bits_source,
  output [16:0] auto_fragmenter_out_a_bits_address,
  output [7:0] auto_fragmenter_out_a_bits_mask,
  output auto_fragmenter_out_a_bits_corrupt,
  output auto_fragmenter_out_d_ready,
  input auto_fragmenter_out_d_valid,
  input [1:0] auto_fragmenter_out_d_bits_size,
  input [8:0] auto_fragmenter_out_d_bits_source,
  input [63:0] auto_fragmenter_out_d_bits_data,
  output auto_tl_in_a_ready,
  input auto_tl_in_a_valid,
  input [2:0] auto_tl_in_a_bits_opcode,
  input [2:0] auto_tl_in_a_bits_param,
  input [2:0] auto_tl_in_a_bits_size,
  input [4:0] auto_tl_in_a_bits_source,
  input [16:0] auto_tl_in_a_bits_address,
  input [7:0] auto_tl_in_a_bits_mask,
  input auto_tl_in_a_bits_corrupt,
  input auto_tl_in_d_ready,
  output auto_tl_in_d_valid,
  output [2:0] auto_tl_in_d_bits_size,
  output [4:0] auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data) ; 
  TLFragmenter_3 fragmenter(.clock(clock),.reset(reset),.auto_in_a_ready(auto_tl_in_a_ready),.auto_in_a_valid(auto_tl_in_a_valid),.auto_in_a_bits_opcode(auto_tl_in_a_bits_opcode),.auto_in_a_bits_param(auto_tl_in_a_bits_param),.auto_in_a_bits_size(auto_tl_in_a_bits_size),.auto_in_a_bits_source(auto_tl_in_a_bits_source),.auto_in_a_bits_address(auto_tl_in_a_bits_address),.auto_in_a_bits_mask(auto_tl_in_a_bits_mask),.auto_in_a_bits_corrupt(auto_tl_in_a_bits_corrupt),.auto_in_d_ready(auto_tl_in_d_ready),.auto_in_d_valid(auto_tl_in_d_valid),.auto_in_d_bits_size(auto_tl_in_d_bits_size),.auto_in_d_bits_source(auto_tl_in_d_bits_source),.auto_in_d_bits_data(auto_tl_in_d_bits_data),.auto_out_a_ready(auto_fragmenter_out_a_ready),.auto_out_a_valid(auto_fragmenter_out_a_valid),.auto_out_a_bits_opcode(auto_fragmenter_out_a_bits_opcode),.auto_out_a_bits_param(auto_fragmenter_out_a_bits_param),.auto_out_a_bits_size(auto_fragmenter_out_a_bits_size),.auto_out_a_bits_source(auto_fragmenter_out_a_bits_source),.auto_out_a_bits_address(auto_fragmenter_out_a_bits_address),.auto_out_a_bits_mask(auto_fragmenter_out_a_bits_mask),.auto_out_a_bits_corrupt(auto_fragmenter_out_a_bits_corrupt),.auto_out_d_ready(auto_fragmenter_out_d_ready),.auto_out_d_valid(auto_fragmenter_out_d_valid),.auto_out_d_bits_size(auto_fragmenter_out_d_bits_size),.auto_out_d_bits_source(auto_fragmenter_out_d_bits_source),.auto_out_d_bits_data(auto_fragmenter_out_d_bits_data)); 
endmodule
 
module PeripheryBus_1 (
  input auto_coupler_to_bootrom_fragmenter_out_a_ready,
  output auto_coupler_to_bootrom_fragmenter_out_a_valid,
  output [2:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode,
  output [2:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_param,
  output [1:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_size,
  output [8:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_source,
  output [16:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_address,
  output [7:0] auto_coupler_to_bootrom_fragmenter_out_a_bits_mask,
  output auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt,
  output auto_coupler_to_bootrom_fragmenter_out_d_ready,
  input auto_coupler_to_bootrom_fragmenter_out_d_valid,
  input [1:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_size,
  input [8:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_source,
  input [63:0] auto_coupler_to_bootrom_fragmenter_out_d_bits_data,
  input auto_coupler_to_debug_fragmenter_out_a_ready,
  output auto_coupler_to_debug_fragmenter_out_a_valid,
  output [2:0] auto_coupler_to_debug_fragmenter_out_a_bits_opcode,
  output [2:0] auto_coupler_to_debug_fragmenter_out_a_bits_param,
  output [1:0] auto_coupler_to_debug_fragmenter_out_a_bits_size,
  output [8:0] auto_coupler_to_debug_fragmenter_out_a_bits_source,
  output [11:0] auto_coupler_to_debug_fragmenter_out_a_bits_address,
  output [7:0] auto_coupler_to_debug_fragmenter_out_a_bits_mask,
  output [63:0] auto_coupler_to_debug_fragmenter_out_a_bits_data,
  output auto_coupler_to_debug_fragmenter_out_a_bits_corrupt,
  output auto_coupler_to_debug_fragmenter_out_d_ready,
  input auto_coupler_to_debug_fragmenter_out_d_valid,
  input [2:0] auto_coupler_to_debug_fragmenter_out_d_bits_opcode,
  input [1:0] auto_coupler_to_debug_fragmenter_out_d_bits_size,
  input [8:0] auto_coupler_to_debug_fragmenter_out_d_bits_source,
  input [63:0] auto_coupler_to_debug_fragmenter_out_d_bits_data,
  input auto_coupler_to_clint_fragmenter_out_a_ready,
  output auto_coupler_to_clint_fragmenter_out_a_valid,
  output [2:0] auto_coupler_to_clint_fragmenter_out_a_bits_opcode,
  output [2:0] auto_coupler_to_clint_fragmenter_out_a_bits_param,
  output [1:0] auto_coupler_to_clint_fragmenter_out_a_bits_size,
  output [8:0] auto_coupler_to_clint_fragmenter_out_a_bits_source,
  output [25:0] auto_coupler_to_clint_fragmenter_out_a_bits_address,
  output [7:0] auto_coupler_to_clint_fragmenter_out_a_bits_mask,
  output [63:0] auto_coupler_to_clint_fragmenter_out_a_bits_data,
  output auto_coupler_to_clint_fragmenter_out_a_bits_corrupt,
  output auto_coupler_to_clint_fragmenter_out_d_ready,
  input auto_coupler_to_clint_fragmenter_out_d_valid,
  input [2:0] auto_coupler_to_clint_fragmenter_out_d_bits_opcode,
  input [1:0] auto_coupler_to_clint_fragmenter_out_d_bits_size,
  input [8:0] auto_coupler_to_clint_fragmenter_out_d_bits_source,
  input [63:0] auto_coupler_to_clint_fragmenter_out_d_bits_data,
  input auto_coupler_to_plic_fragmenter_out_a_ready,
  output auto_coupler_to_plic_fragmenter_out_a_valid,
  output [2:0] auto_coupler_to_plic_fragmenter_out_a_bits_opcode,
  output [2:0] auto_coupler_to_plic_fragmenter_out_a_bits_param,
  output [1:0] auto_coupler_to_plic_fragmenter_out_a_bits_size,
  output [8:0] auto_coupler_to_plic_fragmenter_out_a_bits_source,
  output [27:0] auto_coupler_to_plic_fragmenter_out_a_bits_address,
  output [7:0] auto_coupler_to_plic_fragmenter_out_a_bits_mask,
  output [63:0] auto_coupler_to_plic_fragmenter_out_a_bits_data,
  output auto_coupler_to_plic_fragmenter_out_a_bits_corrupt,
  output auto_coupler_to_plic_fragmenter_out_d_ready,
  input auto_coupler_to_plic_fragmenter_out_d_valid,
  input [2:0] auto_coupler_to_plic_fragmenter_out_d_bits_opcode,
  input [1:0] auto_coupler_to_plic_fragmenter_out_d_bits_size,
  input [8:0] auto_coupler_to_plic_fragmenter_out_d_bits_source,
  input [63:0] auto_coupler_to_plic_fragmenter_out_d_bits_data,
  output auto_fixedClockNode_out_2_clock,
  output auto_fixedClockNode_out_2_reset,
  output auto_fixedClockNode_out_0_clock,
  output auto_fixedClockNode_out_0_reset,
  input auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock,
  input auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset,
  input auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock,
  input auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset,
  output auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock,
  output auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset,
  output auto_bus_xing_in_a_ready,
  input auto_bus_xing_in_a_valid,
  input [2:0] auto_bus_xing_in_a_bits_opcode,
  input [2:0] auto_bus_xing_in_a_bits_param,
  input [3:0] auto_bus_xing_in_a_bits_size,
  input [4:0] auto_bus_xing_in_a_bits_source,
  input [27:0] auto_bus_xing_in_a_bits_address,
  input [7:0] auto_bus_xing_in_a_bits_mask,
  input [63:0] auto_bus_xing_in_a_bits_data,
  input auto_bus_xing_in_a_bits_corrupt,
  input auto_bus_xing_in_d_ready,
  output auto_bus_xing_in_d_valid,
  output [2:0] auto_bus_xing_in_d_bits_opcode,
  output [1:0] auto_bus_xing_in_d_bits_param,
  output [3:0] auto_bus_xing_in_d_bits_size,
  output [4:0] auto_bus_xing_in_d_bits_source,
  output auto_bus_xing_in_d_bits_sink,
  output auto_bus_xing_in_d_bits_denied,
  output [63:0] auto_bus_xing_in_d_bits_data,
  output auto_bus_xing_in_d_bits_corrupt,
  output clock,
  output reset) ; 
   wire _coupler_to_bootrom_auto_tl_in_a_ready ;  
   wire _coupler_to_bootrom_auto_tl_in_d_valid ;  
   wire [2:0] _coupler_to_bootrom_auto_tl_in_d_bits_size ;  
   wire [4:0] _coupler_to_bootrom_auto_tl_in_d_bits_source ;  
   wire [63:0] _coupler_to_bootrom_auto_tl_in_d_bits_data ;  
   wire _coupler_to_debug_auto_tl_in_a_ready ;  
   wire _coupler_to_debug_auto_tl_in_d_valid ;  
   wire [2:0] _coupler_to_debug_auto_tl_in_d_bits_opcode ;  
   wire [2:0] _coupler_to_debug_auto_tl_in_d_bits_size ;  
   wire [4:0] _coupler_to_debug_auto_tl_in_d_bits_source ;  
   wire [63:0] _coupler_to_debug_auto_tl_in_d_bits_data ;  
   wire _coupler_to_clint_auto_tl_in_a_ready ;  
   wire _coupler_to_clint_auto_tl_in_d_valid ;  
   wire [2:0] _coupler_to_clint_auto_tl_in_d_bits_opcode ;  
   wire [2:0] _coupler_to_clint_auto_tl_in_d_bits_size ;  
   wire [4:0] _coupler_to_clint_auto_tl_in_d_bits_source ;  
   wire [63:0] _coupler_to_clint_auto_tl_in_d_bits_data ;  
   wire _coupler_to_plic_auto_tl_in_a_ready ;  
   wire _coupler_to_plic_auto_tl_in_d_valid ;  
   wire [2:0] _coupler_to_plic_auto_tl_in_d_bits_opcode ;  
   wire [2:0] _coupler_to_plic_auto_tl_in_d_bits_size ;  
   wire [4:0] _coupler_to_plic_auto_tl_in_d_bits_source ;  
   wire [63:0] _coupler_to_plic_auto_tl_in_d_bits_data ;  
   wire _wrapped_error_device_auto_buffer_in_a_ready ;  
   wire _wrapped_error_device_auto_buffer_in_d_valid ;  
   wire [2:0] _wrapped_error_device_auto_buffer_in_d_bits_opcode ;  
   wire [1:0] _wrapped_error_device_auto_buffer_in_d_bits_param ;  
   wire [3:0] _wrapped_error_device_auto_buffer_in_d_bits_size ;  
   wire [4:0] _wrapped_error_device_auto_buffer_in_d_bits_source ;  
   wire _wrapped_error_device_auto_buffer_in_d_bits_sink ;  
   wire _wrapped_error_device_auto_buffer_in_d_bits_denied ;  
   wire [63:0] _wrapped_error_device_auto_buffer_in_d_bits_data ;  
   wire _wrapped_error_device_auto_buffer_in_d_bits_corrupt ;  
   wire _atomics_auto_out_a_valid ;  
   wire [2:0] _atomics_auto_out_a_bits_opcode ;  
   wire [2:0] _atomics_auto_out_a_bits_param ;  
   wire [3:0] _atomics_auto_out_a_bits_size ;  
   wire [4:0] _atomics_auto_out_a_bits_source ;  
   wire [27:0] _atomics_auto_out_a_bits_address ;  
   wire [7:0] _atomics_auto_out_a_bits_mask ;  
   wire [63:0] _atomics_auto_out_a_bits_data ;  
   wire _atomics_auto_out_a_bits_corrupt ;  
   wire _atomics_auto_out_d_ready ;  
   wire _buffer_auto_in_a_ready ;  
   wire _buffer_auto_in_d_valid ;  
   wire [2:0] _buffer_auto_in_d_bits_opcode ;  
   wire [1:0] _buffer_auto_in_d_bits_param ;  
   wire [3:0] _buffer_auto_in_d_bits_size ;  
   wire [4:0] _buffer_auto_in_d_bits_source ;  
   wire _buffer_auto_in_d_bits_sink ;  
   wire _buffer_auto_in_d_bits_denied ;  
   wire [63:0] _buffer_auto_in_d_bits_data ;  
   wire _buffer_auto_in_d_bits_corrupt ;  
   wire _buffer_auto_out_a_valid ;  
   wire [2:0] _buffer_auto_out_a_bits_opcode ;  
   wire [2:0] _buffer_auto_out_a_bits_param ;  
   wire [3:0] _buffer_auto_out_a_bits_size ;  
   wire [4:0] _buffer_auto_out_a_bits_source ;  
   wire [27:0] _buffer_auto_out_a_bits_address ;  
   wire [7:0] _buffer_auto_out_a_bits_mask ;  
   wire [63:0] _buffer_auto_out_a_bits_data ;  
   wire _buffer_auto_out_a_bits_corrupt ;  
   wire _buffer_auto_out_d_ready ;  
   wire _out_xbar_auto_in_a_ready ;  
   wire _out_xbar_auto_in_d_valid ;  
   wire [2:0] _out_xbar_auto_in_d_bits_opcode ;  
   wire [1:0] _out_xbar_auto_in_d_bits_param ;  
   wire [3:0] _out_xbar_auto_in_d_bits_size ;  
   wire [4:0] _out_xbar_auto_in_d_bits_source ;  
   wire _out_xbar_auto_in_d_bits_sink ;  
   wire _out_xbar_auto_in_d_bits_denied ;  
   wire [63:0] _out_xbar_auto_in_d_bits_data ;  
   wire _out_xbar_auto_in_d_bits_corrupt ;  
   wire _out_xbar_auto_out_4_a_valid ;  
   wire [2:0] _out_xbar_auto_out_4_a_bits_opcode ;  
   wire [2:0] _out_xbar_auto_out_4_a_bits_param ;  
   wire [2:0] _out_xbar_auto_out_4_a_bits_size ;  
   wire [4:0] _out_xbar_auto_out_4_a_bits_source ;  
   wire [16:0] _out_xbar_auto_out_4_a_bits_address ;  
   wire [7:0] _out_xbar_auto_out_4_a_bits_mask ;  
   wire _out_xbar_auto_out_4_a_bits_corrupt ;  
   wire _out_xbar_auto_out_4_d_ready ;  
   wire _out_xbar_auto_out_3_a_valid ;  
   wire [2:0] _out_xbar_auto_out_3_a_bits_opcode ;  
   wire [2:0] _out_xbar_auto_out_3_a_bits_param ;  
   wire [2:0] _out_xbar_auto_out_3_a_bits_size ;  
   wire [4:0] _out_xbar_auto_out_3_a_bits_source ;  
   wire [11:0] _out_xbar_auto_out_3_a_bits_address ;  
   wire [7:0] _out_xbar_auto_out_3_a_bits_mask ;  
   wire [63:0] _out_xbar_auto_out_3_a_bits_data ;  
   wire _out_xbar_auto_out_3_a_bits_corrupt ;  
   wire _out_xbar_auto_out_3_d_ready ;  
   wire _out_xbar_auto_out_2_a_valid ;  
   wire [2:0] _out_xbar_auto_out_2_a_bits_opcode ;  
   wire [2:0] _out_xbar_auto_out_2_a_bits_param ;  
   wire [2:0] _out_xbar_auto_out_2_a_bits_size ;  
   wire [4:0] _out_xbar_auto_out_2_a_bits_source ;  
   wire [25:0] _out_xbar_auto_out_2_a_bits_address ;  
   wire [7:0] _out_xbar_auto_out_2_a_bits_mask ;  
   wire [63:0] _out_xbar_auto_out_2_a_bits_data ;  
   wire _out_xbar_auto_out_2_a_bits_corrupt ;  
   wire _out_xbar_auto_out_2_d_ready ;  
   wire _out_xbar_auto_out_1_a_valid ;  
   wire [2:0] _out_xbar_auto_out_1_a_bits_opcode ;  
   wire [2:0] _out_xbar_auto_out_1_a_bits_param ;  
   wire [2:0] _out_xbar_auto_out_1_a_bits_size ;  
   wire [4:0] _out_xbar_auto_out_1_a_bits_source ;  
   wire [27:0] _out_xbar_auto_out_1_a_bits_address ;  
   wire [7:0] _out_xbar_auto_out_1_a_bits_mask ;  
   wire [63:0] _out_xbar_auto_out_1_a_bits_data ;  
   wire _out_xbar_auto_out_1_a_bits_corrupt ;  
   wire _out_xbar_auto_out_1_d_ready ;  
   wire _out_xbar_auto_out_0_a_valid ;  
   wire [2:0] _out_xbar_auto_out_0_a_bits_opcode ;  
   wire [2:0] _out_xbar_auto_out_0_a_bits_param ;  
   wire [3:0] _out_xbar_auto_out_0_a_bits_size ;  
   wire [4:0] _out_xbar_auto_out_0_a_bits_source ;  
   wire [13:0] _out_xbar_auto_out_0_a_bits_address ;  
   wire [7:0] _out_xbar_auto_out_0_a_bits_mask ;  
   wire _out_xbar_auto_out_0_a_bits_corrupt ;  
   wire _out_xbar_auto_out_0_d_ready ;  
   wire _fixer_auto_in_a_ready ;  
   wire _fixer_auto_in_d_valid ;  
   wire [2:0] _fixer_auto_in_d_bits_opcode ;  
   wire [1:0] _fixer_auto_in_d_bits_param ;  
   wire [3:0] _fixer_auto_in_d_bits_size ;  
   wire [4:0] _fixer_auto_in_d_bits_source ;  
   wire _fixer_auto_in_d_bits_sink ;  
   wire _fixer_auto_in_d_bits_denied ;  
   wire [63:0] _fixer_auto_in_d_bits_data ;  
   wire _fixer_auto_in_d_bits_corrupt ;  
   wire _fixer_auto_out_a_valid ;  
   wire [2:0] _fixer_auto_out_a_bits_opcode ;  
   wire [2:0] _fixer_auto_out_a_bits_param ;  
   wire [3:0] _fixer_auto_out_a_bits_size ;  
   wire [4:0] _fixer_auto_out_a_bits_source ;  
   wire [27:0] _fixer_auto_out_a_bits_address ;  
   wire [7:0] _fixer_auto_out_a_bits_mask ;  
   wire [63:0] _fixer_auto_out_a_bits_data ;  
   wire _fixer_auto_out_a_bits_corrupt ;  
   wire _fixer_auto_out_d_ready ;  
   wire _fixedClockNode_auto_out_0_clock ;  
   wire _fixedClockNode_auto_out_0_reset ;  
  FixedClockBroadcast_3 fixedClockNode(.auto_in_clock(auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock),.auto_in_reset(auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset),.auto_out_3_clock(auto_fixedClockNode_out_2_clock),.auto_out_3_reset(auto_fixedClockNode_out_2_reset),.auto_out_1_clock(auto_fixedClockNode_out_0_clock),.auto_out_1_reset(auto_fixedClockNode_out_0_reset),.auto_out_0_clock(_fixedClockNode_auto_out_0_clock),.auto_out_0_reset(_fixedClockNode_auto_out_0_reset)); 
  TLFIFOFixer_3 fixer(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_in_a_ready(_fixer_auto_in_a_ready),.auto_in_a_valid(_buffer_auto_out_a_valid),.auto_in_a_bits_opcode(_buffer_auto_out_a_bits_opcode),.auto_in_a_bits_param(_buffer_auto_out_a_bits_param),.auto_in_a_bits_size(_buffer_auto_out_a_bits_size),.auto_in_a_bits_source(_buffer_auto_out_a_bits_source),.auto_in_a_bits_address(_buffer_auto_out_a_bits_address),.auto_in_a_bits_mask(_buffer_auto_out_a_bits_mask),.auto_in_a_bits_data(_buffer_auto_out_a_bits_data),.auto_in_a_bits_corrupt(_buffer_auto_out_a_bits_corrupt),.auto_in_d_ready(_buffer_auto_out_d_ready),.auto_in_d_valid(_fixer_auto_in_d_valid),.auto_in_d_bits_opcode(_fixer_auto_in_d_bits_opcode),.auto_in_d_bits_param(_fixer_auto_in_d_bits_param),.auto_in_d_bits_size(_fixer_auto_in_d_bits_size),.auto_in_d_bits_source(_fixer_auto_in_d_bits_source),.auto_in_d_bits_sink(_fixer_auto_in_d_bits_sink),.auto_in_d_bits_denied(_fixer_auto_in_d_bits_denied),.auto_in_d_bits_data(_fixer_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_fixer_auto_in_d_bits_corrupt),.auto_out_a_ready(_out_xbar_auto_in_a_ready),.auto_out_a_valid(_fixer_auto_out_a_valid),.auto_out_a_bits_opcode(_fixer_auto_out_a_bits_opcode),.auto_out_a_bits_param(_fixer_auto_out_a_bits_param),.auto_out_a_bits_size(_fixer_auto_out_a_bits_size),.auto_out_a_bits_source(_fixer_auto_out_a_bits_source),.auto_out_a_bits_address(_fixer_auto_out_a_bits_address),.auto_out_a_bits_mask(_fixer_auto_out_a_bits_mask),.auto_out_a_bits_data(_fixer_auto_out_a_bits_data),.auto_out_a_bits_corrupt(_fixer_auto_out_a_bits_corrupt),.auto_out_d_ready(_fixer_auto_out_d_ready),.auto_out_d_valid(_out_xbar_auto_in_d_valid),.auto_out_d_bits_opcode(_out_xbar_auto_in_d_bits_opcode),.auto_out_d_bits_param(_out_xbar_auto_in_d_bits_param),.auto_out_d_bits_size(_out_xbar_auto_in_d_bits_size),.auto_out_d_bits_source(_out_xbar_auto_in_d_bits_source),.auto_out_d_bits_sink(_out_xbar_auto_in_d_bits_sink),.auto_out_d_bits_denied(_out_xbar_auto_in_d_bits_denied),.auto_out_d_bits_data(_out_xbar_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_out_xbar_auto_in_d_bits_corrupt)); 
  TLXbar_5 out_xbar(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_in_a_ready(_out_xbar_auto_in_a_ready),.auto_in_a_valid(_fixer_auto_out_a_valid),.auto_in_a_bits_opcode(_fixer_auto_out_a_bits_opcode),.auto_in_a_bits_param(_fixer_auto_out_a_bits_param),.auto_in_a_bits_size(_fixer_auto_out_a_bits_size),.auto_in_a_bits_source(_fixer_auto_out_a_bits_source),.auto_in_a_bits_address(_fixer_auto_out_a_bits_address),.auto_in_a_bits_mask(_fixer_auto_out_a_bits_mask),.auto_in_a_bits_data(_fixer_auto_out_a_bits_data),.auto_in_a_bits_corrupt(_fixer_auto_out_a_bits_corrupt),.auto_in_d_ready(_fixer_auto_out_d_ready),.auto_in_d_valid(_out_xbar_auto_in_d_valid),.auto_in_d_bits_opcode(_out_xbar_auto_in_d_bits_opcode),.auto_in_d_bits_param(_out_xbar_auto_in_d_bits_param),.auto_in_d_bits_size(_out_xbar_auto_in_d_bits_size),.auto_in_d_bits_source(_out_xbar_auto_in_d_bits_source),.auto_in_d_bits_sink(_out_xbar_auto_in_d_bits_sink),.auto_in_d_bits_denied(_out_xbar_auto_in_d_bits_denied),.auto_in_d_bits_data(_out_xbar_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_out_xbar_auto_in_d_bits_corrupt),.auto_out_4_a_ready(_coupler_to_bootrom_auto_tl_in_a_ready),.auto_out_4_a_valid(_out_xbar_auto_out_4_a_valid),.auto_out_4_a_bits_opcode(_out_xbar_auto_out_4_a_bits_opcode),.auto_out_4_a_bits_param(_out_xbar_auto_out_4_a_bits_param),.auto_out_4_a_bits_size(_out_xbar_auto_out_4_a_bits_size),.auto_out_4_a_bits_source(_out_xbar_auto_out_4_a_bits_source),.auto_out_4_a_bits_address(_out_xbar_auto_out_4_a_bits_address),.auto_out_4_a_bits_mask(_out_xbar_auto_out_4_a_bits_mask),.auto_out_4_a_bits_corrupt(_out_xbar_auto_out_4_a_bits_corrupt),.auto_out_4_d_ready(_out_xbar_auto_out_4_d_ready),.auto_out_4_d_valid(_coupler_to_bootrom_auto_tl_in_d_valid),.auto_out_4_d_bits_size(_coupler_to_bootrom_auto_tl_in_d_bits_size),.auto_out_4_d_bits_source(_coupler_to_bootrom_auto_tl_in_d_bits_source),.auto_out_4_d_bits_data(_coupler_to_bootrom_auto_tl_in_d_bits_data),.auto_out_3_a_ready(_coupler_to_debug_auto_tl_in_a_ready),.auto_out_3_a_valid(_out_xbar_auto_out_3_a_valid),.auto_out_3_a_bits_opcode(_out_xbar_auto_out_3_a_bits_opcode),.auto_out_3_a_bits_param(_out_xbar_auto_out_3_a_bits_param),.auto_out_3_a_bits_size(_out_xbar_auto_out_3_a_bits_size),.auto_out_3_a_bits_source(_out_xbar_auto_out_3_a_bits_source),.auto_out_3_a_bits_address(_out_xbar_auto_out_3_a_bits_address),.auto_out_3_a_bits_mask(_out_xbar_auto_out_3_a_bits_mask),.auto_out_3_a_bits_data(_out_xbar_auto_out_3_a_bits_data),.auto_out_3_a_bits_corrupt(_out_xbar_auto_out_3_a_bits_corrupt),.auto_out_3_d_ready(_out_xbar_auto_out_3_d_ready),.auto_out_3_d_valid(_coupler_to_debug_auto_tl_in_d_valid),.auto_out_3_d_bits_opcode(_coupler_to_debug_auto_tl_in_d_bits_opcode),.auto_out_3_d_bits_size(_coupler_to_debug_auto_tl_in_d_bits_size),.auto_out_3_d_bits_source(_coupler_to_debug_auto_tl_in_d_bits_source),.auto_out_3_d_bits_data(_coupler_to_debug_auto_tl_in_d_bits_data),.auto_out_2_a_ready(_coupler_to_clint_auto_tl_in_a_ready),.auto_out_2_a_valid(_out_xbar_auto_out_2_a_valid),.auto_out_2_a_bits_opcode(_out_xbar_auto_out_2_a_bits_opcode),.auto_out_2_a_bits_param(_out_xbar_auto_out_2_a_bits_param),.auto_out_2_a_bits_size(_out_xbar_auto_out_2_a_bits_size),.auto_out_2_a_bits_source(_out_xbar_auto_out_2_a_bits_source),.auto_out_2_a_bits_address(_out_xbar_auto_out_2_a_bits_address),.auto_out_2_a_bits_mask(_out_xbar_auto_out_2_a_bits_mask),.auto_out_2_a_bits_data(_out_xbar_auto_out_2_a_bits_data),.auto_out_2_a_bits_corrupt(_out_xbar_auto_out_2_a_bits_corrupt),.auto_out_2_d_ready(_out_xbar_auto_out_2_d_ready),.auto_out_2_d_valid(_coupler_to_clint_auto_tl_in_d_valid),.auto_out_2_d_bits_opcode(_coupler_to_clint_auto_tl_in_d_bits_opcode),.auto_out_2_d_bits_size(_coupler_to_clint_auto_tl_in_d_bits_size),.auto_out_2_d_bits_source(_coupler_to_clint_auto_tl_in_d_bits_source),.auto_out_2_d_bits_data(_coupler_to_clint_auto_tl_in_d_bits_data),.auto_out_1_a_ready(_coupler_to_plic_auto_tl_in_a_ready),.auto_out_1_a_valid(_out_xbar_auto_out_1_a_valid),.auto_out_1_a_bits_opcode(_out_xbar_auto_out_1_a_bits_opcode),.auto_out_1_a_bits_param(_out_xbar_auto_out_1_a_bits_param),.auto_out_1_a_bits_size(_out_xbar_auto_out_1_a_bits_size),.auto_out_1_a_bits_source(_out_xbar_auto_out_1_a_bits_source),.auto_out_1_a_bits_address(_out_xbar_auto_out_1_a_bits_address),.auto_out_1_a_bits_mask(_out_xbar_auto_out_1_a_bits_mask),.auto_out_1_a_bits_data(_out_xbar_auto_out_1_a_bits_data),.auto_out_1_a_bits_corrupt(_out_xbar_auto_out_1_a_bits_corrupt),.auto_out_1_d_ready(_out_xbar_auto_out_1_d_ready),.auto_out_1_d_valid(_coupler_to_plic_auto_tl_in_d_valid),.auto_out_1_d_bits_opcode(_coupler_to_plic_auto_tl_in_d_bits_opcode),.auto_out_1_d_bits_size(_coupler_to_plic_auto_tl_in_d_bits_size),.auto_out_1_d_bits_source(_coupler_to_plic_auto_tl_in_d_bits_source),.auto_out_1_d_bits_data(_coupler_to_plic_auto_tl_in_d_bits_data),.auto_out_0_a_ready(_wrapped_error_device_auto_buffer_in_a_ready),.auto_out_0_a_valid(_out_xbar_auto_out_0_a_valid),.auto_out_0_a_bits_opcode(_out_xbar_auto_out_0_a_bits_opcode),.auto_out_0_a_bits_param(_out_xbar_auto_out_0_a_bits_param),.auto_out_0_a_bits_size(_out_xbar_auto_out_0_a_bits_size),.auto_out_0_a_bits_source(_out_xbar_auto_out_0_a_bits_source),.auto_out_0_a_bits_address(_out_xbar_auto_out_0_a_bits_address),.auto_out_0_a_bits_mask(_out_xbar_auto_out_0_a_bits_mask),.auto_out_0_a_bits_corrupt(_out_xbar_auto_out_0_a_bits_corrupt),.auto_out_0_d_ready(_out_xbar_auto_out_0_d_ready),.auto_out_0_d_valid(_wrapped_error_device_auto_buffer_in_d_valid),.auto_out_0_d_bits_opcode(_wrapped_error_device_auto_buffer_in_d_bits_opcode),.auto_out_0_d_bits_param(_wrapped_error_device_auto_buffer_in_d_bits_param),.auto_out_0_d_bits_size(_wrapped_error_device_auto_buffer_in_d_bits_size),.auto_out_0_d_bits_source(_wrapped_error_device_auto_buffer_in_d_bits_source),.auto_out_0_d_bits_sink(_wrapped_error_device_auto_buffer_in_d_bits_sink),.auto_out_0_d_bits_denied(_wrapped_error_device_auto_buffer_in_d_bits_denied),.auto_out_0_d_bits_data(_wrapped_error_device_auto_buffer_in_d_bits_data),.auto_out_0_d_bits_corrupt(_wrapped_error_device_auto_buffer_in_d_bits_corrupt)); 
  TLBuffer_4 buffer(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_in_a_ready(_buffer_auto_in_a_ready),.auto_in_a_valid(_atomics_auto_out_a_valid),.auto_in_a_bits_opcode(_atomics_auto_out_a_bits_opcode),.auto_in_a_bits_param(_atomics_auto_out_a_bits_param),.auto_in_a_bits_size(_atomics_auto_out_a_bits_size),.auto_in_a_bits_source(_atomics_auto_out_a_bits_source),.auto_in_a_bits_address(_atomics_auto_out_a_bits_address),.auto_in_a_bits_mask(_atomics_auto_out_a_bits_mask),.auto_in_a_bits_data(_atomics_auto_out_a_bits_data),.auto_in_a_bits_corrupt(_atomics_auto_out_a_bits_corrupt),.auto_in_d_ready(_atomics_auto_out_d_ready),.auto_in_d_valid(_buffer_auto_in_d_valid),.auto_in_d_bits_opcode(_buffer_auto_in_d_bits_opcode),.auto_in_d_bits_param(_buffer_auto_in_d_bits_param),.auto_in_d_bits_size(_buffer_auto_in_d_bits_size),.auto_in_d_bits_source(_buffer_auto_in_d_bits_source),.auto_in_d_bits_sink(_buffer_auto_in_d_bits_sink),.auto_in_d_bits_denied(_buffer_auto_in_d_bits_denied),.auto_in_d_bits_data(_buffer_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt),.auto_out_a_ready(_fixer_auto_in_a_ready),.auto_out_a_valid(_buffer_auto_out_a_valid),.auto_out_a_bits_opcode(_buffer_auto_out_a_bits_opcode),.auto_out_a_bits_param(_buffer_auto_out_a_bits_param),.auto_out_a_bits_size(_buffer_auto_out_a_bits_size),.auto_out_a_bits_source(_buffer_auto_out_a_bits_source),.auto_out_a_bits_address(_buffer_auto_out_a_bits_address),.auto_out_a_bits_mask(_buffer_auto_out_a_bits_mask),.auto_out_a_bits_data(_buffer_auto_out_a_bits_data),.auto_out_a_bits_corrupt(_buffer_auto_out_a_bits_corrupt),.auto_out_d_ready(_buffer_auto_out_d_ready),.auto_out_d_valid(_fixer_auto_in_d_valid),.auto_out_d_bits_opcode(_fixer_auto_in_d_bits_opcode),.auto_out_d_bits_param(_fixer_auto_in_d_bits_param),.auto_out_d_bits_size(_fixer_auto_in_d_bits_size),.auto_out_d_bits_source(_fixer_auto_in_d_bits_source),.auto_out_d_bits_sink(_fixer_auto_in_d_bits_sink),.auto_out_d_bits_denied(_fixer_auto_in_d_bits_denied),.auto_out_d_bits_data(_fixer_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_fixer_auto_in_d_bits_corrupt)); 
  TLAtomicAutomata_1 atomics(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_in_a_ready(auto_bus_xing_in_a_ready),.auto_in_a_valid(auto_bus_xing_in_a_valid),.auto_in_a_bits_opcode(auto_bus_xing_in_a_bits_opcode),.auto_in_a_bits_param(auto_bus_xing_in_a_bits_param),.auto_in_a_bits_size(auto_bus_xing_in_a_bits_size),.auto_in_a_bits_source(auto_bus_xing_in_a_bits_source),.auto_in_a_bits_address(auto_bus_xing_in_a_bits_address),.auto_in_a_bits_mask(auto_bus_xing_in_a_bits_mask),.auto_in_a_bits_data(auto_bus_xing_in_a_bits_data),.auto_in_a_bits_corrupt(auto_bus_xing_in_a_bits_corrupt),.auto_in_d_ready(auto_bus_xing_in_d_ready),.auto_in_d_valid(auto_bus_xing_in_d_valid),.auto_in_d_bits_opcode(auto_bus_xing_in_d_bits_opcode),.auto_in_d_bits_param(auto_bus_xing_in_d_bits_param),.auto_in_d_bits_size(auto_bus_xing_in_d_bits_size),.auto_in_d_bits_source(auto_bus_xing_in_d_bits_source),.auto_in_d_bits_sink(auto_bus_xing_in_d_bits_sink),.auto_in_d_bits_denied(auto_bus_xing_in_d_bits_denied),.auto_in_d_bits_data(auto_bus_xing_in_d_bits_data),.auto_in_d_bits_corrupt(auto_bus_xing_in_d_bits_corrupt),.auto_out_a_ready(_buffer_auto_in_a_ready),.auto_out_a_valid(_atomics_auto_out_a_valid),.auto_out_a_bits_opcode(_atomics_auto_out_a_bits_opcode),.auto_out_a_bits_param(_atomics_auto_out_a_bits_param),.auto_out_a_bits_size(_atomics_auto_out_a_bits_size),.auto_out_a_bits_source(_atomics_auto_out_a_bits_source),.auto_out_a_bits_address(_atomics_auto_out_a_bits_address),.auto_out_a_bits_mask(_atomics_auto_out_a_bits_mask),.auto_out_a_bits_data(_atomics_auto_out_a_bits_data),.auto_out_a_bits_corrupt(_atomics_auto_out_a_bits_corrupt),.auto_out_d_ready(_atomics_auto_out_d_ready),.auto_out_d_valid(_buffer_auto_in_d_valid),.auto_out_d_bits_opcode(_buffer_auto_in_d_bits_opcode),.auto_out_d_bits_param(_buffer_auto_in_d_bits_param),.auto_out_d_bits_size(_buffer_auto_in_d_bits_size),.auto_out_d_bits_source(_buffer_auto_in_d_bits_source),.auto_out_d_bits_sink(_buffer_auto_in_d_bits_sink),.auto_out_d_bits_denied(_buffer_auto_in_d_bits_denied),.auto_out_d_bits_data(_buffer_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt)); 
  ErrorDeviceWrapper wrapped_error_device(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_buffer_in_a_ready(_wrapped_error_device_auto_buffer_in_a_ready),.auto_buffer_in_a_valid(_out_xbar_auto_out_0_a_valid),.auto_buffer_in_a_bits_opcode(_out_xbar_auto_out_0_a_bits_opcode),.auto_buffer_in_a_bits_param(_out_xbar_auto_out_0_a_bits_param),.auto_buffer_in_a_bits_size(_out_xbar_auto_out_0_a_bits_size),.auto_buffer_in_a_bits_source(_out_xbar_auto_out_0_a_bits_source),.auto_buffer_in_a_bits_address(_out_xbar_auto_out_0_a_bits_address),.auto_buffer_in_a_bits_mask(_out_xbar_auto_out_0_a_bits_mask),.auto_buffer_in_a_bits_corrupt(_out_xbar_auto_out_0_a_bits_corrupt),.auto_buffer_in_d_ready(_out_xbar_auto_out_0_d_ready),.auto_buffer_in_d_valid(_wrapped_error_device_auto_buffer_in_d_valid),.auto_buffer_in_d_bits_opcode(_wrapped_error_device_auto_buffer_in_d_bits_opcode),.auto_buffer_in_d_bits_param(_wrapped_error_device_auto_buffer_in_d_bits_param),.auto_buffer_in_d_bits_size(_wrapped_error_device_auto_buffer_in_d_bits_size),.auto_buffer_in_d_bits_source(_wrapped_error_device_auto_buffer_in_d_bits_source),.auto_buffer_in_d_bits_sink(_wrapped_error_device_auto_buffer_in_d_bits_sink),.auto_buffer_in_d_bits_denied(_wrapped_error_device_auto_buffer_in_d_bits_denied),.auto_buffer_in_d_bits_data(_wrapped_error_device_auto_buffer_in_d_bits_data),.auto_buffer_in_d_bits_corrupt(_wrapped_error_device_auto_buffer_in_d_bits_corrupt)); 
  TLInterconnectCoupler_7 coupler_to_plic(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_fragmenter_out_a_ready(auto_coupler_to_plic_fragmenter_out_a_ready),.auto_fragmenter_out_a_valid(auto_coupler_to_plic_fragmenter_out_a_valid),.auto_fragmenter_out_a_bits_opcode(auto_coupler_to_plic_fragmenter_out_a_bits_opcode),.auto_fragmenter_out_a_bits_param(auto_coupler_to_plic_fragmenter_out_a_bits_param),.auto_fragmenter_out_a_bits_size(auto_coupler_to_plic_fragmenter_out_a_bits_size),.auto_fragmenter_out_a_bits_source(auto_coupler_to_plic_fragmenter_out_a_bits_source),.auto_fragmenter_out_a_bits_address(auto_coupler_to_plic_fragmenter_out_a_bits_address),.auto_fragmenter_out_a_bits_mask(auto_coupler_to_plic_fragmenter_out_a_bits_mask),.auto_fragmenter_out_a_bits_data(auto_coupler_to_plic_fragmenter_out_a_bits_data),.auto_fragmenter_out_a_bits_corrupt(auto_coupler_to_plic_fragmenter_out_a_bits_corrupt),.auto_fragmenter_out_d_ready(auto_coupler_to_plic_fragmenter_out_d_ready),.auto_fragmenter_out_d_valid(auto_coupler_to_plic_fragmenter_out_d_valid),.auto_fragmenter_out_d_bits_opcode(auto_coupler_to_plic_fragmenter_out_d_bits_opcode),.auto_fragmenter_out_d_bits_size(auto_coupler_to_plic_fragmenter_out_d_bits_size),.auto_fragmenter_out_d_bits_source(auto_coupler_to_plic_fragmenter_out_d_bits_source),.auto_fragmenter_out_d_bits_data(auto_coupler_to_plic_fragmenter_out_d_bits_data),.auto_tl_in_a_ready(_coupler_to_plic_auto_tl_in_a_ready),.auto_tl_in_a_valid(_out_xbar_auto_out_1_a_valid),.auto_tl_in_a_bits_opcode(_out_xbar_auto_out_1_a_bits_opcode),.auto_tl_in_a_bits_param(_out_xbar_auto_out_1_a_bits_param),.auto_tl_in_a_bits_size(_out_xbar_auto_out_1_a_bits_size),.auto_tl_in_a_bits_source(_out_xbar_auto_out_1_a_bits_source),.auto_tl_in_a_bits_address(_out_xbar_auto_out_1_a_bits_address),.auto_tl_in_a_bits_mask(_out_xbar_auto_out_1_a_bits_mask),.auto_tl_in_a_bits_data(_out_xbar_auto_out_1_a_bits_data),.auto_tl_in_a_bits_corrupt(_out_xbar_auto_out_1_a_bits_corrupt),.auto_tl_in_d_ready(_out_xbar_auto_out_1_d_ready),.auto_tl_in_d_valid(_coupler_to_plic_auto_tl_in_d_valid),.auto_tl_in_d_bits_opcode(_coupler_to_plic_auto_tl_in_d_bits_opcode),.auto_tl_in_d_bits_size(_coupler_to_plic_auto_tl_in_d_bits_size),.auto_tl_in_d_bits_source(_coupler_to_plic_auto_tl_in_d_bits_source),.auto_tl_in_d_bits_data(_coupler_to_plic_auto_tl_in_d_bits_data)); 
  TLInterconnectCoupler_8 coupler_to_clint(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_fragmenter_out_a_ready(auto_coupler_to_clint_fragmenter_out_a_ready),.auto_fragmenter_out_a_valid(auto_coupler_to_clint_fragmenter_out_a_valid),.auto_fragmenter_out_a_bits_opcode(auto_coupler_to_clint_fragmenter_out_a_bits_opcode),.auto_fragmenter_out_a_bits_param(auto_coupler_to_clint_fragmenter_out_a_bits_param),.auto_fragmenter_out_a_bits_size(auto_coupler_to_clint_fragmenter_out_a_bits_size),.auto_fragmenter_out_a_bits_source(auto_coupler_to_clint_fragmenter_out_a_bits_source),.auto_fragmenter_out_a_bits_address(auto_coupler_to_clint_fragmenter_out_a_bits_address),.auto_fragmenter_out_a_bits_mask(auto_coupler_to_clint_fragmenter_out_a_bits_mask),.auto_fragmenter_out_a_bits_data(auto_coupler_to_clint_fragmenter_out_a_bits_data),.auto_fragmenter_out_a_bits_corrupt(auto_coupler_to_clint_fragmenter_out_a_bits_corrupt),.auto_fragmenter_out_d_ready(auto_coupler_to_clint_fragmenter_out_d_ready),.auto_fragmenter_out_d_valid(auto_coupler_to_clint_fragmenter_out_d_valid),.auto_fragmenter_out_d_bits_opcode(auto_coupler_to_clint_fragmenter_out_d_bits_opcode),.auto_fragmenter_out_d_bits_size(auto_coupler_to_clint_fragmenter_out_d_bits_size),.auto_fragmenter_out_d_bits_source(auto_coupler_to_clint_fragmenter_out_d_bits_source),.auto_fragmenter_out_d_bits_data(auto_coupler_to_clint_fragmenter_out_d_bits_data),.auto_tl_in_a_ready(_coupler_to_clint_auto_tl_in_a_ready),.auto_tl_in_a_valid(_out_xbar_auto_out_2_a_valid),.auto_tl_in_a_bits_opcode(_out_xbar_auto_out_2_a_bits_opcode),.auto_tl_in_a_bits_param(_out_xbar_auto_out_2_a_bits_param),.auto_tl_in_a_bits_size(_out_xbar_auto_out_2_a_bits_size),.auto_tl_in_a_bits_source(_out_xbar_auto_out_2_a_bits_source),.auto_tl_in_a_bits_address(_out_xbar_auto_out_2_a_bits_address),.auto_tl_in_a_bits_mask(_out_xbar_auto_out_2_a_bits_mask),.auto_tl_in_a_bits_data(_out_xbar_auto_out_2_a_bits_data),.auto_tl_in_a_bits_corrupt(_out_xbar_auto_out_2_a_bits_corrupt),.auto_tl_in_d_ready(_out_xbar_auto_out_2_d_ready),.auto_tl_in_d_valid(_coupler_to_clint_auto_tl_in_d_valid),.auto_tl_in_d_bits_opcode(_coupler_to_clint_auto_tl_in_d_bits_opcode),.auto_tl_in_d_bits_size(_coupler_to_clint_auto_tl_in_d_bits_size),.auto_tl_in_d_bits_source(_coupler_to_clint_auto_tl_in_d_bits_source),.auto_tl_in_d_bits_data(_coupler_to_clint_auto_tl_in_d_bits_data)); 
  TLInterconnectCoupler_10 coupler_to_debug(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_fragmenter_out_a_ready(auto_coupler_to_debug_fragmenter_out_a_ready),.auto_fragmenter_out_a_valid(auto_coupler_to_debug_fragmenter_out_a_valid),.auto_fragmenter_out_a_bits_opcode(auto_coupler_to_debug_fragmenter_out_a_bits_opcode),.auto_fragmenter_out_a_bits_param(auto_coupler_to_debug_fragmenter_out_a_bits_param),.auto_fragmenter_out_a_bits_size(auto_coupler_to_debug_fragmenter_out_a_bits_size),.auto_fragmenter_out_a_bits_source(auto_coupler_to_debug_fragmenter_out_a_bits_source),.auto_fragmenter_out_a_bits_address(auto_coupler_to_debug_fragmenter_out_a_bits_address),.auto_fragmenter_out_a_bits_mask(auto_coupler_to_debug_fragmenter_out_a_bits_mask),.auto_fragmenter_out_a_bits_data(auto_coupler_to_debug_fragmenter_out_a_bits_data),.auto_fragmenter_out_a_bits_corrupt(auto_coupler_to_debug_fragmenter_out_a_bits_corrupt),.auto_fragmenter_out_d_ready(auto_coupler_to_debug_fragmenter_out_d_ready),.auto_fragmenter_out_d_valid(auto_coupler_to_debug_fragmenter_out_d_valid),.auto_fragmenter_out_d_bits_opcode(auto_coupler_to_debug_fragmenter_out_d_bits_opcode),.auto_fragmenter_out_d_bits_size(auto_coupler_to_debug_fragmenter_out_d_bits_size),.auto_fragmenter_out_d_bits_source(auto_coupler_to_debug_fragmenter_out_d_bits_source),.auto_fragmenter_out_d_bits_data(auto_coupler_to_debug_fragmenter_out_d_bits_data),.auto_tl_in_a_ready(_coupler_to_debug_auto_tl_in_a_ready),.auto_tl_in_a_valid(_out_xbar_auto_out_3_a_valid),.auto_tl_in_a_bits_opcode(_out_xbar_auto_out_3_a_bits_opcode),.auto_tl_in_a_bits_param(_out_xbar_auto_out_3_a_bits_param),.auto_tl_in_a_bits_size(_out_xbar_auto_out_3_a_bits_size),.auto_tl_in_a_bits_source(_out_xbar_auto_out_3_a_bits_source),.auto_tl_in_a_bits_address(_out_xbar_auto_out_3_a_bits_address),.auto_tl_in_a_bits_mask(_out_xbar_auto_out_3_a_bits_mask),.auto_tl_in_a_bits_data(_out_xbar_auto_out_3_a_bits_data),.auto_tl_in_a_bits_corrupt(_out_xbar_auto_out_3_a_bits_corrupt),.auto_tl_in_d_ready(_out_xbar_auto_out_3_d_ready),.auto_tl_in_d_valid(_coupler_to_debug_auto_tl_in_d_valid),.auto_tl_in_d_bits_opcode(_coupler_to_debug_auto_tl_in_d_bits_opcode),.auto_tl_in_d_bits_size(_coupler_to_debug_auto_tl_in_d_bits_size),.auto_tl_in_d_bits_source(_coupler_to_debug_auto_tl_in_d_bits_source),.auto_tl_in_d_bits_data(_coupler_to_debug_auto_tl_in_d_bits_data)); 
  TLInterconnectCoupler_11 coupler_to_bootrom(.clock(_fixedClockNode_auto_out_0_clock),.reset(_fixedClockNode_auto_out_0_reset),.auto_fragmenter_out_a_ready(auto_coupler_to_bootrom_fragmenter_out_a_ready),.auto_fragmenter_out_a_valid(auto_coupler_to_bootrom_fragmenter_out_a_valid),.auto_fragmenter_out_a_bits_opcode(auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode),.auto_fragmenter_out_a_bits_param(auto_coupler_to_bootrom_fragmenter_out_a_bits_param),.auto_fragmenter_out_a_bits_size(auto_coupler_to_bootrom_fragmenter_out_a_bits_size),.auto_fragmenter_out_a_bits_source(auto_coupler_to_bootrom_fragmenter_out_a_bits_source),.auto_fragmenter_out_a_bits_address(auto_coupler_to_bootrom_fragmenter_out_a_bits_address),.auto_fragmenter_out_a_bits_mask(auto_coupler_to_bootrom_fragmenter_out_a_bits_mask),.auto_fragmenter_out_a_bits_corrupt(auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt),.auto_fragmenter_out_d_ready(auto_coupler_to_bootrom_fragmenter_out_d_ready),.auto_fragmenter_out_d_valid(auto_coupler_to_bootrom_fragmenter_out_d_valid),.auto_fragmenter_out_d_bits_size(auto_coupler_to_bootrom_fragmenter_out_d_bits_size),.auto_fragmenter_out_d_bits_source(auto_coupler_to_bootrom_fragmenter_out_d_bits_source),.auto_fragmenter_out_d_bits_data(auto_coupler_to_bootrom_fragmenter_out_d_bits_data),.auto_tl_in_a_ready(_coupler_to_bootrom_auto_tl_in_a_ready),.auto_tl_in_a_valid(_out_xbar_auto_out_4_a_valid),.auto_tl_in_a_bits_opcode(_out_xbar_auto_out_4_a_bits_opcode),.auto_tl_in_a_bits_param(_out_xbar_auto_out_4_a_bits_param),.auto_tl_in_a_bits_size(_out_xbar_auto_out_4_a_bits_size),.auto_tl_in_a_bits_source(_out_xbar_auto_out_4_a_bits_source),.auto_tl_in_a_bits_address(_out_xbar_auto_out_4_a_bits_address),.auto_tl_in_a_bits_mask(_out_xbar_auto_out_4_a_bits_mask),.auto_tl_in_a_bits_corrupt(_out_xbar_auto_out_4_a_bits_corrupt),.auto_tl_in_d_ready(_out_xbar_auto_out_4_d_ready),.auto_tl_in_d_valid(_coupler_to_bootrom_auto_tl_in_d_valid),.auto_tl_in_d_bits_size(_coupler_to_bootrom_auto_tl_in_d_bits_size),.auto_tl_in_d_bits_source(_coupler_to_bootrom_auto_tl_in_d_bits_source),.auto_tl_in_d_bits_data(_coupler_to_bootrom_auto_tl_in_d_bits_data)); 
  assign auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock=auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock; 
  assign auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset=auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset; 
  assign clock=_fixedClockNode_auto_out_0_clock; 
  assign reset=_fixedClockNode_auto_out_0_reset; 
endmodule
 
module TLMonitor_18 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [6:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [2:0] io_in_d_bits_size,
  input [6:0] io_in_d_bits_source,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [6:0] source ;  
   reg [31:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [2:0] size_1 ;  
   reg [6:0] source_1 ;  
   reg denied ;  
   reg [127:0] inflight ;  
   reg [511:0] inflight_opcodes ;  
   reg [511:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [511:0] _GEN_0={503'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_0 ;  
   wire [127:0] _GEN_1={121'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [127:0] _GEN_3={121'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [127:0] inflight_1 ;  
   reg [511:0] inflight_sizes_1 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_4=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_a_bits_param>3'h2 ;  
   wire _GEN_7=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_8=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_9=io_in_a_bits_size!=3'h7&io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_11=io_in_a_bits_mask!=mask ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_18=io_in_d_bits_size<3'h3 ;  
   wire _GEN_19=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_20=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_21=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_22=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_23=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [127:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 128'h1<<_GEN_1:128'h0 ;  
   wire _GEN_24=io_in_d_valid&d_first_1 ;  
   wire _GEN_25=_GEN_24&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_26=_GEN_25&same_cycle_resp&~reset ;  
   wire _GEN_27=_GEN_25&~same_cycle_resp&~reset ;  
   wire _GEN_28=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [127:0] _GEN_29=inflight>>_GEN_1 ;  
   wire [127:0] _GEN_30=inflight>>_GEN_3 ;  
   wire [511:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_0 ;  
   wire [127:0] _GEN_31=inflight_1>>_GEN_3 ;  
   wire [511:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_0 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_29[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~reset&~(_GEN_30[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_25 ? 128'h1<<_GEN_3:128'h0)|a_set_wo_ready==128'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==128'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(_GEN_31[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==128'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/tilelink/CrossingHelper.scala:30:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_32={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_32 ;  
   wire [1026:0] _GEN_33={1018'h0,io_in_a_bits_source,2'h0} ;  
   wire [1038:0] _GEN_34={1030'h0,io_in_d_bits_source,2'h0} ;  
   wire [1038:0] _d_opcodes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_opcodes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_sizes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_11=1039'hF<<_GEN_34 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_35=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_36=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=128'h0;
              inflight_opcodes <=512'h0;
              inflight_sizes <=512'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=128'h0;
              inflight_sizes_1 <=512'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_2 ? 128'h1<<_GEN_1:128'h0))&~(_GEN_35 ? 128'h1<<_GEN_3:128'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_opcodes_clr_T_5[511:0]:512'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_sizes_clr_T_5[511:0]:512'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_36 ? 128'h1<<_GEN_3:128'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_36 ? _d_sizes_clr_T_11[511:0]:512'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLFIFOFixer_4 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [6:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [2:0] auto_in_d_bits_size,
  output [6:0] auto_in_d_bits_source,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [2:0] auto_out_a_bits_size,
  output [6:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [2:0] auto_out_d_bits_size,
  input [6:0] auto_out_d_bits_source,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
  TLMonitor_18 monitor(.clock(clock),.reset(reset),.io_in_a_ready(auto_out_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_out_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source),.io_in_d_bits_denied(auto_out_d_bits_denied),.io_in_d_bits_corrupt(auto_out_d_bits_corrupt)); 
  assign auto_in_a_ready=auto_out_a_ready; 
  assign auto_in_d_valid=auto_out_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source; 
  assign auto_in_d_bits_denied=auto_out_d_bits_denied; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign auto_out_a_valid=auto_in_a_valid; 
  assign auto_out_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_a_bits_size=auto_in_a_bits_size; 
  assign auto_out_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_d_ready=auto_in_d_ready; 
endmodule
 
module TLMonitor_19 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [6:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [2:0] io_in_d_bits_size,
  input [6:0] io_in_d_bits_source,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [6:0] source ;  
   reg [31:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [2:0] size_1 ;  
   reg [6:0] source_1 ;  
   reg denied ;  
   reg [127:0] inflight ;  
   reg [511:0] inflight_opcodes ;  
   reg [511:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [511:0] _GEN_0={503'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_0 ;  
   wire [127:0] _GEN_1={121'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [127:0] _GEN_3={121'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [127:0] inflight_1 ;  
   reg [511:0] inflight_sizes_1 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_4=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_a_bits_param>3'h2 ;  
   wire _GEN_7=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_8=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_9=io_in_a_bits_size!=3'h7&io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_11=io_in_a_bits_mask!=mask ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_18=io_in_d_bits_size<3'h3 ;  
   wire _GEN_19=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_20=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_21=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_22=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_23=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [127:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 128'h1<<_GEN_1:128'h0 ;  
   wire _GEN_24=io_in_d_valid&d_first_1 ;  
   wire _GEN_25=_GEN_24&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_26=_GEN_25&same_cycle_resp&~reset ;  
   wire _GEN_27=_GEN_25&~same_cycle_resp&~reset ;  
   wire _GEN_28=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [127:0] _GEN_29=inflight>>_GEN_1 ;  
   wire [127:0] _GEN_30=inflight>>_GEN_3 ;  
   wire [511:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_0 ;  
   wire [127:0] _GEN_31=inflight_1>>_GEN_3 ;  
   wire [511:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_0 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_29[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~reset&~(_GEN_30[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_25 ? 128'h1<<_GEN_3:128'h0)|a_set_wo_ready==128'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==128'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(_GEN_31[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==128'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/MemoryBus.scala:47:50)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_32={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_32 ;  
   wire [1026:0] _GEN_33={1018'h0,io_in_a_bits_source,2'h0} ;  
   wire [1038:0] _GEN_34={1030'h0,io_in_d_bits_source,2'h0} ;  
   wire [1038:0] _d_opcodes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_opcodes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_sizes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_11=1039'hF<<_GEN_34 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_35=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_36=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=128'h0;
              inflight_opcodes <=512'h0;
              inflight_sizes <=512'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=128'h0;
              inflight_sizes_1 <=512'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_2 ? 128'h1<<_GEN_1:128'h0))&~(_GEN_35 ? 128'h1<<_GEN_3:128'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_opcodes_clr_T_5[511:0]:512'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_sizes_clr_T_5[511:0]:512'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_36 ? 128'h1<<_GEN_3:128'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_36 ? _d_sizes_clr_T_11[511:0]:512'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module ProbePicker (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [6:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [2:0] auto_in_d_bits_size,
  output [6:0] auto_in_d_bits_source,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [2:0] auto_out_a_bits_size,
  output [6:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [2:0] auto_out_d_bits_size,
  input [6:0] auto_out_d_bits_source,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
  TLMonitor_19 monitor(.clock(clock),.reset(reset),.io_in_a_ready(auto_out_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_out_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source),.io_in_d_bits_denied(auto_out_d_bits_denied),.io_in_d_bits_corrupt(auto_out_d_bits_corrupt)); 
  assign auto_in_a_ready=auto_out_a_ready; 
  assign auto_in_d_valid=auto_out_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source; 
  assign auto_in_d_bits_denied=auto_out_d_bits_denied; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign auto_out_a_valid=auto_in_a_valid; 
  assign auto_out_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_a_bits_size=auto_in_a_bits_size; 
  assign auto_out_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_d_ready=auto_in_d_ready; 
endmodule
 
module ram_8x14 (
  input [2:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [13:0] R0_data,
  input [2:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [13:0] W0_data) ; 
   reg [13:0] Memory[0:7] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:14'bx; 
endmodule
 
module Queue_40 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_tl_state_size,
  input [6:0] io_enq_bits_tl_state_source,
  input [2:0] io_enq_bits_extra_id,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_tl_state_size,
  output [6:0] io_deq_bits_tl_state_source,
  output [2:0] io_deq_bits_extra_id) ; 
   wire [13:0] _ram_ext_R0_data ;  
   reg [2:0] enq_ptr_value ;  
   reg [2:0] deq_ptr_value ;  
   reg maybe_full ;  
   wire ptr_match=enq_ptr_value==deq_ptr_value ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              enq_ptr_value <=3'h0;
              deq_ptr_value <=3'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 enq_ptr_value <=enq_ptr_value+3'h1;
              if (do_deq)
                 deq_ptr_value <=deq_ptr_value+3'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_8x14 ram_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(_ram_ext_R0_data),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data({io_enq_bits_extra_id,io_enq_bits_tl_state_source,io_enq_bits_tl_state_size})); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
  assign io_deq_bits_tl_state_size=_ram_ext_R0_data[3:0]; 
  assign io_deq_bits_tl_state_source=_ram_ext_R0_data[10:4]; 
  assign io_deq_bits_extra_id=_ram_ext_R0_data[13:11]; 
endmodule
 
module AXI4UserYanker_2 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [3:0] auto_in_aw_bits_echo_tl_state_size,
  input [6:0] auto_in_aw_bits_echo_tl_state_source,
  input [2:0] auto_in_aw_bits_echo_extra_id,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output [3:0] auto_in_b_bits_echo_tl_state_size,
  output [6:0] auto_in_b_bits_echo_tl_state_source,
  output [2:0] auto_in_b_bits_echo_extra_id,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [3:0] auto_in_ar_bits_echo_tl_state_size,
  input [6:0] auto_in_ar_bits_echo_tl_state_source,
  input [2:0] auto_in_ar_bits_echo_extra_id,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output [3:0] auto_in_r_bits_echo_tl_state_size,
  output [6:0] auto_in_r_bits_echo_tl_state_source,
  output [2:0] auto_in_r_bits_echo_extra_id,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_last) ; 
   wire _Queue_31_io_enq_ready ;  
   wire _Queue_31_io_deq_valid ;  
   wire [3:0] _Queue_31_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_31_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_31_io_deq_bits_extra_id ;  
   wire _Queue_30_io_enq_ready ;  
   wire _Queue_30_io_deq_valid ;  
   wire [3:0] _Queue_30_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_30_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_30_io_deq_bits_extra_id ;  
   wire _Queue_29_io_enq_ready ;  
   wire _Queue_29_io_deq_valid ;  
   wire [3:0] _Queue_29_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_29_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_29_io_deq_bits_extra_id ;  
   wire _Queue_28_io_enq_ready ;  
   wire _Queue_28_io_deq_valid ;  
   wire [3:0] _Queue_28_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_28_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_28_io_deq_bits_extra_id ;  
   wire _Queue_27_io_enq_ready ;  
   wire _Queue_27_io_deq_valid ;  
   wire [3:0] _Queue_27_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_27_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_27_io_deq_bits_extra_id ;  
   wire _Queue_26_io_enq_ready ;  
   wire _Queue_26_io_deq_valid ;  
   wire [3:0] _Queue_26_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_26_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_26_io_deq_bits_extra_id ;  
   wire _Queue_25_io_enq_ready ;  
   wire _Queue_25_io_deq_valid ;  
   wire [3:0] _Queue_25_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_25_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_25_io_deq_bits_extra_id ;  
   wire _Queue_24_io_enq_ready ;  
   wire _Queue_24_io_deq_valid ;  
   wire [3:0] _Queue_24_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_24_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_24_io_deq_bits_extra_id ;  
   wire _Queue_23_io_enq_ready ;  
   wire _Queue_23_io_deq_valid ;  
   wire [3:0] _Queue_23_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_23_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_23_io_deq_bits_extra_id ;  
   wire _Queue_22_io_enq_ready ;  
   wire _Queue_22_io_deq_valid ;  
   wire [3:0] _Queue_22_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_22_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_22_io_deq_bits_extra_id ;  
   wire _Queue_21_io_enq_ready ;  
   wire _Queue_21_io_deq_valid ;  
   wire [3:0] _Queue_21_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_21_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_21_io_deq_bits_extra_id ;  
   wire _Queue_20_io_enq_ready ;  
   wire _Queue_20_io_deq_valid ;  
   wire [3:0] _Queue_20_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_20_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_20_io_deq_bits_extra_id ;  
   wire _Queue_19_io_enq_ready ;  
   wire _Queue_19_io_deq_valid ;  
   wire [3:0] _Queue_19_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_19_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_19_io_deq_bits_extra_id ;  
   wire _Queue_18_io_enq_ready ;  
   wire _Queue_18_io_deq_valid ;  
   wire [3:0] _Queue_18_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_18_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_18_io_deq_bits_extra_id ;  
   wire _Queue_17_io_enq_ready ;  
   wire _Queue_17_io_deq_valid ;  
   wire [3:0] _Queue_17_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_17_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_17_io_deq_bits_extra_id ;  
   wire _Queue_16_io_enq_ready ;  
   wire _Queue_16_io_deq_valid ;  
   wire [3:0] _Queue_16_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_16_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_16_io_deq_bits_extra_id ;  
   wire _Queue_15_io_enq_ready ;  
   wire _Queue_15_io_deq_valid ;  
   wire [3:0] _Queue_15_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_15_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_15_io_deq_bits_extra_id ;  
   wire _Queue_14_io_enq_ready ;  
   wire _Queue_14_io_deq_valid ;  
   wire [3:0] _Queue_14_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_14_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_14_io_deq_bits_extra_id ;  
   wire _Queue_13_io_enq_ready ;  
   wire _Queue_13_io_deq_valid ;  
   wire [3:0] _Queue_13_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_13_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_13_io_deq_bits_extra_id ;  
   wire _Queue_12_io_enq_ready ;  
   wire _Queue_12_io_deq_valid ;  
   wire [3:0] _Queue_12_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_12_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_12_io_deq_bits_extra_id ;  
   wire _Queue_11_io_enq_ready ;  
   wire _Queue_11_io_deq_valid ;  
   wire [3:0] _Queue_11_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_11_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_11_io_deq_bits_extra_id ;  
   wire _Queue_10_io_enq_ready ;  
   wire _Queue_10_io_deq_valid ;  
   wire [3:0] _Queue_10_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_10_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_10_io_deq_bits_extra_id ;  
   wire _Queue_9_io_enq_ready ;  
   wire _Queue_9_io_deq_valid ;  
   wire [3:0] _Queue_9_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_9_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_9_io_deq_bits_extra_id ;  
   wire _Queue_8_io_enq_ready ;  
   wire _Queue_8_io_deq_valid ;  
   wire [3:0] _Queue_8_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_8_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_8_io_deq_bits_extra_id ;  
   wire _Queue_7_io_enq_ready ;  
   wire _Queue_7_io_deq_valid ;  
   wire [3:0] _Queue_7_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_7_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_7_io_deq_bits_extra_id ;  
   wire _Queue_6_io_enq_ready ;  
   wire _Queue_6_io_deq_valid ;  
   wire [3:0] _Queue_6_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_6_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_6_io_deq_bits_extra_id ;  
   wire _Queue_5_io_enq_ready ;  
   wire _Queue_5_io_deq_valid ;  
   wire [3:0] _Queue_5_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_5_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_5_io_deq_bits_extra_id ;  
   wire _Queue_4_io_enq_ready ;  
   wire _Queue_4_io_deq_valid ;  
   wire [3:0] _Queue_4_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_4_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_4_io_deq_bits_extra_id ;  
   wire _Queue_3_io_enq_ready ;  
   wire _Queue_3_io_deq_valid ;  
   wire [3:0] _Queue_3_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_3_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_3_io_deq_bits_extra_id ;  
   wire _Queue_2_io_enq_ready ;  
   wire _Queue_2_io_deq_valid ;  
   wire [3:0] _Queue_2_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_2_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_2_io_deq_bits_extra_id ;  
   wire _Queue_1_io_enq_ready ;  
   wire _Queue_1_io_deq_valid ;  
   wire [3:0] _Queue_1_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_1_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_1_io_deq_bits_extra_id ;  
   wire _Queue_io_enq_ready ;  
   wire _Queue_io_deq_valid ;  
   wire [3:0] _Queue_io_deq_bits_tl_state_size ;  
   wire [6:0] _Queue_io_deq_bits_tl_state_source ;  
   wire [2:0] _Queue_io_deq_bits_extra_id ;  
   reg casez_tmp ;  
  always @(*)
       begin 
         casez (auto_in_ar_bits_id)
          4 'b0000:
             casez_tmp =_Queue_io_enq_ready;
          4 'b0001:
             casez_tmp =_Queue_1_io_enq_ready;
          4 'b0010:
             casez_tmp =_Queue_2_io_enq_ready;
          4 'b0011:
             casez_tmp =_Queue_3_io_enq_ready;
          4 'b0100:
             casez_tmp =_Queue_4_io_enq_ready;
          4 'b0101:
             casez_tmp =_Queue_5_io_enq_ready;
          4 'b0110:
             casez_tmp =_Queue_6_io_enq_ready;
          4 'b0111:
             casez_tmp =_Queue_7_io_enq_ready;
          4 'b1000:
             casez_tmp =_Queue_8_io_enq_ready;
          4 'b1001:
             casez_tmp =_Queue_9_io_enq_ready;
          4 'b1010:
             casez_tmp =_Queue_10_io_enq_ready;
          4 'b1011:
             casez_tmp =_Queue_11_io_enq_ready;
          4 'b1100:
             casez_tmp =_Queue_12_io_enq_ready;
          4 'b1101:
             casez_tmp =_Queue_13_io_enq_ready;
          4 'b1110:
             casez_tmp =_Queue_14_io_enq_ready;
          default :
             casez_tmp =_Queue_15_io_enq_ready;
         endcase 
       end
  
   reg casez_tmp_0 ;  
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp_0 =_Queue_io_deq_valid;
          4 'b0001:
             casez_tmp_0 =_Queue_1_io_deq_valid;
          4 'b0010:
             casez_tmp_0 =_Queue_2_io_deq_valid;
          4 'b0011:
             casez_tmp_0 =_Queue_3_io_deq_valid;
          4 'b0100:
             casez_tmp_0 =_Queue_4_io_deq_valid;
          4 'b0101:
             casez_tmp_0 =_Queue_5_io_deq_valid;
          4 'b0110:
             casez_tmp_0 =_Queue_6_io_deq_valid;
          4 'b0111:
             casez_tmp_0 =_Queue_7_io_deq_valid;
          4 'b1000:
             casez_tmp_0 =_Queue_8_io_deq_valid;
          4 'b1001:
             casez_tmp_0 =_Queue_9_io_deq_valid;
          4 'b1010:
             casez_tmp_0 =_Queue_10_io_deq_valid;
          4 'b1011:
             casez_tmp_0 =_Queue_11_io_deq_valid;
          4 'b1100:
             casez_tmp_0 =_Queue_12_io_deq_valid;
          4 'b1101:
             casez_tmp_0 =_Queue_13_io_deq_valid;
          4 'b1110:
             casez_tmp_0 =_Queue_14_io_deq_valid;
          default :
             casez_tmp_0 =_Queue_15_io_deq_valid;
         endcase 
       end
  
   reg [3:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp_1 =_Queue_io_deq_bits_tl_state_size;
          4 'b0001:
             casez_tmp_1 =_Queue_1_io_deq_bits_tl_state_size;
          4 'b0010:
             casez_tmp_1 =_Queue_2_io_deq_bits_tl_state_size;
          4 'b0011:
             casez_tmp_1 =_Queue_3_io_deq_bits_tl_state_size;
          4 'b0100:
             casez_tmp_1 =_Queue_4_io_deq_bits_tl_state_size;
          4 'b0101:
             casez_tmp_1 =_Queue_5_io_deq_bits_tl_state_size;
          4 'b0110:
             casez_tmp_1 =_Queue_6_io_deq_bits_tl_state_size;
          4 'b0111:
             casez_tmp_1 =_Queue_7_io_deq_bits_tl_state_size;
          4 'b1000:
             casez_tmp_1 =_Queue_8_io_deq_bits_tl_state_size;
          4 'b1001:
             casez_tmp_1 =_Queue_9_io_deq_bits_tl_state_size;
          4 'b1010:
             casez_tmp_1 =_Queue_10_io_deq_bits_tl_state_size;
          4 'b1011:
             casez_tmp_1 =_Queue_11_io_deq_bits_tl_state_size;
          4 'b1100:
             casez_tmp_1 =_Queue_12_io_deq_bits_tl_state_size;
          4 'b1101:
             casez_tmp_1 =_Queue_13_io_deq_bits_tl_state_size;
          4 'b1110:
             casez_tmp_1 =_Queue_14_io_deq_bits_tl_state_size;
          default :
             casez_tmp_1 =_Queue_15_io_deq_bits_tl_state_size;
         endcase 
       end
  
   reg [6:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp_2 =_Queue_io_deq_bits_tl_state_source;
          4 'b0001:
             casez_tmp_2 =_Queue_1_io_deq_bits_tl_state_source;
          4 'b0010:
             casez_tmp_2 =_Queue_2_io_deq_bits_tl_state_source;
          4 'b0011:
             casez_tmp_2 =_Queue_3_io_deq_bits_tl_state_source;
          4 'b0100:
             casez_tmp_2 =_Queue_4_io_deq_bits_tl_state_source;
          4 'b0101:
             casez_tmp_2 =_Queue_5_io_deq_bits_tl_state_source;
          4 'b0110:
             casez_tmp_2 =_Queue_6_io_deq_bits_tl_state_source;
          4 'b0111:
             casez_tmp_2 =_Queue_7_io_deq_bits_tl_state_source;
          4 'b1000:
             casez_tmp_2 =_Queue_8_io_deq_bits_tl_state_source;
          4 'b1001:
             casez_tmp_2 =_Queue_9_io_deq_bits_tl_state_source;
          4 'b1010:
             casez_tmp_2 =_Queue_10_io_deq_bits_tl_state_source;
          4 'b1011:
             casez_tmp_2 =_Queue_11_io_deq_bits_tl_state_source;
          4 'b1100:
             casez_tmp_2 =_Queue_12_io_deq_bits_tl_state_source;
          4 'b1101:
             casez_tmp_2 =_Queue_13_io_deq_bits_tl_state_source;
          4 'b1110:
             casez_tmp_2 =_Queue_14_io_deq_bits_tl_state_source;
          default :
             casez_tmp_2 =_Queue_15_io_deq_bits_tl_state_source;
         endcase 
       end
  
   reg [2:0] casez_tmp_3 ;  
  always @(*)
       begin 
         casez (auto_out_r_bits_id)
          4 'b0000:
             casez_tmp_3 =_Queue_io_deq_bits_extra_id;
          4 'b0001:
             casez_tmp_3 =_Queue_1_io_deq_bits_extra_id;
          4 'b0010:
             casez_tmp_3 =_Queue_2_io_deq_bits_extra_id;
          4 'b0011:
             casez_tmp_3 =_Queue_3_io_deq_bits_extra_id;
          4 'b0100:
             casez_tmp_3 =_Queue_4_io_deq_bits_extra_id;
          4 'b0101:
             casez_tmp_3 =_Queue_5_io_deq_bits_extra_id;
          4 'b0110:
             casez_tmp_3 =_Queue_6_io_deq_bits_extra_id;
          4 'b0111:
             casez_tmp_3 =_Queue_7_io_deq_bits_extra_id;
          4 'b1000:
             casez_tmp_3 =_Queue_8_io_deq_bits_extra_id;
          4 'b1001:
             casez_tmp_3 =_Queue_9_io_deq_bits_extra_id;
          4 'b1010:
             casez_tmp_3 =_Queue_10_io_deq_bits_extra_id;
          4 'b1011:
             casez_tmp_3 =_Queue_11_io_deq_bits_extra_id;
          4 'b1100:
             casez_tmp_3 =_Queue_12_io_deq_bits_extra_id;
          4 'b1101:
             casez_tmp_3 =_Queue_13_io_deq_bits_extra_id;
          4 'b1110:
             casez_tmp_3 =_Queue_14_io_deq_bits_extra_id;
          default :
             casez_tmp_3 =_Queue_15_io_deq_bits_extra_id;
         endcase 
       end
  
   wire _GEN=auto_out_r_valid&auto_in_r_ready ;  
   wire _GEN_0=auto_in_ar_valid&auto_out_ar_ready ;  
   reg casez_tmp_4 ;  
  always @(*)
       begin 
         casez (auto_in_aw_bits_id)
          4 'b0000:
             casez_tmp_4 =_Queue_16_io_enq_ready;
          4 'b0001:
             casez_tmp_4 =_Queue_17_io_enq_ready;
          4 'b0010:
             casez_tmp_4 =_Queue_18_io_enq_ready;
          4 'b0011:
             casez_tmp_4 =_Queue_19_io_enq_ready;
          4 'b0100:
             casez_tmp_4 =_Queue_20_io_enq_ready;
          4 'b0101:
             casez_tmp_4 =_Queue_21_io_enq_ready;
          4 'b0110:
             casez_tmp_4 =_Queue_22_io_enq_ready;
          4 'b0111:
             casez_tmp_4 =_Queue_23_io_enq_ready;
          4 'b1000:
             casez_tmp_4 =_Queue_24_io_enq_ready;
          4 'b1001:
             casez_tmp_4 =_Queue_25_io_enq_ready;
          4 'b1010:
             casez_tmp_4 =_Queue_26_io_enq_ready;
          4 'b1011:
             casez_tmp_4 =_Queue_27_io_enq_ready;
          4 'b1100:
             casez_tmp_4 =_Queue_28_io_enq_ready;
          4 'b1101:
             casez_tmp_4 =_Queue_29_io_enq_ready;
          4 'b1110:
             casez_tmp_4 =_Queue_30_io_enq_ready;
          default :
             casez_tmp_4 =_Queue_31_io_enq_ready;
         endcase 
       end
  
   reg casez_tmp_5 ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp_5 =_Queue_16_io_deq_valid;
          4 'b0001:
             casez_tmp_5 =_Queue_17_io_deq_valid;
          4 'b0010:
             casez_tmp_5 =_Queue_18_io_deq_valid;
          4 'b0011:
             casez_tmp_5 =_Queue_19_io_deq_valid;
          4 'b0100:
             casez_tmp_5 =_Queue_20_io_deq_valid;
          4 'b0101:
             casez_tmp_5 =_Queue_21_io_deq_valid;
          4 'b0110:
             casez_tmp_5 =_Queue_22_io_deq_valid;
          4 'b0111:
             casez_tmp_5 =_Queue_23_io_deq_valid;
          4 'b1000:
             casez_tmp_5 =_Queue_24_io_deq_valid;
          4 'b1001:
             casez_tmp_5 =_Queue_25_io_deq_valid;
          4 'b1010:
             casez_tmp_5 =_Queue_26_io_deq_valid;
          4 'b1011:
             casez_tmp_5 =_Queue_27_io_deq_valid;
          4 'b1100:
             casez_tmp_5 =_Queue_28_io_deq_valid;
          4 'b1101:
             casez_tmp_5 =_Queue_29_io_deq_valid;
          4 'b1110:
             casez_tmp_5 =_Queue_30_io_deq_valid;
          default :
             casez_tmp_5 =_Queue_31_io_deq_valid;
         endcase 
       end
  
  always @( posedge clock)
       begin 
         if (~reset&~(~auto_out_r_valid|casez_tmp_0))
            begin 
              if (1)$display("Assertion failed\n    at UserYanker.scala:66 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
              if (1)$display("");
            end 
         if (~reset&~(~auto_out_b_valid|casez_tmp_5))
            begin 
              if (1)$display("Assertion failed\n    at UserYanker.scala:95 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
              if (1)$display("");
            end 
       end
  
   reg [3:0] casez_tmp_6 ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp_6 =_Queue_16_io_deq_bits_tl_state_size;
          4 'b0001:
             casez_tmp_6 =_Queue_17_io_deq_bits_tl_state_size;
          4 'b0010:
             casez_tmp_6 =_Queue_18_io_deq_bits_tl_state_size;
          4 'b0011:
             casez_tmp_6 =_Queue_19_io_deq_bits_tl_state_size;
          4 'b0100:
             casez_tmp_6 =_Queue_20_io_deq_bits_tl_state_size;
          4 'b0101:
             casez_tmp_6 =_Queue_21_io_deq_bits_tl_state_size;
          4 'b0110:
             casez_tmp_6 =_Queue_22_io_deq_bits_tl_state_size;
          4 'b0111:
             casez_tmp_6 =_Queue_23_io_deq_bits_tl_state_size;
          4 'b1000:
             casez_tmp_6 =_Queue_24_io_deq_bits_tl_state_size;
          4 'b1001:
             casez_tmp_6 =_Queue_25_io_deq_bits_tl_state_size;
          4 'b1010:
             casez_tmp_6 =_Queue_26_io_deq_bits_tl_state_size;
          4 'b1011:
             casez_tmp_6 =_Queue_27_io_deq_bits_tl_state_size;
          4 'b1100:
             casez_tmp_6 =_Queue_28_io_deq_bits_tl_state_size;
          4 'b1101:
             casez_tmp_6 =_Queue_29_io_deq_bits_tl_state_size;
          4 'b1110:
             casez_tmp_6 =_Queue_30_io_deq_bits_tl_state_size;
          default :
             casez_tmp_6 =_Queue_31_io_deq_bits_tl_state_size;
         endcase 
       end
  
   reg [6:0] casez_tmp_7 ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp_7 =_Queue_16_io_deq_bits_tl_state_source;
          4 'b0001:
             casez_tmp_7 =_Queue_17_io_deq_bits_tl_state_source;
          4 'b0010:
             casez_tmp_7 =_Queue_18_io_deq_bits_tl_state_source;
          4 'b0011:
             casez_tmp_7 =_Queue_19_io_deq_bits_tl_state_source;
          4 'b0100:
             casez_tmp_7 =_Queue_20_io_deq_bits_tl_state_source;
          4 'b0101:
             casez_tmp_7 =_Queue_21_io_deq_bits_tl_state_source;
          4 'b0110:
             casez_tmp_7 =_Queue_22_io_deq_bits_tl_state_source;
          4 'b0111:
             casez_tmp_7 =_Queue_23_io_deq_bits_tl_state_source;
          4 'b1000:
             casez_tmp_7 =_Queue_24_io_deq_bits_tl_state_source;
          4 'b1001:
             casez_tmp_7 =_Queue_25_io_deq_bits_tl_state_source;
          4 'b1010:
             casez_tmp_7 =_Queue_26_io_deq_bits_tl_state_source;
          4 'b1011:
             casez_tmp_7 =_Queue_27_io_deq_bits_tl_state_source;
          4 'b1100:
             casez_tmp_7 =_Queue_28_io_deq_bits_tl_state_source;
          4 'b1101:
             casez_tmp_7 =_Queue_29_io_deq_bits_tl_state_source;
          4 'b1110:
             casez_tmp_7 =_Queue_30_io_deq_bits_tl_state_source;
          default :
             casez_tmp_7 =_Queue_31_io_deq_bits_tl_state_source;
         endcase 
       end
  
   reg [2:0] casez_tmp_8 ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp_8 =_Queue_16_io_deq_bits_extra_id;
          4 'b0001:
             casez_tmp_8 =_Queue_17_io_deq_bits_extra_id;
          4 'b0010:
             casez_tmp_8 =_Queue_18_io_deq_bits_extra_id;
          4 'b0011:
             casez_tmp_8 =_Queue_19_io_deq_bits_extra_id;
          4 'b0100:
             casez_tmp_8 =_Queue_20_io_deq_bits_extra_id;
          4 'b0101:
             casez_tmp_8 =_Queue_21_io_deq_bits_extra_id;
          4 'b0110:
             casez_tmp_8 =_Queue_22_io_deq_bits_extra_id;
          4 'b0111:
             casez_tmp_8 =_Queue_23_io_deq_bits_extra_id;
          4 'b1000:
             casez_tmp_8 =_Queue_24_io_deq_bits_extra_id;
          4 'b1001:
             casez_tmp_8 =_Queue_25_io_deq_bits_extra_id;
          4 'b1010:
             casez_tmp_8 =_Queue_26_io_deq_bits_extra_id;
          4 'b1011:
             casez_tmp_8 =_Queue_27_io_deq_bits_extra_id;
          4 'b1100:
             casez_tmp_8 =_Queue_28_io_deq_bits_extra_id;
          4 'b1101:
             casez_tmp_8 =_Queue_29_io_deq_bits_extra_id;
          4 'b1110:
             casez_tmp_8 =_Queue_30_io_deq_bits_extra_id;
          default :
             casez_tmp_8 =_Queue_31_io_deq_bits_extra_id;
         endcase 
       end
  
   wire _GEN_1=auto_out_b_valid&auto_in_b_ready ;  
   wire _GEN_2=auto_in_aw_valid&auto_out_aw_ready ;  
  Queue_40 Queue(.clock(clock),.reset(reset),.io_enq_ready(_Queue_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h0),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h0&auto_out_r_bits_last),.io_deq_valid(_Queue_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_io_deq_bits_extra_id)); 
  Queue_40 Queue_1(.clock(clock),.reset(reset),.io_enq_ready(_Queue_1_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h1),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h1&auto_out_r_bits_last),.io_deq_valid(_Queue_1_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_1_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_1_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_1_io_deq_bits_extra_id)); 
  Queue_40 Queue_2(.clock(clock),.reset(reset),.io_enq_ready(_Queue_2_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h2),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h2&auto_out_r_bits_last),.io_deq_valid(_Queue_2_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_2_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_2_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_2_io_deq_bits_extra_id)); 
  Queue_40 Queue_3(.clock(clock),.reset(reset),.io_enq_ready(_Queue_3_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h3),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h3&auto_out_r_bits_last),.io_deq_valid(_Queue_3_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_3_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_3_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_3_io_deq_bits_extra_id)); 
  Queue_40 Queue_4(.clock(clock),.reset(reset),.io_enq_ready(_Queue_4_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h4),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h4&auto_out_r_bits_last),.io_deq_valid(_Queue_4_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_4_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_4_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_4_io_deq_bits_extra_id)); 
  Queue_40 Queue_5(.clock(clock),.reset(reset),.io_enq_ready(_Queue_5_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h5),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h5&auto_out_r_bits_last),.io_deq_valid(_Queue_5_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_5_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_5_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_5_io_deq_bits_extra_id)); 
  Queue_40 Queue_6(.clock(clock),.reset(reset),.io_enq_ready(_Queue_6_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h6),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h6&auto_out_r_bits_last),.io_deq_valid(_Queue_6_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_6_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_6_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_6_io_deq_bits_extra_id)); 
  Queue_40 Queue_7(.clock(clock),.reset(reset),.io_enq_ready(_Queue_7_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h7),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h7&auto_out_r_bits_last),.io_deq_valid(_Queue_7_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_7_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_7_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_7_io_deq_bits_extra_id)); 
  Queue_40 Queue_8(.clock(clock),.reset(reset),.io_enq_ready(_Queue_8_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h8),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h8&auto_out_r_bits_last),.io_deq_valid(_Queue_8_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_8_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_8_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_8_io_deq_bits_extra_id)); 
  Queue_40 Queue_9(.clock(clock),.reset(reset),.io_enq_ready(_Queue_9_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'h9),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'h9&auto_out_r_bits_last),.io_deq_valid(_Queue_9_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_9_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_9_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_9_io_deq_bits_extra_id)); 
  Queue_40 Queue_10(.clock(clock),.reset(reset),.io_enq_ready(_Queue_10_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'hA),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'hA&auto_out_r_bits_last),.io_deq_valid(_Queue_10_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_10_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_10_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_10_io_deq_bits_extra_id)); 
  Queue_40 Queue_11(.clock(clock),.reset(reset),.io_enq_ready(_Queue_11_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'hB),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'hB&auto_out_r_bits_last),.io_deq_valid(_Queue_11_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_11_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_11_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_11_io_deq_bits_extra_id)); 
  Queue_40 Queue_12(.clock(clock),.reset(reset),.io_enq_ready(_Queue_12_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'hC),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'hC&auto_out_r_bits_last),.io_deq_valid(_Queue_12_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_12_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_12_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_12_io_deq_bits_extra_id)); 
  Queue_40 Queue_13(.clock(clock),.reset(reset),.io_enq_ready(_Queue_13_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'hD),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'hD&auto_out_r_bits_last),.io_deq_valid(_Queue_13_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_13_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_13_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_13_io_deq_bits_extra_id)); 
  Queue_40 Queue_14(.clock(clock),.reset(reset),.io_enq_ready(_Queue_14_io_enq_ready),.io_enq_valid(_GEN_0&auto_in_ar_bits_id==4'hE),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&auto_out_r_bits_id==4'hE&auto_out_r_bits_last),.io_deq_valid(_Queue_14_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_14_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_14_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_14_io_deq_bits_extra_id)); 
  Queue_40 Queue_15(.clock(clock),.reset(reset),.io_enq_ready(_Queue_15_io_enq_ready),.io_enq_valid(_GEN_0&(&auto_in_ar_bits_id)),.io_enq_bits_tl_state_size(auto_in_ar_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_ar_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_ar_bits_echo_extra_id),.io_deq_ready(_GEN&(&auto_out_r_bits_id)&auto_out_r_bits_last),.io_deq_valid(_Queue_15_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_15_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_15_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_15_io_deq_bits_extra_id)); 
  Queue_40 Queue_16(.clock(clock),.reset(reset),.io_enq_ready(_Queue_16_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h0),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h0),.io_deq_valid(_Queue_16_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_16_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_16_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_16_io_deq_bits_extra_id)); 
  Queue_40 Queue_17(.clock(clock),.reset(reset),.io_enq_ready(_Queue_17_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h1),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h1),.io_deq_valid(_Queue_17_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_17_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_17_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_17_io_deq_bits_extra_id)); 
  Queue_40 Queue_18(.clock(clock),.reset(reset),.io_enq_ready(_Queue_18_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h2),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h2),.io_deq_valid(_Queue_18_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_18_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_18_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_18_io_deq_bits_extra_id)); 
  Queue_40 Queue_19(.clock(clock),.reset(reset),.io_enq_ready(_Queue_19_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h3),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h3),.io_deq_valid(_Queue_19_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_19_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_19_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_19_io_deq_bits_extra_id)); 
  Queue_40 Queue_20(.clock(clock),.reset(reset),.io_enq_ready(_Queue_20_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h4),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h4),.io_deq_valid(_Queue_20_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_20_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_20_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_20_io_deq_bits_extra_id)); 
  Queue_40 Queue_21(.clock(clock),.reset(reset),.io_enq_ready(_Queue_21_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h5),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h5),.io_deq_valid(_Queue_21_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_21_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_21_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_21_io_deq_bits_extra_id)); 
  Queue_40 Queue_22(.clock(clock),.reset(reset),.io_enq_ready(_Queue_22_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h6),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h6),.io_deq_valid(_Queue_22_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_22_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_22_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_22_io_deq_bits_extra_id)); 
  Queue_40 Queue_23(.clock(clock),.reset(reset),.io_enq_ready(_Queue_23_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h7),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h7),.io_deq_valid(_Queue_23_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_23_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_23_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_23_io_deq_bits_extra_id)); 
  Queue_40 Queue_24(.clock(clock),.reset(reset),.io_enq_ready(_Queue_24_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h8),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h8),.io_deq_valid(_Queue_24_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_24_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_24_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_24_io_deq_bits_extra_id)); 
  Queue_40 Queue_25(.clock(clock),.reset(reset),.io_enq_ready(_Queue_25_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'h9),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'h9),.io_deq_valid(_Queue_25_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_25_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_25_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_25_io_deq_bits_extra_id)); 
  Queue_40 Queue_26(.clock(clock),.reset(reset),.io_enq_ready(_Queue_26_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'hA),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'hA),.io_deq_valid(_Queue_26_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_26_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_26_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_26_io_deq_bits_extra_id)); 
  Queue_40 Queue_27(.clock(clock),.reset(reset),.io_enq_ready(_Queue_27_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'hB),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'hB),.io_deq_valid(_Queue_27_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_27_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_27_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_27_io_deq_bits_extra_id)); 
  Queue_40 Queue_28(.clock(clock),.reset(reset),.io_enq_ready(_Queue_28_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'hC),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'hC),.io_deq_valid(_Queue_28_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_28_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_28_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_28_io_deq_bits_extra_id)); 
  Queue_40 Queue_29(.clock(clock),.reset(reset),.io_enq_ready(_Queue_29_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'hD),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'hD),.io_deq_valid(_Queue_29_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_29_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_29_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_29_io_deq_bits_extra_id)); 
  Queue_40 Queue_30(.clock(clock),.reset(reset),.io_enq_ready(_Queue_30_io_enq_ready),.io_enq_valid(_GEN_2&auto_in_aw_bits_id==4'hE),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&auto_out_b_bits_id==4'hE),.io_deq_valid(_Queue_30_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_30_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_30_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_30_io_deq_bits_extra_id)); 
  Queue_40 Queue_31(.clock(clock),.reset(reset),.io_enq_ready(_Queue_31_io_enq_ready),.io_enq_valid(_GEN_2&(&auto_in_aw_bits_id)),.io_enq_bits_tl_state_size(auto_in_aw_bits_echo_tl_state_size),.io_enq_bits_tl_state_source(auto_in_aw_bits_echo_tl_state_source),.io_enq_bits_extra_id(auto_in_aw_bits_echo_extra_id),.io_deq_ready(_GEN_1&(&auto_out_b_bits_id)),.io_deq_valid(_Queue_31_io_deq_valid),.io_deq_bits_tl_state_size(_Queue_31_io_deq_bits_tl_state_size),.io_deq_bits_tl_state_source(_Queue_31_io_deq_bits_tl_state_source),.io_deq_bits_extra_id(_Queue_31_io_deq_bits_extra_id)); 
  assign auto_in_aw_ready=auto_out_aw_ready&casez_tmp_4; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_b_bits_echo_tl_state_size=casez_tmp_6; 
  assign auto_in_b_bits_echo_tl_state_source=casez_tmp_7; 
  assign auto_in_b_bits_echo_extra_id=casez_tmp_8; 
  assign auto_in_ar_ready=auto_out_ar_ready&casez_tmp; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_echo_tl_state_size=casez_tmp_1; 
  assign auto_in_r_bits_echo_tl_state_source=casez_tmp_2; 
  assign auto_in_r_bits_echo_extra_id=casez_tmp_3; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid&casez_tmp_4; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid&casez_tmp; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module AXI4IdIndexer_2 (
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [6:0] auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [3:0] auto_in_aw_bits_echo_tl_state_size,
  input [6:0] auto_in_aw_bits_echo_tl_state_source,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [6:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output [3:0] auto_in_b_bits_echo_tl_state_size,
  output [6:0] auto_in_b_bits_echo_tl_state_source,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [6:0] auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [3:0] auto_in_ar_bits_echo_tl_state_size,
  input [6:0] auto_in_ar_bits_echo_tl_state_source,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [6:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output [3:0] auto_in_r_bits_echo_tl_state_size,
  output [6:0] auto_in_r_bits_echo_tl_state_source,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [3:0] auto_out_aw_bits_echo_tl_state_size,
  output [6:0] auto_out_aw_bits_echo_tl_state_source,
  output [2:0] auto_out_aw_bits_echo_extra_id,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input [3:0] auto_out_b_bits_echo_tl_state_size,
  input [6:0] auto_out_b_bits_echo_tl_state_source,
  input [2:0] auto_out_b_bits_echo_extra_id,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [3:0] auto_out_ar_bits_echo_tl_state_size,
  output [6:0] auto_out_ar_bits_echo_tl_state_source,
  output [2:0] auto_out_ar_bits_echo_extra_id,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input [3:0] auto_out_r_bits_echo_tl_state_size,
  input [6:0] auto_out_r_bits_echo_tl_state_source,
  input [2:0] auto_out_r_bits_echo_extra_id,
  input auto_out_r_bits_last) ; 
  assign auto_in_aw_ready=auto_out_aw_ready; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id={auto_out_b_bits_echo_extra_id,auto_out_b_bits_id}; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_b_bits_echo_tl_state_size=auto_out_b_bits_echo_tl_state_size; 
  assign auto_in_b_bits_echo_tl_state_source=auto_out_b_bits_echo_tl_state_source; 
  assign auto_in_ar_ready=auto_out_ar_ready; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id={auto_out_r_bits_echo_extra_id,auto_out_r_bits_id}; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_echo_tl_state_size=auto_out_r_bits_echo_tl_state_size; 
  assign auto_in_r_bits_echo_tl_state_source=auto_out_r_bits_echo_tl_state_source; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id[3:0]; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_aw_bits_echo_tl_state_size=auto_in_aw_bits_echo_tl_state_size; 
  assign auto_out_aw_bits_echo_tl_state_source=auto_in_aw_bits_echo_tl_state_source; 
  assign auto_out_aw_bits_echo_extra_id=auto_in_aw_bits_id[6:4]; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id[3:0]; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_ar_bits_echo_tl_state_size=auto_in_ar_bits_echo_tl_state_size; 
  assign auto_out_ar_bits_echo_tl_state_source=auto_in_ar_bits_echo_tl_state_source; 
  assign auto_out_ar_bits_echo_extra_id=auto_in_ar_bits_id[6:4]; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module TLMonitor_20 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [6:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [2:0] io_in_d_bits_size,
  input [6:0] io_in_d_bits_source,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [6:0] source ;  
   reg [31:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [2:0] size_1 ;  
   reg [6:0] source_1 ;  
   reg denied ;  
   reg [127:0] inflight ;  
   reg [511:0] inflight_opcodes ;  
   reg [511:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [511:0] _GEN_0={503'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_0 ;  
   wire [127:0] _GEN_1={121'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [127:0] _GEN_3={121'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [127:0] inflight_1 ;  
   reg [511:0] inflight_sizes_1 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_4=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_a_bits_param>3'h2 ;  
   wire _GEN_7=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_8=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_9=io_in_a_bits_size!=3'h7&io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_11=io_in_a_bits_mask!=mask ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_18=io_in_d_bits_size<3'h3 ;  
   wire _GEN_19=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_20=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_21=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_22=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_23=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [127:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 128'h1<<_GEN_1:128'h0 ;  
   wire _GEN_24=io_in_d_valid&d_first_1 ;  
   wire _GEN_25=_GEN_24&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_26=_GEN_25&same_cycle_resp&~reset ;  
   wire _GEN_27=_GEN_25&~same_cycle_resp&~reset ;  
   wire _GEN_28=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [127:0] _GEN_29=inflight>>_GEN_1 ;  
   wire [127:0] _GEN_30=inflight>>_GEN_3 ;  
   wire [511:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_0 ;  
   wire [127:0] _GEN_31=inflight_1>>_GEN_3 ;  
   wire [511:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_0 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_29[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~reset&~(_GEN_30[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_25 ? 128'h1<<_GEN_3:128'h0)|a_set_wo_ready==128'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==128'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(_GEN_31[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==128'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/Ports.scala:91:9)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_32={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_32 ;  
   wire [1026:0] _GEN_33={1018'h0,io_in_a_bits_source,2'h0} ;  
   wire [1038:0] _GEN_34={1030'h0,io_in_d_bits_source,2'h0} ;  
   wire [1038:0] _d_opcodes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_opcodes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_sizes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_11=1039'hF<<_GEN_34 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_35=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_36=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=128'h0;
              inflight_opcodes <=512'h0;
              inflight_sizes <=512'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=128'h0;
              inflight_sizes_1 <=512'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_2 ? 128'h1<<_GEN_1:128'h0))&~(_GEN_35 ? 128'h1<<_GEN_3:128'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_opcodes_clr_T_5[511:0]:512'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_sizes_clr_T_5[511:0]:512'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_36 ? 128'h1<<_GEN_3:128'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_36 ? _d_sizes_clr_T_11[511:0]:512'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module Queue_73 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [6:0] io_enq_bits_id,
  input [31:0] io_enq_bits_addr,
  input [7:0] io_enq_bits_len,
  input [2:0] io_enq_bits_size,
  input [3:0] io_enq_bits_echo_tl_state_size,
  input [6:0] io_enq_bits_echo_tl_state_source,
  input io_enq_bits_wen,
  input io_deq_ready,
  output io_deq_valid,
  output [6:0] io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [3:0] io_deq_bits_echo_tl_state_size,
  output [6:0] io_deq_bits_echo_tl_state_source,
  output io_deq_bits_wen) ; 
   reg ram_wen ;  
   reg [2:0] ram_size ;  
   reg [7:0] ram_len ;  
   reg [31:0] ram_addr ;  
   reg [6:0] ram_id ;  
   reg [10:0] ram_echo ;  
   reg full ;  
   wire io_enq_ready_0=io_deq_ready|~full ;  
   wire do_enq=io_enq_ready_0&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_wen <=io_enq_bits_wen;
              ram_size <=io_enq_bits_size;
              ram_len <=io_enq_bits_len;
              ram_addr <=io_enq_bits_addr;
              ram_id <=io_enq_bits_id;
              ram_echo <={io_enq_bits_echo_tl_state_source,io_enq_bits_echo_tl_state_size};
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(io_deq_ready&full)))
               full <=do_enq;
       end
  
  assign io_enq_ready=io_enq_ready_0; 
  assign io_deq_valid=full; 
  assign io_deq_bits_id=ram_id; 
  assign io_deq_bits_addr=ram_addr; 
  assign io_deq_bits_len=ram_len; 
  assign io_deq_bits_size=ram_size; 
  assign io_deq_bits_echo_tl_state_size=ram_echo[3:0]; 
  assign io_deq_bits_echo_tl_state_source=ram_echo[10:4]; 
  assign io_deq_bits_wen=ram_wen; 
endmodule
 
module TLToAXI4_1 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [6:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [2:0] auto_in_d_bits_size,
  output [6:0] auto_in_d_bits_source,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [6:0] auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [3:0] auto_out_aw_bits_echo_tl_state_size,
  output [6:0] auto_out_aw_bits_echo_tl_state_source,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [6:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input [3:0] auto_out_b_bits_echo_tl_state_size,
  input [6:0] auto_out_b_bits_echo_tl_state_source,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [6:0] auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [3:0] auto_out_ar_bits_echo_tl_state_size,
  output [6:0] auto_out_ar_bits_echo_tl_state_source,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [6:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input [3:0] auto_out_r_bits_echo_tl_state_size,
  input [6:0] auto_out_r_bits_echo_tl_state_source,
  input auto_out_r_bits_last) ; 
   reg count_128 ;  
   reg count_127 ;  
   reg count_126 ;  
   reg count_125 ;  
   reg count_124 ;  
   reg count_123 ;  
   reg count_122 ;  
   reg count_121 ;  
   reg count_120 ;  
   reg count_119 ;  
   reg count_118 ;  
   reg count_117 ;  
   reg count_116 ;  
   reg count_115 ;  
   reg count_114 ;  
   reg count_113 ;  
   reg count_112 ;  
   reg count_111 ;  
   reg count_110 ;  
   reg count_109 ;  
   reg count_108 ;  
   reg count_107 ;  
   reg count_106 ;  
   reg count_105 ;  
   reg count_104 ;  
   reg count_103 ;  
   reg count_102 ;  
   reg count_101 ;  
   reg count_100 ;  
   reg count_99 ;  
   reg count_98 ;  
   reg count_97 ;  
   reg count_96 ;  
   reg count_95 ;  
   reg count_94 ;  
   reg count_93 ;  
   reg count_92 ;  
   reg count_91 ;  
   reg count_90 ;  
   reg count_89 ;  
   reg count_88 ;  
   reg count_87 ;  
   reg count_86 ;  
   reg count_85 ;  
   reg count_84 ;  
   reg count_83 ;  
   reg count_82 ;  
   reg count_81 ;  
   reg count_80 ;  
   reg count_79 ;  
   reg count_78 ;  
   reg count_77 ;  
   reg count_76 ;  
   reg count_75 ;  
   reg count_74 ;  
   reg count_73 ;  
   reg count_72 ;  
   reg count_71 ;  
   reg count_70 ;  
   reg count_69 ;  
   reg count_68 ;  
   reg count_67 ;  
   reg count_66 ;  
   reg count_65 ;  
   reg count_64 ;  
   reg count_63 ;  
   reg count_62 ;  
   reg count_61 ;  
   reg count_60 ;  
   reg count_59 ;  
   reg count_58 ;  
   reg count_57 ;  
   reg count_56 ;  
   reg count_55 ;  
   reg count_54 ;  
   reg count_53 ;  
   reg count_52 ;  
   reg count_51 ;  
   reg count_50 ;  
   reg count_49 ;  
   reg count_48 ;  
   reg count_47 ;  
   reg count_46 ;  
   reg count_45 ;  
   reg count_44 ;  
   reg count_43 ;  
   reg count_42 ;  
   reg count_41 ;  
   reg count_40 ;  
   reg count_39 ;  
   reg count_38 ;  
   reg count_37 ;  
   reg count_36 ;  
   reg count_35 ;  
   reg count_34 ;  
   reg count_33 ;  
   reg count_32 ;  
   reg count_31 ;  
   reg count_30 ;  
   reg count_29 ;  
   reg count_28 ;  
   reg count_27 ;  
   reg count_26 ;  
   reg count_25 ;  
   reg count_24 ;  
   reg count_23 ;  
   reg count_22 ;  
   reg count_21 ;  
   reg count_20 ;  
   reg count_19 ;  
   reg count_18 ;  
   reg count_17 ;  
   reg count_16 ;  
   reg count_15 ;  
   reg count_14 ;  
   reg count_13 ;  
   reg count_12 ;  
   reg count_11 ;  
   reg count_10 ;  
   reg count_9 ;  
   reg count_8 ;  
   reg count_7 ;  
   reg count_6 ;  
   reg count_5 ;  
   reg count_4 ;  
   reg count_3 ;  
   reg count_2 ;  
   reg count_1 ;  
   wire _queue_arw_deq_q_io_enq_ready ;  
   wire _queue_arw_deq_q_io_deq_valid ;  
   wire [6:0] _queue_arw_deq_q_io_deq_bits_id ;  
   wire [31:0] _queue_arw_deq_q_io_deq_bits_addr ;  
   wire [7:0] _queue_arw_deq_q_io_deq_bits_len ;  
   wire [2:0] _queue_arw_deq_q_io_deq_bits_size ;  
   wire [3:0] _queue_arw_deq_q_io_deq_bits_echo_tl_state_size ;  
   wire [6:0] _queue_arw_deq_q_io_deq_bits_echo_tl_state_source ;  
   wire _queue_arw_deq_q_io_deq_bits_wen ;  
   wire _nodeOut_w_deq_q_io_enq_ready ;  
   wire [12:0] _beats1_decode_T_1=13'h3F<<auto_in_a_bits_size ;  
   wire [2:0] beats1=auto_in_a_bits_opcode[2] ? 3'h0:~(_beats1_decode_T_1[5:3]) ;  
   reg [2:0] counter ;  
   wire a_first=counter==3'h0 ;  
   wire a_last=counter==3'h1|beats1==3'h0 ;  
   reg doneAW ;  
   reg [6:0] casez_tmp ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_source)
          7 'b0000000:
             casez_tmp =7'h0;
          7 'b0000001:
             casez_tmp =7'h1;
          7 'b0000010:
             casez_tmp =7'h2;
          7 'b0000011:
             casez_tmp =7'h3;
          7 'b0000100:
             casez_tmp =7'h4;
          7 'b0000101:
             casez_tmp =7'h5;
          7 'b0000110:
             casez_tmp =7'h6;
          7 'b0000111:
             casez_tmp =7'h7;
          7 'b0001000:
             casez_tmp =7'h8;
          7 'b0001001:
             casez_tmp =7'h9;
          7 'b0001010:
             casez_tmp =7'hA;
          7 'b0001011:
             casez_tmp =7'hB;
          7 'b0001100:
             casez_tmp =7'hC;
          7 'b0001101:
             casez_tmp =7'hD;
          7 'b0001110:
             casez_tmp =7'hE;
          7 'b0001111:
             casez_tmp =7'hF;
          7 'b0010000:
             casez_tmp =7'h10;
          7 'b0010001:
             casez_tmp =7'h11;
          7 'b0010010:
             casez_tmp =7'h12;
          7 'b0010011:
             casez_tmp =7'h13;
          7 'b0010100:
             casez_tmp =7'h14;
          7 'b0010101:
             casez_tmp =7'h15;
          7 'b0010110:
             casez_tmp =7'h16;
          7 'b0010111:
             casez_tmp =7'h17;
          7 'b0011000:
             casez_tmp =7'h18;
          7 'b0011001:
             casez_tmp =7'h19;
          7 'b0011010:
             casez_tmp =7'h1A;
          7 'b0011011:
             casez_tmp =7'h1B;
          7 'b0011100:
             casez_tmp =7'h1C;
          7 'b0011101:
             casez_tmp =7'h1D;
          7 'b0011110:
             casez_tmp =7'h1E;
          7 'b0011111:
             casez_tmp =7'h1F;
          7 'b0100000:
             casez_tmp =7'h20;
          7 'b0100001:
             casez_tmp =7'h21;
          7 'b0100010:
             casez_tmp =7'h22;
          7 'b0100011:
             casez_tmp =7'h23;
          7 'b0100100:
             casez_tmp =7'h24;
          7 'b0100101:
             casez_tmp =7'h25;
          7 'b0100110:
             casez_tmp =7'h26;
          7 'b0100111:
             casez_tmp =7'h27;
          7 'b0101000:
             casez_tmp =7'h28;
          7 'b0101001:
             casez_tmp =7'h29;
          7 'b0101010:
             casez_tmp =7'h2A;
          7 'b0101011:
             casez_tmp =7'h2B;
          7 'b0101100:
             casez_tmp =7'h2C;
          7 'b0101101:
             casez_tmp =7'h2D;
          7 'b0101110:
             casez_tmp =7'h2E;
          7 'b0101111:
             casez_tmp =7'h2F;
          7 'b0110000:
             casez_tmp =7'h30;
          7 'b0110001:
             casez_tmp =7'h31;
          7 'b0110010:
             casez_tmp =7'h32;
          7 'b0110011:
             casez_tmp =7'h33;
          7 'b0110100:
             casez_tmp =7'h34;
          7 'b0110101:
             casez_tmp =7'h35;
          7 'b0110110:
             casez_tmp =7'h36;
          7 'b0110111:
             casez_tmp =7'h37;
          7 'b0111000:
             casez_tmp =7'h38;
          7 'b0111001:
             casez_tmp =7'h39;
          7 'b0111010:
             casez_tmp =7'h3A;
          7 'b0111011:
             casez_tmp =7'h3B;
          7 'b0111100:
             casez_tmp =7'h3C;
          7 'b0111101:
             casez_tmp =7'h3D;
          7 'b0111110:
             casez_tmp =7'h3E;
          7 'b0111111:
             casez_tmp =7'h3F;
          7 'b1000000:
             casez_tmp =7'h40;
          7 'b1000001:
             casez_tmp =7'h41;
          7 'b1000010:
             casez_tmp =7'h42;
          7 'b1000011:
             casez_tmp =7'h43;
          7 'b1000100:
             casez_tmp =7'h44;
          7 'b1000101:
             casez_tmp =7'h45;
          7 'b1000110:
             casez_tmp =7'h46;
          7 'b1000111:
             casez_tmp =7'h47;
          7 'b1001000:
             casez_tmp =7'h48;
          7 'b1001001:
             casez_tmp =7'h49;
          7 'b1001010:
             casez_tmp =7'h4A;
          7 'b1001011:
             casez_tmp =7'h4B;
          7 'b1001100:
             casez_tmp =7'h4C;
          7 'b1001101:
             casez_tmp =7'h4D;
          7 'b1001110:
             casez_tmp =7'h4E;
          7 'b1001111:
             casez_tmp =7'h4F;
          7 'b1010000:
             casez_tmp =7'h50;
          7 'b1010001:
             casez_tmp =7'h51;
          7 'b1010010:
             casez_tmp =7'h52;
          7 'b1010011:
             casez_tmp =7'h53;
          7 'b1010100:
             casez_tmp =7'h54;
          7 'b1010101:
             casez_tmp =7'h55;
          7 'b1010110:
             casez_tmp =7'h56;
          7 'b1010111:
             casez_tmp =7'h57;
          7 'b1011000:
             casez_tmp =7'h58;
          7 'b1011001:
             casez_tmp =7'h59;
          7 'b1011010:
             casez_tmp =7'h5A;
          7 'b1011011:
             casez_tmp =7'h5B;
          7 'b1011100:
             casez_tmp =7'h5C;
          7 'b1011101:
             casez_tmp =7'h5D;
          7 'b1011110:
             casez_tmp =7'h5E;
          7 'b1011111:
             casez_tmp =7'h5F;
          7 'b1100000:
             casez_tmp =7'h60;
          7 'b1100001:
             casez_tmp =7'h61;
          7 'b1100010:
             casez_tmp =7'h62;
          7 'b1100011:
             casez_tmp =7'h63;
          7 'b1100100:
             casez_tmp =7'h64;
          7 'b1100101:
             casez_tmp =7'h65;
          7 'b1100110:
             casez_tmp =7'h66;
          7 'b1100111:
             casez_tmp =7'h67;
          7 'b1101000:
             casez_tmp =7'h68;
          7 'b1101001:
             casez_tmp =7'h69;
          7 'b1101010:
             casez_tmp =7'h6A;
          7 'b1101011:
             casez_tmp =7'h6B;
          7 'b1101100:
             casez_tmp =7'h6C;
          7 'b1101101:
             casez_tmp =7'h6D;
          7 'b1101110:
             casez_tmp =7'h6E;
          7 'b1101111:
             casez_tmp =7'h6F;
          7 'b1110000:
             casez_tmp =7'h70;
          7 'b1110001:
             casez_tmp =7'h71;
          7 'b1110010:
             casez_tmp =7'h72;
          7 'b1110011:
             casez_tmp =7'h73;
          7 'b1110100:
             casez_tmp =7'h74;
          7 'b1110101:
             casez_tmp =7'h75;
          7 'b1110110:
             casez_tmp =7'h76;
          7 'b1110111:
             casez_tmp =7'h77;
          7 'b1111000:
             casez_tmp =7'h78;
          7 'b1111001:
             casez_tmp =7'h79;
          7 'b1111010:
             casez_tmp =7'h7A;
          7 'b1111011:
             casez_tmp =7'h7B;
          7 'b1111100:
             casez_tmp =7'h7C;
          7 'b1111101:
             casez_tmp =7'h7D;
          7 'b1111110:
             casez_tmp =7'h7E;
          default :
             casez_tmp =7'h7F;
         endcase 
       end
  
   wire [17:0] _out_arw_bits_len_T_1=18'h7FF<<auto_in_a_bits_size ;  
   reg casez_tmp_0 ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_source)
          7 'b0000000:
             casez_tmp_0 =count_1;
          7 'b0000001:
             casez_tmp_0 =count_2;
          7 'b0000010:
             casez_tmp_0 =count_3;
          7 'b0000011:
             casez_tmp_0 =count_4;
          7 'b0000100:
             casez_tmp_0 =count_5;
          7 'b0000101:
             casez_tmp_0 =count_6;
          7 'b0000110:
             casez_tmp_0 =count_7;
          7 'b0000111:
             casez_tmp_0 =count_8;
          7 'b0001000:
             casez_tmp_0 =count_9;
          7 'b0001001:
             casez_tmp_0 =count_10;
          7 'b0001010:
             casez_tmp_0 =count_11;
          7 'b0001011:
             casez_tmp_0 =count_12;
          7 'b0001100:
             casez_tmp_0 =count_13;
          7 'b0001101:
             casez_tmp_0 =count_14;
          7 'b0001110:
             casez_tmp_0 =count_15;
          7 'b0001111:
             casez_tmp_0 =count_16;
          7 'b0010000:
             casez_tmp_0 =count_17;
          7 'b0010001:
             casez_tmp_0 =count_18;
          7 'b0010010:
             casez_tmp_0 =count_19;
          7 'b0010011:
             casez_tmp_0 =count_20;
          7 'b0010100:
             casez_tmp_0 =count_21;
          7 'b0010101:
             casez_tmp_0 =count_22;
          7 'b0010110:
             casez_tmp_0 =count_23;
          7 'b0010111:
             casez_tmp_0 =count_24;
          7 'b0011000:
             casez_tmp_0 =count_25;
          7 'b0011001:
             casez_tmp_0 =count_26;
          7 'b0011010:
             casez_tmp_0 =count_27;
          7 'b0011011:
             casez_tmp_0 =count_28;
          7 'b0011100:
             casez_tmp_0 =count_29;
          7 'b0011101:
             casez_tmp_0 =count_30;
          7 'b0011110:
             casez_tmp_0 =count_31;
          7 'b0011111:
             casez_tmp_0 =count_32;
          7 'b0100000:
             casez_tmp_0 =count_33;
          7 'b0100001:
             casez_tmp_0 =count_34;
          7 'b0100010:
             casez_tmp_0 =count_35;
          7 'b0100011:
             casez_tmp_0 =count_36;
          7 'b0100100:
             casez_tmp_0 =count_37;
          7 'b0100101:
             casez_tmp_0 =count_38;
          7 'b0100110:
             casez_tmp_0 =count_39;
          7 'b0100111:
             casez_tmp_0 =count_40;
          7 'b0101000:
             casez_tmp_0 =count_41;
          7 'b0101001:
             casez_tmp_0 =count_42;
          7 'b0101010:
             casez_tmp_0 =count_43;
          7 'b0101011:
             casez_tmp_0 =count_44;
          7 'b0101100:
             casez_tmp_0 =count_45;
          7 'b0101101:
             casez_tmp_0 =count_46;
          7 'b0101110:
             casez_tmp_0 =count_47;
          7 'b0101111:
             casez_tmp_0 =count_48;
          7 'b0110000:
             casez_tmp_0 =count_49;
          7 'b0110001:
             casez_tmp_0 =count_50;
          7 'b0110010:
             casez_tmp_0 =count_51;
          7 'b0110011:
             casez_tmp_0 =count_52;
          7 'b0110100:
             casez_tmp_0 =count_53;
          7 'b0110101:
             casez_tmp_0 =count_54;
          7 'b0110110:
             casez_tmp_0 =count_55;
          7 'b0110111:
             casez_tmp_0 =count_56;
          7 'b0111000:
             casez_tmp_0 =count_57;
          7 'b0111001:
             casez_tmp_0 =count_58;
          7 'b0111010:
             casez_tmp_0 =count_59;
          7 'b0111011:
             casez_tmp_0 =count_60;
          7 'b0111100:
             casez_tmp_0 =count_61;
          7 'b0111101:
             casez_tmp_0 =count_62;
          7 'b0111110:
             casez_tmp_0 =count_63;
          7 'b0111111:
             casez_tmp_0 =count_64;
          7 'b1000000:
             casez_tmp_0 =count_65;
          7 'b1000001:
             casez_tmp_0 =count_66;
          7 'b1000010:
             casez_tmp_0 =count_67;
          7 'b1000011:
             casez_tmp_0 =count_68;
          7 'b1000100:
             casez_tmp_0 =count_69;
          7 'b1000101:
             casez_tmp_0 =count_70;
          7 'b1000110:
             casez_tmp_0 =count_71;
          7 'b1000111:
             casez_tmp_0 =count_72;
          7 'b1001000:
             casez_tmp_0 =count_73;
          7 'b1001001:
             casez_tmp_0 =count_74;
          7 'b1001010:
             casez_tmp_0 =count_75;
          7 'b1001011:
             casez_tmp_0 =count_76;
          7 'b1001100:
             casez_tmp_0 =count_77;
          7 'b1001101:
             casez_tmp_0 =count_78;
          7 'b1001110:
             casez_tmp_0 =count_79;
          7 'b1001111:
             casez_tmp_0 =count_80;
          7 'b1010000:
             casez_tmp_0 =count_81;
          7 'b1010001:
             casez_tmp_0 =count_82;
          7 'b1010010:
             casez_tmp_0 =count_83;
          7 'b1010011:
             casez_tmp_0 =count_84;
          7 'b1010100:
             casez_tmp_0 =count_85;
          7 'b1010101:
             casez_tmp_0 =count_86;
          7 'b1010110:
             casez_tmp_0 =count_87;
          7 'b1010111:
             casez_tmp_0 =count_88;
          7 'b1011000:
             casez_tmp_0 =count_89;
          7 'b1011001:
             casez_tmp_0 =count_90;
          7 'b1011010:
             casez_tmp_0 =count_91;
          7 'b1011011:
             casez_tmp_0 =count_92;
          7 'b1011100:
             casez_tmp_0 =count_93;
          7 'b1011101:
             casez_tmp_0 =count_94;
          7 'b1011110:
             casez_tmp_0 =count_95;
          7 'b1011111:
             casez_tmp_0 =count_96;
          7 'b1100000:
             casez_tmp_0 =count_97;
          7 'b1100001:
             casez_tmp_0 =count_98;
          7 'b1100010:
             casez_tmp_0 =count_99;
          7 'b1100011:
             casez_tmp_0 =count_100;
          7 'b1100100:
             casez_tmp_0 =count_101;
          7 'b1100101:
             casez_tmp_0 =count_102;
          7 'b1100110:
             casez_tmp_0 =count_103;
          7 'b1100111:
             casez_tmp_0 =count_104;
          7 'b1101000:
             casez_tmp_0 =count_105;
          7 'b1101001:
             casez_tmp_0 =count_106;
          7 'b1101010:
             casez_tmp_0 =count_107;
          7 'b1101011:
             casez_tmp_0 =count_108;
          7 'b1101100:
             casez_tmp_0 =count_109;
          7 'b1101101:
             casez_tmp_0 =count_110;
          7 'b1101110:
             casez_tmp_0 =count_111;
          7 'b1101111:
             casez_tmp_0 =count_112;
          7 'b1110000:
             casez_tmp_0 =count_113;
          7 'b1110001:
             casez_tmp_0 =count_114;
          7 'b1110010:
             casez_tmp_0 =count_115;
          7 'b1110011:
             casez_tmp_0 =count_116;
          7 'b1110100:
             casez_tmp_0 =count_117;
          7 'b1110101:
             casez_tmp_0 =count_118;
          7 'b1110110:
             casez_tmp_0 =count_119;
          7 'b1110111:
             casez_tmp_0 =count_120;
          7 'b1111000:
             casez_tmp_0 =count_121;
          7 'b1111001:
             casez_tmp_0 =count_122;
          7 'b1111010:
             casez_tmp_0 =count_123;
          7 'b1111011:
             casez_tmp_0 =count_124;
          7 'b1111100:
             casez_tmp_0 =count_125;
          7 'b1111101:
             casez_tmp_0 =count_126;
          7 'b1111110:
             casez_tmp_0 =count_127;
          default :
             casez_tmp_0 =count_128;
         endcase 
       end
  
   wire stall=casez_tmp_0&a_first ;  
   wire _out_w_valid_T_3=doneAW|_queue_arw_deq_q_io_enq_ready ;  
   wire nodeIn_a_ready=~stall&(auto_in_a_bits_opcode[2] ? _queue_arw_deq_q_io_enq_ready:_out_w_valid_T_3&_nodeOut_w_deq_q_io_enq_ready) ;  
   wire out_arw_valid=~stall&auto_in_a_valid&(auto_in_a_bits_opcode[2]|~doneAW&_nodeOut_w_deq_q_io_enq_ready) ;  
   reg r_holds_d ;  
   reg [2:0] b_delay ;  
   wire r_wins=auto_out_r_valid&b_delay!=3'h7|r_holds_d ;  
   wire nodeOut_r_ready=auto_in_d_ready&r_wins ;  
   wire nodeOut_b_ready=auto_in_d_ready&~r_wins ;  
   wire nodeIn_d_valid=r_wins ? auto_out_r_valid:auto_out_b_valid ;  
   reg r_first ;  
   reg r_denied_r ;  
   wire r_denied=r_first ? (&auto_out_r_bits_resp):r_denied_r ;  
   wire [2:0] nodeIn_d_bits_opcode={2'h0,r_wins} ;  
   wire [2:0] nodeIn_d_bits_size=r_wins ? auto_out_r_bits_echo_tl_state_size[2:0]:auto_out_b_bits_echo_tl_state_size[2:0] ;  
   wire [6:0] nodeIn_d_bits_source=r_wins ? auto_out_r_bits_echo_tl_state_source:auto_out_b_bits_echo_tl_state_source ;  
   wire nodeIn_d_bits_denied=r_wins ? r_denied:(|auto_out_b_bits_resp) ;  
   wire nodeIn_d_bits_corrupt=r_wins&((|auto_out_r_bits_resp)|r_denied) ;  
   wire [6:0] d_sel_shiftAmount=r_wins ? auto_out_r_bits_id:auto_out_b_bits_id ;  
   wire d_last=~r_wins|auto_out_r_bits_last ;  
   wire _inc_T_127=_queue_arw_deq_q_io_enq_ready&out_arw_valid ;  
   wire inc=casez_tmp==7'h0&_inc_T_127 ;  
   wire _dec_T_255=auto_in_d_ready&nodeIn_d_valid ;  
   wire dec=d_sel_shiftAmount==7'h0&d_last&_dec_T_255 ;  
   wire inc_1=casez_tmp==7'h1&_inc_T_127 ;  
   wire dec_1=d_sel_shiftAmount==7'h1&d_last&_dec_T_255 ;  
   wire inc_2=casez_tmp==7'h2&_inc_T_127 ;  
   wire dec_2=d_sel_shiftAmount==7'h2&d_last&_dec_T_255 ;  
   wire inc_3=casez_tmp==7'h3&_inc_T_127 ;  
   wire dec_3=d_sel_shiftAmount==7'h3&d_last&_dec_T_255 ;  
   wire inc_4=casez_tmp==7'h4&_inc_T_127 ;  
   wire dec_4=d_sel_shiftAmount==7'h4&d_last&_dec_T_255 ;  
   wire inc_5=casez_tmp==7'h5&_inc_T_127 ;  
   wire dec_5=d_sel_shiftAmount==7'h5&d_last&_dec_T_255 ;  
   wire inc_6=casez_tmp==7'h6&_inc_T_127 ;  
   wire dec_6=d_sel_shiftAmount==7'h6&d_last&_dec_T_255 ;  
   wire inc_7=casez_tmp==7'h7&_inc_T_127 ;  
   wire dec_7=d_sel_shiftAmount==7'h7&d_last&_dec_T_255 ;  
   wire inc_8=casez_tmp==7'h8&_inc_T_127 ;  
   wire dec_8=d_sel_shiftAmount==7'h8&d_last&_dec_T_255 ;  
   wire inc_9=casez_tmp==7'h9&_inc_T_127 ;  
   wire dec_9=d_sel_shiftAmount==7'h9&d_last&_dec_T_255 ;  
   wire inc_10=casez_tmp==7'hA&_inc_T_127 ;  
   wire dec_10=d_sel_shiftAmount==7'hA&d_last&_dec_T_255 ;  
   wire inc_11=casez_tmp==7'hB&_inc_T_127 ;  
   wire dec_11=d_sel_shiftAmount==7'hB&d_last&_dec_T_255 ;  
   wire inc_12=casez_tmp==7'hC&_inc_T_127 ;  
   wire dec_12=d_sel_shiftAmount==7'hC&d_last&_dec_T_255 ;  
   wire inc_13=casez_tmp==7'hD&_inc_T_127 ;  
   wire dec_13=d_sel_shiftAmount==7'hD&d_last&_dec_T_255 ;  
   wire inc_14=casez_tmp==7'hE&_inc_T_127 ;  
   wire dec_14=d_sel_shiftAmount==7'hE&d_last&_dec_T_255 ;  
   wire inc_15=casez_tmp==7'hF&_inc_T_127 ;  
   wire dec_15=d_sel_shiftAmount==7'hF&d_last&_dec_T_255 ;  
   wire inc_16=casez_tmp==7'h10&_inc_T_127 ;  
   wire dec_16=d_sel_shiftAmount==7'h10&d_last&_dec_T_255 ;  
   wire inc_17=casez_tmp==7'h11&_inc_T_127 ;  
   wire dec_17=d_sel_shiftAmount==7'h11&d_last&_dec_T_255 ;  
   wire inc_18=casez_tmp==7'h12&_inc_T_127 ;  
   wire dec_18=d_sel_shiftAmount==7'h12&d_last&_dec_T_255 ;  
   wire inc_19=casez_tmp==7'h13&_inc_T_127 ;  
   wire dec_19=d_sel_shiftAmount==7'h13&d_last&_dec_T_255 ;  
   wire inc_20=casez_tmp==7'h14&_inc_T_127 ;  
   wire dec_20=d_sel_shiftAmount==7'h14&d_last&_dec_T_255 ;  
   wire inc_21=casez_tmp==7'h15&_inc_T_127 ;  
   wire dec_21=d_sel_shiftAmount==7'h15&d_last&_dec_T_255 ;  
   wire inc_22=casez_tmp==7'h16&_inc_T_127 ;  
   wire dec_22=d_sel_shiftAmount==7'h16&d_last&_dec_T_255 ;  
   wire inc_23=casez_tmp==7'h17&_inc_T_127 ;  
   wire dec_23=d_sel_shiftAmount==7'h17&d_last&_dec_T_255 ;  
   wire inc_24=casez_tmp==7'h18&_inc_T_127 ;  
   wire dec_24=d_sel_shiftAmount==7'h18&d_last&_dec_T_255 ;  
   wire inc_25=casez_tmp==7'h19&_inc_T_127 ;  
   wire dec_25=d_sel_shiftAmount==7'h19&d_last&_dec_T_255 ;  
   wire inc_26=casez_tmp==7'h1A&_inc_T_127 ;  
   wire dec_26=d_sel_shiftAmount==7'h1A&d_last&_dec_T_255 ;  
   wire inc_27=casez_tmp==7'h1B&_inc_T_127 ;  
   wire dec_27=d_sel_shiftAmount==7'h1B&d_last&_dec_T_255 ;  
   wire inc_28=casez_tmp==7'h1C&_inc_T_127 ;  
   wire dec_28=d_sel_shiftAmount==7'h1C&d_last&_dec_T_255 ;  
   wire inc_29=casez_tmp==7'h1D&_inc_T_127 ;  
   wire dec_29=d_sel_shiftAmount==7'h1D&d_last&_dec_T_255 ;  
   wire inc_30=casez_tmp==7'h1E&_inc_T_127 ;  
   wire dec_30=d_sel_shiftAmount==7'h1E&d_last&_dec_T_255 ;  
   wire inc_31=casez_tmp==7'h1F&_inc_T_127 ;  
   wire dec_31=d_sel_shiftAmount==7'h1F&d_last&_dec_T_255 ;  
   wire inc_32=casez_tmp==7'h20&_inc_T_127 ;  
   wire dec_32=d_sel_shiftAmount==7'h20&d_last&_dec_T_255 ;  
   wire inc_33=casez_tmp==7'h21&_inc_T_127 ;  
   wire dec_33=d_sel_shiftAmount==7'h21&d_last&_dec_T_255 ;  
   wire inc_34=casez_tmp==7'h22&_inc_T_127 ;  
   wire dec_34=d_sel_shiftAmount==7'h22&d_last&_dec_T_255 ;  
   wire inc_35=casez_tmp==7'h23&_inc_T_127 ;  
   wire dec_35=d_sel_shiftAmount==7'h23&d_last&_dec_T_255 ;  
   wire inc_36=casez_tmp==7'h24&_inc_T_127 ;  
   wire dec_36=d_sel_shiftAmount==7'h24&d_last&_dec_T_255 ;  
   wire inc_37=casez_tmp==7'h25&_inc_T_127 ;  
   wire dec_37=d_sel_shiftAmount==7'h25&d_last&_dec_T_255 ;  
   wire inc_38=casez_tmp==7'h26&_inc_T_127 ;  
   wire dec_38=d_sel_shiftAmount==7'h26&d_last&_dec_T_255 ;  
   wire inc_39=casez_tmp==7'h27&_inc_T_127 ;  
   wire dec_39=d_sel_shiftAmount==7'h27&d_last&_dec_T_255 ;  
   wire inc_40=casez_tmp==7'h28&_inc_T_127 ;  
   wire dec_40=d_sel_shiftAmount==7'h28&d_last&_dec_T_255 ;  
   wire inc_41=casez_tmp==7'h29&_inc_T_127 ;  
   wire dec_41=d_sel_shiftAmount==7'h29&d_last&_dec_T_255 ;  
   wire inc_42=casez_tmp==7'h2A&_inc_T_127 ;  
   wire dec_42=d_sel_shiftAmount==7'h2A&d_last&_dec_T_255 ;  
   wire inc_43=casez_tmp==7'h2B&_inc_T_127 ;  
   wire dec_43=d_sel_shiftAmount==7'h2B&d_last&_dec_T_255 ;  
   wire inc_44=casez_tmp==7'h2C&_inc_T_127 ;  
   wire dec_44=d_sel_shiftAmount==7'h2C&d_last&_dec_T_255 ;  
   wire inc_45=casez_tmp==7'h2D&_inc_T_127 ;  
   wire dec_45=d_sel_shiftAmount==7'h2D&d_last&_dec_T_255 ;  
   wire inc_46=casez_tmp==7'h2E&_inc_T_127 ;  
   wire dec_46=d_sel_shiftAmount==7'h2E&d_last&_dec_T_255 ;  
   wire inc_47=casez_tmp==7'h2F&_inc_T_127 ;  
   wire dec_47=d_sel_shiftAmount==7'h2F&d_last&_dec_T_255 ;  
   wire inc_48=casez_tmp==7'h30&_inc_T_127 ;  
   wire dec_48=d_sel_shiftAmount==7'h30&d_last&_dec_T_255 ;  
   wire inc_49=casez_tmp==7'h31&_inc_T_127 ;  
   wire dec_49=d_sel_shiftAmount==7'h31&d_last&_dec_T_255 ;  
   wire inc_50=casez_tmp==7'h32&_inc_T_127 ;  
   wire dec_50=d_sel_shiftAmount==7'h32&d_last&_dec_T_255 ;  
   wire inc_51=casez_tmp==7'h33&_inc_T_127 ;  
   wire dec_51=d_sel_shiftAmount==7'h33&d_last&_dec_T_255 ;  
   wire inc_52=casez_tmp==7'h34&_inc_T_127 ;  
   wire dec_52=d_sel_shiftAmount==7'h34&d_last&_dec_T_255 ;  
   wire inc_53=casez_tmp==7'h35&_inc_T_127 ;  
   wire dec_53=d_sel_shiftAmount==7'h35&d_last&_dec_T_255 ;  
   wire inc_54=casez_tmp==7'h36&_inc_T_127 ;  
   wire dec_54=d_sel_shiftAmount==7'h36&d_last&_dec_T_255 ;  
   wire inc_55=casez_tmp==7'h37&_inc_T_127 ;  
   wire dec_55=d_sel_shiftAmount==7'h37&d_last&_dec_T_255 ;  
   wire inc_56=casez_tmp==7'h38&_inc_T_127 ;  
   wire dec_56=d_sel_shiftAmount==7'h38&d_last&_dec_T_255 ;  
   wire inc_57=casez_tmp==7'h39&_inc_T_127 ;  
   wire dec_57=d_sel_shiftAmount==7'h39&d_last&_dec_T_255 ;  
   wire inc_58=casez_tmp==7'h3A&_inc_T_127 ;  
   wire dec_58=d_sel_shiftAmount==7'h3A&d_last&_dec_T_255 ;  
   wire inc_59=casez_tmp==7'h3B&_inc_T_127 ;  
   wire dec_59=d_sel_shiftAmount==7'h3B&d_last&_dec_T_255 ;  
   wire inc_60=casez_tmp==7'h3C&_inc_T_127 ;  
   wire dec_60=d_sel_shiftAmount==7'h3C&d_last&_dec_T_255 ;  
   wire inc_61=casez_tmp==7'h3D&_inc_T_127 ;  
   wire dec_61=d_sel_shiftAmount==7'h3D&d_last&_dec_T_255 ;  
   wire inc_62=casez_tmp==7'h3E&_inc_T_127 ;  
   wire dec_62=d_sel_shiftAmount==7'h3E&d_last&_dec_T_255 ;  
   wire inc_63=casez_tmp==7'h3F&_inc_T_127 ;  
   wire dec_63=d_sel_shiftAmount==7'h3F&d_last&_dec_T_255 ;  
   wire inc_64=casez_tmp==7'h40&_inc_T_127 ;  
   wire dec_64=d_sel_shiftAmount==7'h40&d_last&_dec_T_255 ;  
   wire inc_65=casez_tmp==7'h41&_inc_T_127 ;  
   wire dec_65=d_sel_shiftAmount==7'h41&d_last&_dec_T_255 ;  
   wire inc_66=casez_tmp==7'h42&_inc_T_127 ;  
   wire dec_66=d_sel_shiftAmount==7'h42&d_last&_dec_T_255 ;  
   wire inc_67=casez_tmp==7'h43&_inc_T_127 ;  
   wire dec_67=d_sel_shiftAmount==7'h43&d_last&_dec_T_255 ;  
   wire inc_68=casez_tmp==7'h44&_inc_T_127 ;  
   wire dec_68=d_sel_shiftAmount==7'h44&d_last&_dec_T_255 ;  
   wire inc_69=casez_tmp==7'h45&_inc_T_127 ;  
   wire dec_69=d_sel_shiftAmount==7'h45&d_last&_dec_T_255 ;  
   wire inc_70=casez_tmp==7'h46&_inc_T_127 ;  
   wire dec_70=d_sel_shiftAmount==7'h46&d_last&_dec_T_255 ;  
   wire inc_71=casez_tmp==7'h47&_inc_T_127 ;  
   wire dec_71=d_sel_shiftAmount==7'h47&d_last&_dec_T_255 ;  
   wire inc_72=casez_tmp==7'h48&_inc_T_127 ;  
   wire dec_72=d_sel_shiftAmount==7'h48&d_last&_dec_T_255 ;  
   wire inc_73=casez_tmp==7'h49&_inc_T_127 ;  
   wire dec_73=d_sel_shiftAmount==7'h49&d_last&_dec_T_255 ;  
   wire inc_74=casez_tmp==7'h4A&_inc_T_127 ;  
   wire dec_74=d_sel_shiftAmount==7'h4A&d_last&_dec_T_255 ;  
   wire inc_75=casez_tmp==7'h4B&_inc_T_127 ;  
   wire dec_75=d_sel_shiftAmount==7'h4B&d_last&_dec_T_255 ;  
   wire inc_76=casez_tmp==7'h4C&_inc_T_127 ;  
   wire dec_76=d_sel_shiftAmount==7'h4C&d_last&_dec_T_255 ;  
   wire inc_77=casez_tmp==7'h4D&_inc_T_127 ;  
   wire dec_77=d_sel_shiftAmount==7'h4D&d_last&_dec_T_255 ;  
   wire inc_78=casez_tmp==7'h4E&_inc_T_127 ;  
   wire dec_78=d_sel_shiftAmount==7'h4E&d_last&_dec_T_255 ;  
   wire inc_79=casez_tmp==7'h4F&_inc_T_127 ;  
   wire dec_79=d_sel_shiftAmount==7'h4F&d_last&_dec_T_255 ;  
   wire inc_80=casez_tmp==7'h50&_inc_T_127 ;  
   wire dec_80=d_sel_shiftAmount==7'h50&d_last&_dec_T_255 ;  
   wire inc_81=casez_tmp==7'h51&_inc_T_127 ;  
   wire dec_81=d_sel_shiftAmount==7'h51&d_last&_dec_T_255 ;  
   wire inc_82=casez_tmp==7'h52&_inc_T_127 ;  
   wire dec_82=d_sel_shiftAmount==7'h52&d_last&_dec_T_255 ;  
   wire inc_83=casez_tmp==7'h53&_inc_T_127 ;  
   wire dec_83=d_sel_shiftAmount==7'h53&d_last&_dec_T_255 ;  
   wire inc_84=casez_tmp==7'h54&_inc_T_127 ;  
   wire dec_84=d_sel_shiftAmount==7'h54&d_last&_dec_T_255 ;  
   wire inc_85=casez_tmp==7'h55&_inc_T_127 ;  
   wire dec_85=d_sel_shiftAmount==7'h55&d_last&_dec_T_255 ;  
   wire inc_86=casez_tmp==7'h56&_inc_T_127 ;  
   wire dec_86=d_sel_shiftAmount==7'h56&d_last&_dec_T_255 ;  
   wire inc_87=casez_tmp==7'h57&_inc_T_127 ;  
   wire dec_87=d_sel_shiftAmount==7'h57&d_last&_dec_T_255 ;  
   wire inc_88=casez_tmp==7'h58&_inc_T_127 ;  
   wire dec_88=d_sel_shiftAmount==7'h58&d_last&_dec_T_255 ;  
   wire inc_89=casez_tmp==7'h59&_inc_T_127 ;  
   wire dec_89=d_sel_shiftAmount==7'h59&d_last&_dec_T_255 ;  
   wire inc_90=casez_tmp==7'h5A&_inc_T_127 ;  
   wire dec_90=d_sel_shiftAmount==7'h5A&d_last&_dec_T_255 ;  
   wire inc_91=casez_tmp==7'h5B&_inc_T_127 ;  
   wire dec_91=d_sel_shiftAmount==7'h5B&d_last&_dec_T_255 ;  
   wire inc_92=casez_tmp==7'h5C&_inc_T_127 ;  
   wire dec_92=d_sel_shiftAmount==7'h5C&d_last&_dec_T_255 ;  
   wire inc_93=casez_tmp==7'h5D&_inc_T_127 ;  
   wire dec_93=d_sel_shiftAmount==7'h5D&d_last&_dec_T_255 ;  
   wire inc_94=casez_tmp==7'h5E&_inc_T_127 ;  
   wire dec_94=d_sel_shiftAmount==7'h5E&d_last&_dec_T_255 ;  
   wire inc_95=casez_tmp==7'h5F&_inc_T_127 ;  
   wire dec_95=d_sel_shiftAmount==7'h5F&d_last&_dec_T_255 ;  
   wire inc_96=casez_tmp==7'h60&_inc_T_127 ;  
   wire dec_96=d_sel_shiftAmount==7'h60&d_last&_dec_T_255 ;  
   wire inc_97=casez_tmp==7'h61&_inc_T_127 ;  
   wire dec_97=d_sel_shiftAmount==7'h61&d_last&_dec_T_255 ;  
   wire inc_98=casez_tmp==7'h62&_inc_T_127 ;  
   wire dec_98=d_sel_shiftAmount==7'h62&d_last&_dec_T_255 ;  
   wire inc_99=casez_tmp==7'h63&_inc_T_127 ;  
   wire dec_99=d_sel_shiftAmount==7'h63&d_last&_dec_T_255 ;  
   wire inc_100=casez_tmp==7'h64&_inc_T_127 ;  
   wire dec_100=d_sel_shiftAmount==7'h64&d_last&_dec_T_255 ;  
   wire inc_101=casez_tmp==7'h65&_inc_T_127 ;  
   wire dec_101=d_sel_shiftAmount==7'h65&d_last&_dec_T_255 ;  
   wire inc_102=casez_tmp==7'h66&_inc_T_127 ;  
   wire dec_102=d_sel_shiftAmount==7'h66&d_last&_dec_T_255 ;  
   wire inc_103=casez_tmp==7'h67&_inc_T_127 ;  
   wire dec_103=d_sel_shiftAmount==7'h67&d_last&_dec_T_255 ;  
   wire inc_104=casez_tmp==7'h68&_inc_T_127 ;  
   wire dec_104=d_sel_shiftAmount==7'h68&d_last&_dec_T_255 ;  
   wire inc_105=casez_tmp==7'h69&_inc_T_127 ;  
   wire dec_105=d_sel_shiftAmount==7'h69&d_last&_dec_T_255 ;  
   wire inc_106=casez_tmp==7'h6A&_inc_T_127 ;  
   wire dec_106=d_sel_shiftAmount==7'h6A&d_last&_dec_T_255 ;  
   wire inc_107=casez_tmp==7'h6B&_inc_T_127 ;  
   wire dec_107=d_sel_shiftAmount==7'h6B&d_last&_dec_T_255 ;  
   wire inc_108=casez_tmp==7'h6C&_inc_T_127 ;  
   wire dec_108=d_sel_shiftAmount==7'h6C&d_last&_dec_T_255 ;  
   wire inc_109=casez_tmp==7'h6D&_inc_T_127 ;  
   wire dec_109=d_sel_shiftAmount==7'h6D&d_last&_dec_T_255 ;  
   wire inc_110=casez_tmp==7'h6E&_inc_T_127 ;  
   wire dec_110=d_sel_shiftAmount==7'h6E&d_last&_dec_T_255 ;  
   wire inc_111=casez_tmp==7'h6F&_inc_T_127 ;  
   wire dec_111=d_sel_shiftAmount==7'h6F&d_last&_dec_T_255 ;  
   wire inc_112=casez_tmp==7'h70&_inc_T_127 ;  
   wire dec_112=d_sel_shiftAmount==7'h70&d_last&_dec_T_255 ;  
   wire inc_113=casez_tmp==7'h71&_inc_T_127 ;  
   wire dec_113=d_sel_shiftAmount==7'h71&d_last&_dec_T_255 ;  
   wire inc_114=casez_tmp==7'h72&_inc_T_127 ;  
   wire dec_114=d_sel_shiftAmount==7'h72&d_last&_dec_T_255 ;  
   wire inc_115=casez_tmp==7'h73&_inc_T_127 ;  
   wire dec_115=d_sel_shiftAmount==7'h73&d_last&_dec_T_255 ;  
   wire inc_116=casez_tmp==7'h74&_inc_T_127 ;  
   wire dec_116=d_sel_shiftAmount==7'h74&d_last&_dec_T_255 ;  
   wire inc_117=casez_tmp==7'h75&_inc_T_127 ;  
   wire dec_117=d_sel_shiftAmount==7'h75&d_last&_dec_T_255 ;  
   wire inc_118=casez_tmp==7'h76&_inc_T_127 ;  
   wire dec_118=d_sel_shiftAmount==7'h76&d_last&_dec_T_255 ;  
   wire inc_119=casez_tmp==7'h77&_inc_T_127 ;  
   wire dec_119=d_sel_shiftAmount==7'h77&d_last&_dec_T_255 ;  
   wire inc_120=casez_tmp==7'h78&_inc_T_127 ;  
   wire dec_120=d_sel_shiftAmount==7'h78&d_last&_dec_T_255 ;  
   wire inc_121=casez_tmp==7'h79&_inc_T_127 ;  
   wire dec_121=d_sel_shiftAmount==7'h79&d_last&_dec_T_255 ;  
   wire inc_122=casez_tmp==7'h7A&_inc_T_127 ;  
   wire dec_122=d_sel_shiftAmount==7'h7A&d_last&_dec_T_255 ;  
   wire inc_123=casez_tmp==7'h7B&_inc_T_127 ;  
   wire dec_123=d_sel_shiftAmount==7'h7B&d_last&_dec_T_255 ;  
   wire inc_124=casez_tmp==7'h7C&_inc_T_127 ;  
   wire dec_124=d_sel_shiftAmount==7'h7C&d_last&_dec_T_255 ;  
   wire inc_125=casez_tmp==7'h7D&_inc_T_127 ;  
   wire dec_125=d_sel_shiftAmount==7'h7D&d_last&_dec_T_255 ;  
   wire inc_126=casez_tmp==7'h7E&_inc_T_127 ;  
   wire dec_126=d_sel_shiftAmount==7'h7E&d_last&_dec_T_255 ;  
   wire inc_127=(&casez_tmp)&_inc_T_127 ;  
   wire dec_127=(&d_sel_shiftAmount)&d_last&_dec_T_255 ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~dec|count_1))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc|~count_1))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_1|count_2))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_1|~count_2))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_2|count_3))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_2|~count_3))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_3|count_4))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_3|~count_4))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_4|count_5))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_4|~count_5))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_5|count_6))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_5|~count_6))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_6|count_7))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_6|~count_7))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_7|count_8))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_7|~count_8))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_8|count_9))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_8|~count_9))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_9|count_10))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_9|~count_10))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_10|count_11))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_10|~count_11))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_11|count_12))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_11|~count_12))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_12|count_13))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_12|~count_13))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_13|count_14))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_13|~count_14))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_14|count_15))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_14|~count_15))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_15|count_16))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_15|~count_16))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_16|count_17))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_16|~count_17))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_17|count_18))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_17|~count_18))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_18|count_19))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_18|~count_19))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_19|count_20))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_19|~count_20))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_20|count_21))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_20|~count_21))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_21|count_22))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_21|~count_22))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_22|count_23))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_22|~count_23))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_23|count_24))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_23|~count_24))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_24|count_25))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_24|~count_25))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_25|count_26))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_25|~count_26))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_26|count_27))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_26|~count_27))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_27|count_28))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_27|~count_28))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_28|count_29))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_28|~count_29))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_29|count_30))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_29|~count_30))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_30|count_31))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_30|~count_31))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_31|count_32))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_31|~count_32))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_32|count_33))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_32|~count_33))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_33|count_34))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_33|~count_34))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_34|count_35))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_34|~count_35))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_35|count_36))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_35|~count_36))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_36|count_37))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_36|~count_37))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_37|count_38))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_37|~count_38))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_38|count_39))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_38|~count_39))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_39|count_40))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_39|~count_40))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_40|count_41))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_40|~count_41))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_41|count_42))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_41|~count_42))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_42|count_43))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_42|~count_43))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_43|count_44))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_43|~count_44))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_44|count_45))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_44|~count_45))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_45|count_46))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_45|~count_46))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_46|count_47))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_46|~count_47))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_47|count_48))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_47|~count_48))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_48|count_49))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_48|~count_49))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_49|count_50))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_49|~count_50))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_50|count_51))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_50|~count_51))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_51|count_52))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_51|~count_52))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_52|count_53))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_52|~count_53))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_53|count_54))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_53|~count_54))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_54|count_55))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_54|~count_55))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_55|count_56))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_55|~count_56))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_56|count_57))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_56|~count_57))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_57|count_58))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_57|~count_58))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_58|count_59))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_58|~count_59))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_59|count_60))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_59|~count_60))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_60|count_61))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_60|~count_61))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_61|count_62))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_61|~count_62))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_62|count_63))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_62|~count_63))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_63|count_64))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_63|~count_64))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_64|count_65))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_64|~count_65))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_65|count_66))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_65|~count_66))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_66|count_67))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_66|~count_67))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_67|count_68))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_67|~count_68))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_68|count_69))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_68|~count_69))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_69|count_70))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_69|~count_70))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_70|count_71))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_70|~count_71))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_71|count_72))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_71|~count_72))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_72|count_73))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_72|~count_73))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_73|count_74))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_73|~count_74))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_74|count_75))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_74|~count_75))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_75|count_76))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_75|~count_76))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_76|count_77))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_76|~count_77))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_77|count_78))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_77|~count_78))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_78|count_79))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_78|~count_79))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_79|count_80))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_79|~count_80))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_80|count_81))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_80|~count_81))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_81|count_82))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_81|~count_82))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_82|count_83))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_82|~count_83))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_83|count_84))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_83|~count_84))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_84|count_85))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_84|~count_85))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_85|count_86))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_85|~count_86))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_86|count_87))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_86|~count_87))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_87|count_88))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_87|~count_88))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_88|count_89))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_88|~count_89))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_89|count_90))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_89|~count_90))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_90|count_91))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_90|~count_91))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_91|count_92))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_91|~count_92))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_92|count_93))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_92|~count_93))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_93|count_94))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_93|~count_94))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_94|count_95))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_94|~count_95))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_95|count_96))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_95|~count_96))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_96|count_97))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_96|~count_97))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_97|count_98))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_97|~count_98))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_98|count_99))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_98|~count_99))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_99|count_100))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_99|~count_100))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_100|count_101))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_100|~count_101))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_101|count_102))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_101|~count_102))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_102|count_103))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_102|~count_103))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_103|count_104))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_103|~count_104))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_104|count_105))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_104|~count_105))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_105|count_106))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_105|~count_106))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_106|count_107))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_106|~count_107))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_107|count_108))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_107|~count_108))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_108|count_109))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_108|~count_109))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_109|count_110))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_109|~count_110))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_110|count_111))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_110|~count_111))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_111|count_112))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_111|~count_112))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_112|count_113))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_112|~count_113))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_113|count_114))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_113|~count_114))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_114|count_115))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_114|~count_115))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_115|count_116))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_115|~count_116))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_116|count_117))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_116|~count_117))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_117|count_118))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_117|~count_118))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_118|count_119))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_118|~count_119))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_119|count_120))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_119|~count_120))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_120|count_121))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_120|~count_121))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_121|count_122))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_121|~count_122))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_122|count_123))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_122|~count_123))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_123|count_124))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_123|~count_124))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_124|count_125))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_124|~count_125))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_125|count_126))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_125|~count_126))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_126|count_127))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_126|~count_127))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~dec_127|count_128))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:273 assert (!dec || count =/= 0.U)        // underflow\n");
              if (1)$display("");
            end 
         if (~reset&~(~inc_127|~count_128))
            begin 
              if (1)$display("Assertion failed\n    at ToAXI4.scala:274 assert (!inc || count =/= maxCount.U) // overflow\n");
              if (1)$display("");
            end 
       end
  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              counter <=3'h0;
              doneAW <=1'h0;
              r_holds_d <=1'h0;
              r_first <=1'h1;
              count_1 <=1'h0;
              count_2 <=1'h0;
              count_3 <=1'h0;
              count_4 <=1'h0;
              count_5 <=1'h0;
              count_6 <=1'h0;
              count_7 <=1'h0;
              count_8 <=1'h0;
              count_9 <=1'h0;
              count_10 <=1'h0;
              count_11 <=1'h0;
              count_12 <=1'h0;
              count_13 <=1'h0;
              count_14 <=1'h0;
              count_15 <=1'h0;
              count_16 <=1'h0;
              count_17 <=1'h0;
              count_18 <=1'h0;
              count_19 <=1'h0;
              count_20 <=1'h0;
              count_21 <=1'h0;
              count_22 <=1'h0;
              count_23 <=1'h0;
              count_24 <=1'h0;
              count_25 <=1'h0;
              count_26 <=1'h0;
              count_27 <=1'h0;
              count_28 <=1'h0;
              count_29 <=1'h0;
              count_30 <=1'h0;
              count_31 <=1'h0;
              count_32 <=1'h0;
              count_33 <=1'h0;
              count_34 <=1'h0;
              count_35 <=1'h0;
              count_36 <=1'h0;
              count_37 <=1'h0;
              count_38 <=1'h0;
              count_39 <=1'h0;
              count_40 <=1'h0;
              count_41 <=1'h0;
              count_42 <=1'h0;
              count_43 <=1'h0;
              count_44 <=1'h0;
              count_45 <=1'h0;
              count_46 <=1'h0;
              count_47 <=1'h0;
              count_48 <=1'h0;
              count_49 <=1'h0;
              count_50 <=1'h0;
              count_51 <=1'h0;
              count_52 <=1'h0;
              count_53 <=1'h0;
              count_54 <=1'h0;
              count_55 <=1'h0;
              count_56 <=1'h0;
              count_57 <=1'h0;
              count_58 <=1'h0;
              count_59 <=1'h0;
              count_60 <=1'h0;
              count_61 <=1'h0;
              count_62 <=1'h0;
              count_63 <=1'h0;
              count_64 <=1'h0;
              count_65 <=1'h0;
              count_66 <=1'h0;
              count_67 <=1'h0;
              count_68 <=1'h0;
              count_69 <=1'h0;
              count_70 <=1'h0;
              count_71 <=1'h0;
              count_72 <=1'h0;
              count_73 <=1'h0;
              count_74 <=1'h0;
              count_75 <=1'h0;
              count_76 <=1'h0;
              count_77 <=1'h0;
              count_78 <=1'h0;
              count_79 <=1'h0;
              count_80 <=1'h0;
              count_81 <=1'h0;
              count_82 <=1'h0;
              count_83 <=1'h0;
              count_84 <=1'h0;
              count_85 <=1'h0;
              count_86 <=1'h0;
              count_87 <=1'h0;
              count_88 <=1'h0;
              count_89 <=1'h0;
              count_90 <=1'h0;
              count_91 <=1'h0;
              count_92 <=1'h0;
              count_93 <=1'h0;
              count_94 <=1'h0;
              count_95 <=1'h0;
              count_96 <=1'h0;
              count_97 <=1'h0;
              count_98 <=1'h0;
              count_99 <=1'h0;
              count_100 <=1'h0;
              count_101 <=1'h0;
              count_102 <=1'h0;
              count_103 <=1'h0;
              count_104 <=1'h0;
              count_105 <=1'h0;
              count_106 <=1'h0;
              count_107 <=1'h0;
              count_108 <=1'h0;
              count_109 <=1'h0;
              count_110 <=1'h0;
              count_111 <=1'h0;
              count_112 <=1'h0;
              count_113 <=1'h0;
              count_114 <=1'h0;
              count_115 <=1'h0;
              count_116 <=1'h0;
              count_117 <=1'h0;
              count_118 <=1'h0;
              count_119 <=1'h0;
              count_120 <=1'h0;
              count_121 <=1'h0;
              count_122 <=1'h0;
              count_123 <=1'h0;
              count_124 <=1'h0;
              count_125 <=1'h0;
              count_126 <=1'h0;
              count_127 <=1'h0;
              count_128 <=1'h0;
            end 
          else 
            begin 
              if (nodeIn_a_ready&auto_in_a_valid)
                 begin 
                   if (a_first)
                      counter <=beats1;
                    else 
                      counter <=counter-3'h1;
                   doneAW <=~a_last;
                 end 
              if (nodeOut_r_ready&auto_out_r_valid)
                 begin 
                   r_holds_d <=~auto_out_r_bits_last;
                   r_first <=auto_out_r_bits_last;
                 end 
              count_1 <=count_1+inc-dec;
              count_2 <=count_2+inc_1-dec_1;
              count_3 <=count_3+inc_2-dec_2;
              count_4 <=count_4+inc_3-dec_3;
              count_5 <=count_5+inc_4-dec_4;
              count_6 <=count_6+inc_5-dec_5;
              count_7 <=count_7+inc_6-dec_6;
              count_8 <=count_8+inc_7-dec_7;
              count_9 <=count_9+inc_8-dec_8;
              count_10 <=count_10+inc_9-dec_9;
              count_11 <=count_11+inc_10-dec_10;
              count_12 <=count_12+inc_11-dec_11;
              count_13 <=count_13+inc_12-dec_12;
              count_14 <=count_14+inc_13-dec_13;
              count_15 <=count_15+inc_14-dec_14;
              count_16 <=count_16+inc_15-dec_15;
              count_17 <=count_17+inc_16-dec_16;
              count_18 <=count_18+inc_17-dec_17;
              count_19 <=count_19+inc_18-dec_18;
              count_20 <=count_20+inc_19-dec_19;
              count_21 <=count_21+inc_20-dec_20;
              count_22 <=count_22+inc_21-dec_21;
              count_23 <=count_23+inc_22-dec_22;
              count_24 <=count_24+inc_23-dec_23;
              count_25 <=count_25+inc_24-dec_24;
              count_26 <=count_26+inc_25-dec_25;
              count_27 <=count_27+inc_26-dec_26;
              count_28 <=count_28+inc_27-dec_27;
              count_29 <=count_29+inc_28-dec_28;
              count_30 <=count_30+inc_29-dec_29;
              count_31 <=count_31+inc_30-dec_30;
              count_32 <=count_32+inc_31-dec_31;
              count_33 <=count_33+inc_32-dec_32;
              count_34 <=count_34+inc_33-dec_33;
              count_35 <=count_35+inc_34-dec_34;
              count_36 <=count_36+inc_35-dec_35;
              count_37 <=count_37+inc_36-dec_36;
              count_38 <=count_38+inc_37-dec_37;
              count_39 <=count_39+inc_38-dec_38;
              count_40 <=count_40+inc_39-dec_39;
              count_41 <=count_41+inc_40-dec_40;
              count_42 <=count_42+inc_41-dec_41;
              count_43 <=count_43+inc_42-dec_42;
              count_44 <=count_44+inc_43-dec_43;
              count_45 <=count_45+inc_44-dec_44;
              count_46 <=count_46+inc_45-dec_45;
              count_47 <=count_47+inc_46-dec_46;
              count_48 <=count_48+inc_47-dec_47;
              count_49 <=count_49+inc_48-dec_48;
              count_50 <=count_50+inc_49-dec_49;
              count_51 <=count_51+inc_50-dec_50;
              count_52 <=count_52+inc_51-dec_51;
              count_53 <=count_53+inc_52-dec_52;
              count_54 <=count_54+inc_53-dec_53;
              count_55 <=count_55+inc_54-dec_54;
              count_56 <=count_56+inc_55-dec_55;
              count_57 <=count_57+inc_56-dec_56;
              count_58 <=count_58+inc_57-dec_57;
              count_59 <=count_59+inc_58-dec_58;
              count_60 <=count_60+inc_59-dec_59;
              count_61 <=count_61+inc_60-dec_60;
              count_62 <=count_62+inc_61-dec_61;
              count_63 <=count_63+inc_62-dec_62;
              count_64 <=count_64+inc_63-dec_63;
              count_65 <=count_65+inc_64-dec_64;
              count_66 <=count_66+inc_65-dec_65;
              count_67 <=count_67+inc_66-dec_66;
              count_68 <=count_68+inc_67-dec_67;
              count_69 <=count_69+inc_68-dec_68;
              count_70 <=count_70+inc_69-dec_69;
              count_71 <=count_71+inc_70-dec_70;
              count_72 <=count_72+inc_71-dec_71;
              count_73 <=count_73+inc_72-dec_72;
              count_74 <=count_74+inc_73-dec_73;
              count_75 <=count_75+inc_74-dec_74;
              count_76 <=count_76+inc_75-dec_75;
              count_77 <=count_77+inc_76-dec_76;
              count_78 <=count_78+inc_77-dec_77;
              count_79 <=count_79+inc_78-dec_78;
              count_80 <=count_80+inc_79-dec_79;
              count_81 <=count_81+inc_80-dec_80;
              count_82 <=count_82+inc_81-dec_81;
              count_83 <=count_83+inc_82-dec_82;
              count_84 <=count_84+inc_83-dec_83;
              count_85 <=count_85+inc_84-dec_84;
              count_86 <=count_86+inc_85-dec_85;
              count_87 <=count_87+inc_86-dec_86;
              count_88 <=count_88+inc_87-dec_87;
              count_89 <=count_89+inc_88-dec_88;
              count_90 <=count_90+inc_89-dec_89;
              count_91 <=count_91+inc_90-dec_90;
              count_92 <=count_92+inc_91-dec_91;
              count_93 <=count_93+inc_92-dec_92;
              count_94 <=count_94+inc_93-dec_93;
              count_95 <=count_95+inc_94-dec_94;
              count_96 <=count_96+inc_95-dec_95;
              count_97 <=count_97+inc_96-dec_96;
              count_98 <=count_98+inc_97-dec_97;
              count_99 <=count_99+inc_98-dec_98;
              count_100 <=count_100+inc_99-dec_99;
              count_101 <=count_101+inc_100-dec_100;
              count_102 <=count_102+inc_101-dec_101;
              count_103 <=count_103+inc_102-dec_102;
              count_104 <=count_104+inc_103-dec_103;
              count_105 <=count_105+inc_104-dec_104;
              count_106 <=count_106+inc_105-dec_105;
              count_107 <=count_107+inc_106-dec_106;
              count_108 <=count_108+inc_107-dec_107;
              count_109 <=count_109+inc_108-dec_108;
              count_110 <=count_110+inc_109-dec_109;
              count_111 <=count_111+inc_110-dec_110;
              count_112 <=count_112+inc_111-dec_111;
              count_113 <=count_113+inc_112-dec_112;
              count_114 <=count_114+inc_113-dec_113;
              count_115 <=count_115+inc_114-dec_114;
              count_116 <=count_116+inc_115-dec_115;
              count_117 <=count_117+inc_116-dec_116;
              count_118 <=count_118+inc_117-dec_117;
              count_119 <=count_119+inc_118-dec_118;
              count_120 <=count_120+inc_119-dec_119;
              count_121 <=count_121+inc_120-dec_120;
              count_122 <=count_122+inc_121-dec_121;
              count_123 <=count_123+inc_122-dec_122;
              count_124 <=count_124+inc_123-dec_123;
              count_125 <=count_125+inc_124-dec_124;
              count_126 <=count_126+inc_125-dec_125;
              count_127 <=count_127+inc_126-dec_126;
              count_128 <=count_128+inc_127-dec_127;
            end 
         if (auto_out_b_valid&~nodeOut_b_ready)
            b_delay <=b_delay+3'h1;
          else 
            b_delay <=3'h0;
         if (r_first)
            r_denied_r <=&auto_out_r_bits_resp;
       end
  
  TLMonitor_20 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(nodeIn_d_bits_opcode),.io_in_d_bits_size(nodeIn_d_bits_size),.io_in_d_bits_source(nodeIn_d_bits_source),.io_in_d_bits_denied(nodeIn_d_bits_denied),.io_in_d_bits_corrupt(nodeIn_d_bits_corrupt)); 
  Queue_20 nodeOut_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_w_deq_q_io_enq_ready),.io_enq_valid(~stall&auto_in_a_valid&~(auto_in_a_bits_opcode[2])&_out_w_valid_T_3),.io_enq_bits_data(auto_in_a_bits_data),.io_enq_bits_strb(auto_in_a_bits_mask),.io_enq_bits_last(a_last),.io_deq_ready(auto_out_w_ready),.io_deq_valid(auto_out_w_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last(auto_out_w_bits_last)); 
  Queue_73 queue_arw_deq_q(.clock(clock),.reset(reset),.io_enq_ready(_queue_arw_deq_q_io_enq_ready),.io_enq_valid(out_arw_valid),.io_enq_bits_id(casez_tmp),.io_enq_bits_addr(auto_in_a_bits_address),.io_enq_bits_len(~(_out_arw_bits_len_T_1[10:3])),.io_enq_bits_size(auto_in_a_bits_size>3'h2 ? 3'h3:auto_in_a_bits_size),.io_enq_bits_echo_tl_state_size({1'h0,auto_in_a_bits_size}),.io_enq_bits_echo_tl_state_source(auto_in_a_bits_source),.io_enq_bits_wen(~(auto_in_a_bits_opcode[2])),.io_deq_ready(_queue_arw_deq_q_io_deq_bits_wen ? auto_out_aw_ready:auto_out_ar_ready),.io_deq_valid(_queue_arw_deq_q_io_deq_valid),.io_deq_bits_id(_queue_arw_deq_q_io_deq_bits_id),.io_deq_bits_addr(_queue_arw_deq_q_io_deq_bits_addr),.io_deq_bits_len(_queue_arw_deq_q_io_deq_bits_len),.io_deq_bits_size(_queue_arw_deq_q_io_deq_bits_size),.io_deq_bits_echo_tl_state_size(_queue_arw_deq_q_io_deq_bits_echo_tl_state_size),.io_deq_bits_echo_tl_state_source(_queue_arw_deq_q_io_deq_bits_echo_tl_state_source),.io_deq_bits_wen(_queue_arw_deq_q_io_deq_bits_wen)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=nodeIn_d_bits_opcode; 
  assign auto_in_d_bits_size=nodeIn_d_bits_size; 
  assign auto_in_d_bits_source=nodeIn_d_bits_source; 
  assign auto_in_d_bits_denied=nodeIn_d_bits_denied; 
  assign auto_in_d_bits_data=auto_out_r_bits_data; 
  assign auto_in_d_bits_corrupt=nodeIn_d_bits_corrupt; 
  assign auto_out_aw_valid=_queue_arw_deq_q_io_deq_valid&_queue_arw_deq_q_io_deq_bits_wen; 
  assign auto_out_aw_bits_id=_queue_arw_deq_q_io_deq_bits_id; 
  assign auto_out_aw_bits_addr=_queue_arw_deq_q_io_deq_bits_addr; 
  assign auto_out_aw_bits_len=_queue_arw_deq_q_io_deq_bits_len; 
  assign auto_out_aw_bits_size=_queue_arw_deq_q_io_deq_bits_size; 
  assign auto_out_aw_bits_echo_tl_state_size=_queue_arw_deq_q_io_deq_bits_echo_tl_state_size; 
  assign auto_out_aw_bits_echo_tl_state_source=_queue_arw_deq_q_io_deq_bits_echo_tl_state_source; 
  assign auto_out_b_ready=nodeOut_b_ready; 
  assign auto_out_ar_valid=_queue_arw_deq_q_io_deq_valid&~_queue_arw_deq_q_io_deq_bits_wen; 
  assign auto_out_ar_bits_id=_queue_arw_deq_q_io_deq_bits_id; 
  assign auto_out_ar_bits_addr=_queue_arw_deq_q_io_deq_bits_addr; 
  assign auto_out_ar_bits_len=_queue_arw_deq_q_io_deq_bits_len; 
  assign auto_out_ar_bits_size=_queue_arw_deq_q_io_deq_bits_size; 
  assign auto_out_ar_bits_echo_tl_state_size=_queue_arw_deq_q_io_deq_bits_echo_tl_state_size; 
  assign auto_out_ar_bits_echo_tl_state_source=_queue_arw_deq_q_io_deq_bits_echo_tl_state_source; 
  assign auto_out_r_ready=nodeOut_r_ready; 
endmodule
 
module TLInterconnectCoupler_12 (
  input clock,
  input reset,
  output auto_widget_in_a_ready,
  input auto_widget_in_a_valid,
  input [2:0] auto_widget_in_a_bits_opcode,
  input [2:0] auto_widget_in_a_bits_param,
  input [2:0] auto_widget_in_a_bits_size,
  input [6:0] auto_widget_in_a_bits_source,
  input [31:0] auto_widget_in_a_bits_address,
  input [7:0] auto_widget_in_a_bits_mask,
  input [63:0] auto_widget_in_a_bits_data,
  input auto_widget_in_d_ready,
  output auto_widget_in_d_valid,
  output [2:0] auto_widget_in_d_bits_opcode,
  output [2:0] auto_widget_in_d_bits_size,
  output [6:0] auto_widget_in_d_bits_source,
  output auto_widget_in_d_bits_denied,
  output [63:0] auto_widget_in_d_bits_data,
  output auto_widget_in_d_bits_corrupt,
  input auto_axi4yank_out_aw_ready,
  output auto_axi4yank_out_aw_valid,
  output [3:0] auto_axi4yank_out_aw_bits_id,
  output [31:0] auto_axi4yank_out_aw_bits_addr,
  output [7:0] auto_axi4yank_out_aw_bits_len,
  output [2:0] auto_axi4yank_out_aw_bits_size,
  input auto_axi4yank_out_w_ready,
  output auto_axi4yank_out_w_valid,
  output [63:0] auto_axi4yank_out_w_bits_data,
  output [7:0] auto_axi4yank_out_w_bits_strb,
  output auto_axi4yank_out_w_bits_last,
  output auto_axi4yank_out_b_ready,
  input auto_axi4yank_out_b_valid,
  input [3:0] auto_axi4yank_out_b_bits_id,
  input [1:0] auto_axi4yank_out_b_bits_resp,
  input auto_axi4yank_out_ar_ready,
  output auto_axi4yank_out_ar_valid,
  output [3:0] auto_axi4yank_out_ar_bits_id,
  output [31:0] auto_axi4yank_out_ar_bits_addr,
  output [7:0] auto_axi4yank_out_ar_bits_len,
  output [2:0] auto_axi4yank_out_ar_bits_size,
  output auto_axi4yank_out_r_ready,
  input auto_axi4yank_out_r_valid,
  input [3:0] auto_axi4yank_out_r_bits_id,
  input [63:0] auto_axi4yank_out_r_bits_data,
  input [1:0] auto_axi4yank_out_r_bits_resp,
  input auto_axi4yank_out_r_bits_last,
  output auto_tl_in_a_ready,
  input auto_tl_in_a_valid,
  input [2:0] auto_tl_in_a_bits_opcode,
  input [2:0] auto_tl_in_a_bits_param,
  input [2:0] auto_tl_in_a_bits_size,
  input [6:0] auto_tl_in_a_bits_source,
  input [31:0] auto_tl_in_a_bits_address,
  input [7:0] auto_tl_in_a_bits_mask,
  input [63:0] auto_tl_in_a_bits_data,
  input auto_tl_in_d_ready,
  output auto_tl_in_d_valid,
  output [2:0] auto_tl_in_d_bits_opcode,
  output [2:0] auto_tl_in_d_bits_size,
  output [6:0] auto_tl_in_d_bits_source,
  output auto_tl_in_d_bits_denied,
  output [63:0] auto_tl_in_d_bits_data,
  output auto_tl_in_d_bits_corrupt,
  input auto_tl_out_a_ready,
  output auto_tl_out_a_valid,
  output [2:0] auto_tl_out_a_bits_opcode,
  output [2:0] auto_tl_out_a_bits_param,
  output [2:0] auto_tl_out_a_bits_size,
  output [6:0] auto_tl_out_a_bits_source,
  output [31:0] auto_tl_out_a_bits_address,
  output [7:0] auto_tl_out_a_bits_mask,
  output [63:0] auto_tl_out_a_bits_data,
  output auto_tl_out_d_ready,
  input auto_tl_out_d_valid,
  input [2:0] auto_tl_out_d_bits_opcode,
  input [2:0] auto_tl_out_d_bits_size,
  input [6:0] auto_tl_out_d_bits_source,
  input auto_tl_out_d_bits_denied,
  input [63:0] auto_tl_out_d_bits_data,
  input auto_tl_out_d_bits_corrupt) ; 
   wire _tl2axi4_auto_out_aw_valid ;  
   wire [6:0] _tl2axi4_auto_out_aw_bits_id ;  
   wire [31:0] _tl2axi4_auto_out_aw_bits_addr ;  
   wire [7:0] _tl2axi4_auto_out_aw_bits_len ;  
   wire [2:0] _tl2axi4_auto_out_aw_bits_size ;  
   wire [3:0] _tl2axi4_auto_out_aw_bits_echo_tl_state_size ;  
   wire [6:0] _tl2axi4_auto_out_aw_bits_echo_tl_state_source ;  
   wire _tl2axi4_auto_out_w_valid ;  
   wire [63:0] _tl2axi4_auto_out_w_bits_data ;  
   wire [7:0] _tl2axi4_auto_out_w_bits_strb ;  
   wire _tl2axi4_auto_out_w_bits_last ;  
   wire _tl2axi4_auto_out_b_ready ;  
   wire _tl2axi4_auto_out_ar_valid ;  
   wire [6:0] _tl2axi4_auto_out_ar_bits_id ;  
   wire [31:0] _tl2axi4_auto_out_ar_bits_addr ;  
   wire [7:0] _tl2axi4_auto_out_ar_bits_len ;  
   wire [2:0] _tl2axi4_auto_out_ar_bits_size ;  
   wire [3:0] _tl2axi4_auto_out_ar_bits_echo_tl_state_size ;  
   wire [6:0] _tl2axi4_auto_out_ar_bits_echo_tl_state_source ;  
   wire _tl2axi4_auto_out_r_ready ;  
   wire _axi4index_auto_in_aw_ready ;  
   wire _axi4index_auto_in_w_ready ;  
   wire _axi4index_auto_in_b_valid ;  
   wire [6:0] _axi4index_auto_in_b_bits_id ;  
   wire [1:0] _axi4index_auto_in_b_bits_resp ;  
   wire [3:0] _axi4index_auto_in_b_bits_echo_tl_state_size ;  
   wire [6:0] _axi4index_auto_in_b_bits_echo_tl_state_source ;  
   wire _axi4index_auto_in_ar_ready ;  
   wire _axi4index_auto_in_r_valid ;  
   wire [6:0] _axi4index_auto_in_r_bits_id ;  
   wire [63:0] _axi4index_auto_in_r_bits_data ;  
   wire [1:0] _axi4index_auto_in_r_bits_resp ;  
   wire [3:0] _axi4index_auto_in_r_bits_echo_tl_state_size ;  
   wire [6:0] _axi4index_auto_in_r_bits_echo_tl_state_source ;  
   wire _axi4index_auto_in_r_bits_last ;  
   wire _axi4index_auto_out_aw_valid ;  
   wire [3:0] _axi4index_auto_out_aw_bits_id ;  
   wire [31:0] _axi4index_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4index_auto_out_aw_bits_len ;  
   wire [2:0] _axi4index_auto_out_aw_bits_size ;  
   wire [3:0] _axi4index_auto_out_aw_bits_echo_tl_state_size ;  
   wire [6:0] _axi4index_auto_out_aw_bits_echo_tl_state_source ;  
   wire [2:0] _axi4index_auto_out_aw_bits_echo_extra_id ;  
   wire _axi4index_auto_out_w_valid ;  
   wire [63:0] _axi4index_auto_out_w_bits_data ;  
   wire [7:0] _axi4index_auto_out_w_bits_strb ;  
   wire _axi4index_auto_out_w_bits_last ;  
   wire _axi4index_auto_out_b_ready ;  
   wire _axi4index_auto_out_ar_valid ;  
   wire [3:0] _axi4index_auto_out_ar_bits_id ;  
   wire [31:0] _axi4index_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4index_auto_out_ar_bits_len ;  
   wire [2:0] _axi4index_auto_out_ar_bits_size ;  
   wire [3:0] _axi4index_auto_out_ar_bits_echo_tl_state_size ;  
   wire [6:0] _axi4index_auto_out_ar_bits_echo_tl_state_source ;  
   wire [2:0] _axi4index_auto_out_ar_bits_echo_extra_id ;  
   wire _axi4index_auto_out_r_ready ;  
   wire _axi4yank_auto_in_aw_ready ;  
   wire _axi4yank_auto_in_w_ready ;  
   wire _axi4yank_auto_in_b_valid ;  
   wire [3:0] _axi4yank_auto_in_b_bits_id ;  
   wire [1:0] _axi4yank_auto_in_b_bits_resp ;  
   wire [3:0] _axi4yank_auto_in_b_bits_echo_tl_state_size ;  
   wire [6:0] _axi4yank_auto_in_b_bits_echo_tl_state_source ;  
   wire [2:0] _axi4yank_auto_in_b_bits_echo_extra_id ;  
   wire _axi4yank_auto_in_ar_ready ;  
   wire _axi4yank_auto_in_r_valid ;  
   wire [3:0] _axi4yank_auto_in_r_bits_id ;  
   wire [63:0] _axi4yank_auto_in_r_bits_data ;  
   wire [1:0] _axi4yank_auto_in_r_bits_resp ;  
   wire [3:0] _axi4yank_auto_in_r_bits_echo_tl_state_size ;  
   wire [6:0] _axi4yank_auto_in_r_bits_echo_tl_state_source ;  
   wire [2:0] _axi4yank_auto_in_r_bits_echo_extra_id ;  
   wire _axi4yank_auto_in_r_bits_last ;  
  AXI4UserYanker_2 axi4yank(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4yank_auto_in_aw_ready),.auto_in_aw_valid(_axi4index_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4index_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4index_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4index_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4index_auto_out_aw_bits_size),.auto_in_aw_bits_echo_tl_state_size(_axi4index_auto_out_aw_bits_echo_tl_state_size),.auto_in_aw_bits_echo_tl_state_source(_axi4index_auto_out_aw_bits_echo_tl_state_source),.auto_in_aw_bits_echo_extra_id(_axi4index_auto_out_aw_bits_echo_extra_id),.auto_in_w_ready(_axi4yank_auto_in_w_ready),.auto_in_w_valid(_axi4index_auto_out_w_valid),.auto_in_w_bits_data(_axi4index_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4index_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4index_auto_out_w_bits_last),.auto_in_b_ready(_axi4index_auto_out_b_ready),.auto_in_b_valid(_axi4yank_auto_in_b_valid),.auto_in_b_bits_id(_axi4yank_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4yank_auto_in_b_bits_resp),.auto_in_b_bits_echo_tl_state_size(_axi4yank_auto_in_b_bits_echo_tl_state_size),.auto_in_b_bits_echo_tl_state_source(_axi4yank_auto_in_b_bits_echo_tl_state_source),.auto_in_b_bits_echo_extra_id(_axi4yank_auto_in_b_bits_echo_extra_id),.auto_in_ar_ready(_axi4yank_auto_in_ar_ready),.auto_in_ar_valid(_axi4index_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4index_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4index_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4index_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4index_auto_out_ar_bits_size),.auto_in_ar_bits_echo_tl_state_size(_axi4index_auto_out_ar_bits_echo_tl_state_size),.auto_in_ar_bits_echo_tl_state_source(_axi4index_auto_out_ar_bits_echo_tl_state_source),.auto_in_ar_bits_echo_extra_id(_axi4index_auto_out_ar_bits_echo_extra_id),.auto_in_r_ready(_axi4index_auto_out_r_ready),.auto_in_r_valid(_axi4yank_auto_in_r_valid),.auto_in_r_bits_id(_axi4yank_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4yank_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4yank_auto_in_r_bits_resp),.auto_in_r_bits_echo_tl_state_size(_axi4yank_auto_in_r_bits_echo_tl_state_size),.auto_in_r_bits_echo_tl_state_source(_axi4yank_auto_in_r_bits_echo_tl_state_source),.auto_in_r_bits_echo_extra_id(_axi4yank_auto_in_r_bits_echo_extra_id),.auto_in_r_bits_last(_axi4yank_auto_in_r_bits_last),.auto_out_aw_ready(auto_axi4yank_out_aw_ready),.auto_out_aw_valid(auto_axi4yank_out_aw_valid),.auto_out_aw_bits_id(auto_axi4yank_out_aw_bits_id),.auto_out_aw_bits_addr(auto_axi4yank_out_aw_bits_addr),.auto_out_aw_bits_len(auto_axi4yank_out_aw_bits_len),.auto_out_aw_bits_size(auto_axi4yank_out_aw_bits_size),.auto_out_w_ready(auto_axi4yank_out_w_ready),.auto_out_w_valid(auto_axi4yank_out_w_valid),.auto_out_w_bits_data(auto_axi4yank_out_w_bits_data),.auto_out_w_bits_strb(auto_axi4yank_out_w_bits_strb),.auto_out_w_bits_last(auto_axi4yank_out_w_bits_last),.auto_out_b_ready(auto_axi4yank_out_b_ready),.auto_out_b_valid(auto_axi4yank_out_b_valid),.auto_out_b_bits_id(auto_axi4yank_out_b_bits_id),.auto_out_b_bits_resp(auto_axi4yank_out_b_bits_resp),.auto_out_ar_ready(auto_axi4yank_out_ar_ready),.auto_out_ar_valid(auto_axi4yank_out_ar_valid),.auto_out_ar_bits_id(auto_axi4yank_out_ar_bits_id),.auto_out_ar_bits_addr(auto_axi4yank_out_ar_bits_addr),.auto_out_ar_bits_len(auto_axi4yank_out_ar_bits_len),.auto_out_ar_bits_size(auto_axi4yank_out_ar_bits_size),.auto_out_r_ready(auto_axi4yank_out_r_ready),.auto_out_r_valid(auto_axi4yank_out_r_valid),.auto_out_r_bits_id(auto_axi4yank_out_r_bits_id),.auto_out_r_bits_data(auto_axi4yank_out_r_bits_data),.auto_out_r_bits_resp(auto_axi4yank_out_r_bits_resp),.auto_out_r_bits_last(auto_axi4yank_out_r_bits_last)); 
  AXI4IdIndexer_2 axi4index(.auto_in_aw_ready(_axi4index_auto_in_aw_ready),.auto_in_aw_valid(_tl2axi4_auto_out_aw_valid),.auto_in_aw_bits_id(_tl2axi4_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_tl2axi4_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_tl2axi4_auto_out_aw_bits_len),.auto_in_aw_bits_size(_tl2axi4_auto_out_aw_bits_size),.auto_in_aw_bits_echo_tl_state_size(_tl2axi4_auto_out_aw_bits_echo_tl_state_size),.auto_in_aw_bits_echo_tl_state_source(_tl2axi4_auto_out_aw_bits_echo_tl_state_source),.auto_in_w_ready(_axi4index_auto_in_w_ready),.auto_in_w_valid(_tl2axi4_auto_out_w_valid),.auto_in_w_bits_data(_tl2axi4_auto_out_w_bits_data),.auto_in_w_bits_strb(_tl2axi4_auto_out_w_bits_strb),.auto_in_w_bits_last(_tl2axi4_auto_out_w_bits_last),.auto_in_b_ready(_tl2axi4_auto_out_b_ready),.auto_in_b_valid(_axi4index_auto_in_b_valid),.auto_in_b_bits_id(_axi4index_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4index_auto_in_b_bits_resp),.auto_in_b_bits_echo_tl_state_size(_axi4index_auto_in_b_bits_echo_tl_state_size),.auto_in_b_bits_echo_tl_state_source(_axi4index_auto_in_b_bits_echo_tl_state_source),.auto_in_ar_ready(_axi4index_auto_in_ar_ready),.auto_in_ar_valid(_tl2axi4_auto_out_ar_valid),.auto_in_ar_bits_id(_tl2axi4_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_tl2axi4_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_tl2axi4_auto_out_ar_bits_len),.auto_in_ar_bits_size(_tl2axi4_auto_out_ar_bits_size),.auto_in_ar_bits_echo_tl_state_size(_tl2axi4_auto_out_ar_bits_echo_tl_state_size),.auto_in_ar_bits_echo_tl_state_source(_tl2axi4_auto_out_ar_bits_echo_tl_state_source),.auto_in_r_ready(_tl2axi4_auto_out_r_ready),.auto_in_r_valid(_axi4index_auto_in_r_valid),.auto_in_r_bits_id(_axi4index_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4index_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4index_auto_in_r_bits_resp),.auto_in_r_bits_echo_tl_state_size(_axi4index_auto_in_r_bits_echo_tl_state_size),.auto_in_r_bits_echo_tl_state_source(_axi4index_auto_in_r_bits_echo_tl_state_source),.auto_in_r_bits_last(_axi4index_auto_in_r_bits_last),.auto_out_aw_ready(_axi4yank_auto_in_aw_ready),.auto_out_aw_valid(_axi4index_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4index_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4index_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4index_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4index_auto_out_aw_bits_size),.auto_out_aw_bits_echo_tl_state_size(_axi4index_auto_out_aw_bits_echo_tl_state_size),.auto_out_aw_bits_echo_tl_state_source(_axi4index_auto_out_aw_bits_echo_tl_state_source),.auto_out_aw_bits_echo_extra_id(_axi4index_auto_out_aw_bits_echo_extra_id),.auto_out_w_ready(_axi4yank_auto_in_w_ready),.auto_out_w_valid(_axi4index_auto_out_w_valid),.auto_out_w_bits_data(_axi4index_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4index_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4index_auto_out_w_bits_last),.auto_out_b_ready(_axi4index_auto_out_b_ready),.auto_out_b_valid(_axi4yank_auto_in_b_valid),.auto_out_b_bits_id(_axi4yank_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4yank_auto_in_b_bits_resp),.auto_out_b_bits_echo_tl_state_size(_axi4yank_auto_in_b_bits_echo_tl_state_size),.auto_out_b_bits_echo_tl_state_source(_axi4yank_auto_in_b_bits_echo_tl_state_source),.auto_out_b_bits_echo_extra_id(_axi4yank_auto_in_b_bits_echo_extra_id),.auto_out_ar_ready(_axi4yank_auto_in_ar_ready),.auto_out_ar_valid(_axi4index_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4index_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4index_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4index_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4index_auto_out_ar_bits_size),.auto_out_ar_bits_echo_tl_state_size(_axi4index_auto_out_ar_bits_echo_tl_state_size),.auto_out_ar_bits_echo_tl_state_source(_axi4index_auto_out_ar_bits_echo_tl_state_source),.auto_out_ar_bits_echo_extra_id(_axi4index_auto_out_ar_bits_echo_extra_id),.auto_out_r_ready(_axi4index_auto_out_r_ready),.auto_out_r_valid(_axi4yank_auto_in_r_valid),.auto_out_r_bits_id(_axi4yank_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4yank_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4yank_auto_in_r_bits_resp),.auto_out_r_bits_echo_tl_state_size(_axi4yank_auto_in_r_bits_echo_tl_state_size),.auto_out_r_bits_echo_tl_state_source(_axi4yank_auto_in_r_bits_echo_tl_state_source),.auto_out_r_bits_echo_extra_id(_axi4yank_auto_in_r_bits_echo_extra_id),.auto_out_r_bits_last(_axi4yank_auto_in_r_bits_last)); 
  TLToAXI4_1 tl2axi4(.clock(clock),.reset(reset),.auto_in_a_ready(auto_widget_in_a_ready),.auto_in_a_valid(auto_widget_in_a_valid),.auto_in_a_bits_opcode(auto_widget_in_a_bits_opcode),.auto_in_a_bits_param(auto_widget_in_a_bits_param),.auto_in_a_bits_size(auto_widget_in_a_bits_size),.auto_in_a_bits_source(auto_widget_in_a_bits_source),.auto_in_a_bits_address(auto_widget_in_a_bits_address),.auto_in_a_bits_mask(auto_widget_in_a_bits_mask),.auto_in_a_bits_data(auto_widget_in_a_bits_data),.auto_in_d_ready(auto_widget_in_d_ready),.auto_in_d_valid(auto_widget_in_d_valid),.auto_in_d_bits_opcode(auto_widget_in_d_bits_opcode),.auto_in_d_bits_size(auto_widget_in_d_bits_size),.auto_in_d_bits_source(auto_widget_in_d_bits_source),.auto_in_d_bits_denied(auto_widget_in_d_bits_denied),.auto_in_d_bits_data(auto_widget_in_d_bits_data),.auto_in_d_bits_corrupt(auto_widget_in_d_bits_corrupt),.auto_out_aw_ready(_axi4index_auto_in_aw_ready),.auto_out_aw_valid(_tl2axi4_auto_out_aw_valid),.auto_out_aw_bits_id(_tl2axi4_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_tl2axi4_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_tl2axi4_auto_out_aw_bits_len),.auto_out_aw_bits_size(_tl2axi4_auto_out_aw_bits_size),.auto_out_aw_bits_echo_tl_state_size(_tl2axi4_auto_out_aw_bits_echo_tl_state_size),.auto_out_aw_bits_echo_tl_state_source(_tl2axi4_auto_out_aw_bits_echo_tl_state_source),.auto_out_w_ready(_axi4index_auto_in_w_ready),.auto_out_w_valid(_tl2axi4_auto_out_w_valid),.auto_out_w_bits_data(_tl2axi4_auto_out_w_bits_data),.auto_out_w_bits_strb(_tl2axi4_auto_out_w_bits_strb),.auto_out_w_bits_last(_tl2axi4_auto_out_w_bits_last),.auto_out_b_ready(_tl2axi4_auto_out_b_ready),.auto_out_b_valid(_axi4index_auto_in_b_valid),.auto_out_b_bits_id(_axi4index_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4index_auto_in_b_bits_resp),.auto_out_b_bits_echo_tl_state_size(_axi4index_auto_in_b_bits_echo_tl_state_size),.auto_out_b_bits_echo_tl_state_source(_axi4index_auto_in_b_bits_echo_tl_state_source),.auto_out_ar_ready(_axi4index_auto_in_ar_ready),.auto_out_ar_valid(_tl2axi4_auto_out_ar_valid),.auto_out_ar_bits_id(_tl2axi4_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_tl2axi4_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_tl2axi4_auto_out_ar_bits_len),.auto_out_ar_bits_size(_tl2axi4_auto_out_ar_bits_size),.auto_out_ar_bits_echo_tl_state_size(_tl2axi4_auto_out_ar_bits_echo_tl_state_size),.auto_out_ar_bits_echo_tl_state_source(_tl2axi4_auto_out_ar_bits_echo_tl_state_source),.auto_out_r_ready(_tl2axi4_auto_out_r_ready),.auto_out_r_valid(_axi4index_auto_in_r_valid),.auto_out_r_bits_id(_axi4index_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4index_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4index_auto_in_r_bits_resp),.auto_out_r_bits_echo_tl_state_size(_axi4index_auto_in_r_bits_echo_tl_state_size),.auto_out_r_bits_echo_tl_state_source(_axi4index_auto_in_r_bits_echo_tl_state_source),.auto_out_r_bits_last(_axi4index_auto_in_r_bits_last)); 
  assign auto_tl_in_a_ready=auto_tl_out_a_ready; 
  assign auto_tl_in_d_valid=auto_tl_out_d_valid; 
  assign auto_tl_in_d_bits_opcode=auto_tl_out_d_bits_opcode; 
  assign auto_tl_in_d_bits_size=auto_tl_out_d_bits_size; 
  assign auto_tl_in_d_bits_source=auto_tl_out_d_bits_source; 
  assign auto_tl_in_d_bits_denied=auto_tl_out_d_bits_denied; 
  assign auto_tl_in_d_bits_data=auto_tl_out_d_bits_data; 
  assign auto_tl_in_d_bits_corrupt=auto_tl_out_d_bits_corrupt; 
  assign auto_tl_out_a_valid=auto_tl_in_a_valid; 
  assign auto_tl_out_a_bits_opcode=auto_tl_in_a_bits_opcode; 
  assign auto_tl_out_a_bits_param=auto_tl_in_a_bits_param; 
  assign auto_tl_out_a_bits_size=auto_tl_in_a_bits_size; 
  assign auto_tl_out_a_bits_source=auto_tl_in_a_bits_source; 
  assign auto_tl_out_a_bits_address=auto_tl_in_a_bits_address; 
  assign auto_tl_out_a_bits_mask=auto_tl_in_a_bits_mask; 
  assign auto_tl_out_a_bits_data=auto_tl_in_a_bits_data; 
  assign auto_tl_out_d_ready=auto_tl_in_d_ready; 
endmodule
 
module MemoryBus (
  input auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready,
  output auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid,
  output [3:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id,
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr,
  output [7:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len,
  output [2:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size,
  input auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready,
  output auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid,
  output [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data,
  output [7:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb,
  output auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last,
  output auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready,
  input auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid,
  input [3:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id,
  input [1:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp,
  input auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready,
  output auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid,
  output [3:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id,
  output [31:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr,
  output [7:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len,
  output [2:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size,
  output auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready,
  input auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid,
  input [3:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id,
  input [63:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data,
  input [1:0] auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp,
  input auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last,
  input auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock,
  input auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset,
  output auto_bus_xing_in_a_ready,
  input auto_bus_xing_in_a_valid,
  input [2:0] auto_bus_xing_in_a_bits_opcode,
  input [2:0] auto_bus_xing_in_a_bits_param,
  input [2:0] auto_bus_xing_in_a_bits_size,
  input [6:0] auto_bus_xing_in_a_bits_source,
  input [31:0] auto_bus_xing_in_a_bits_address,
  input [7:0] auto_bus_xing_in_a_bits_mask,
  input [63:0] auto_bus_xing_in_a_bits_data,
  input auto_bus_xing_in_d_ready,
  output auto_bus_xing_in_d_valid,
  output [2:0] auto_bus_xing_in_d_bits_opcode,
  output [2:0] auto_bus_xing_in_d_bits_size,
  output [6:0] auto_bus_xing_in_d_bits_source,
  output auto_bus_xing_in_d_bits_denied,
  output [63:0] auto_bus_xing_in_d_bits_data,
  output auto_bus_xing_in_d_bits_corrupt) ; 
   wire _coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_ready ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_valid ;  
   wire [2:0] _coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_opcode ;  
   wire [2:0] _coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_size ;  
   wire [6:0] _coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_source ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_denied ;  
   wire [63:0] _coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_data ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_corrupt ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid ;  
   wire [2:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode ;  
   wire [2:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size ;  
   wire [6:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied ;  
   wire [63:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_valid ;  
   wire [2:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_opcode ;  
   wire [2:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_param ;  
   wire [2:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_size ;  
   wire [6:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_source ;  
   wire [31:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_address ;  
   wire [7:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_mask ;  
   wire [63:0] _coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_data ;  
   wire _coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_ready ;  
   wire _picker_auto_in_a_ready ;  
   wire _picker_auto_in_d_valid ;  
   wire [2:0] _picker_auto_in_d_bits_opcode ;  
   wire [2:0] _picker_auto_in_d_bits_size ;  
   wire [6:0] _picker_auto_in_d_bits_source ;  
   wire _picker_auto_in_d_bits_denied ;  
   wire [63:0] _picker_auto_in_d_bits_data ;  
   wire _picker_auto_in_d_bits_corrupt ;  
   wire _picker_auto_out_a_valid ;  
   wire [2:0] _picker_auto_out_a_bits_opcode ;  
   wire [2:0] _picker_auto_out_a_bits_param ;  
   wire [2:0] _picker_auto_out_a_bits_size ;  
   wire [6:0] _picker_auto_out_a_bits_source ;  
   wire [31:0] _picker_auto_out_a_bits_address ;  
   wire [7:0] _picker_auto_out_a_bits_mask ;  
   wire [63:0] _picker_auto_out_a_bits_data ;  
   wire _picker_auto_out_d_ready ;  
   wire _fixer_auto_out_a_valid ;  
   wire [2:0] _fixer_auto_out_a_bits_opcode ;  
   wire [2:0] _fixer_auto_out_a_bits_param ;  
   wire [2:0] _fixer_auto_out_a_bits_size ;  
   wire [6:0] _fixer_auto_out_a_bits_source ;  
   wire [31:0] _fixer_auto_out_a_bits_address ;  
   wire [7:0] _fixer_auto_out_a_bits_mask ;  
   wire [63:0] _fixer_auto_out_a_bits_data ;  
   wire _fixer_auto_out_d_ready ;  
  TLFIFOFixer_4 fixer(.clock(auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),.reset(auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),.auto_in_a_ready(auto_bus_xing_in_a_ready),.auto_in_a_valid(auto_bus_xing_in_a_valid),.auto_in_a_bits_opcode(auto_bus_xing_in_a_bits_opcode),.auto_in_a_bits_param(auto_bus_xing_in_a_bits_param),.auto_in_a_bits_size(auto_bus_xing_in_a_bits_size),.auto_in_a_bits_source(auto_bus_xing_in_a_bits_source),.auto_in_a_bits_address(auto_bus_xing_in_a_bits_address),.auto_in_a_bits_mask(auto_bus_xing_in_a_bits_mask),.auto_in_a_bits_data(auto_bus_xing_in_a_bits_data),.auto_in_d_ready(auto_bus_xing_in_d_ready),.auto_in_d_valid(auto_bus_xing_in_d_valid),.auto_in_d_bits_opcode(auto_bus_xing_in_d_bits_opcode),.auto_in_d_bits_size(auto_bus_xing_in_d_bits_size),.auto_in_d_bits_source(auto_bus_xing_in_d_bits_source),.auto_in_d_bits_denied(auto_bus_xing_in_d_bits_denied),.auto_in_d_bits_data(auto_bus_xing_in_d_bits_data),.auto_in_d_bits_corrupt(auto_bus_xing_in_d_bits_corrupt),.auto_out_a_ready(_picker_auto_in_a_ready),.auto_out_a_valid(_fixer_auto_out_a_valid),.auto_out_a_bits_opcode(_fixer_auto_out_a_bits_opcode),.auto_out_a_bits_param(_fixer_auto_out_a_bits_param),.auto_out_a_bits_size(_fixer_auto_out_a_bits_size),.auto_out_a_bits_source(_fixer_auto_out_a_bits_source),.auto_out_a_bits_address(_fixer_auto_out_a_bits_address),.auto_out_a_bits_mask(_fixer_auto_out_a_bits_mask),.auto_out_a_bits_data(_fixer_auto_out_a_bits_data),.auto_out_d_ready(_fixer_auto_out_d_ready),.auto_out_d_valid(_picker_auto_in_d_valid),.auto_out_d_bits_opcode(_picker_auto_in_d_bits_opcode),.auto_out_d_bits_size(_picker_auto_in_d_bits_size),.auto_out_d_bits_source(_picker_auto_in_d_bits_source),.auto_out_d_bits_denied(_picker_auto_in_d_bits_denied),.auto_out_d_bits_data(_picker_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_picker_auto_in_d_bits_corrupt)); 
  ProbePicker picker(.clock(auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),.reset(auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),.auto_in_a_ready(_picker_auto_in_a_ready),.auto_in_a_valid(_fixer_auto_out_a_valid),.auto_in_a_bits_opcode(_fixer_auto_out_a_bits_opcode),.auto_in_a_bits_param(_fixer_auto_out_a_bits_param),.auto_in_a_bits_size(_fixer_auto_out_a_bits_size),.auto_in_a_bits_source(_fixer_auto_out_a_bits_source),.auto_in_a_bits_address(_fixer_auto_out_a_bits_address),.auto_in_a_bits_mask(_fixer_auto_out_a_bits_mask),.auto_in_a_bits_data(_fixer_auto_out_a_bits_data),.auto_in_d_ready(_fixer_auto_out_d_ready),.auto_in_d_valid(_picker_auto_in_d_valid),.auto_in_d_bits_opcode(_picker_auto_in_d_bits_opcode),.auto_in_d_bits_size(_picker_auto_in_d_bits_size),.auto_in_d_bits_source(_picker_auto_in_d_bits_source),.auto_in_d_bits_denied(_picker_auto_in_d_bits_denied),.auto_in_d_bits_data(_picker_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_picker_auto_in_d_bits_corrupt),.auto_out_a_ready(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready),.auto_out_a_valid(_picker_auto_out_a_valid),.auto_out_a_bits_opcode(_picker_auto_out_a_bits_opcode),.auto_out_a_bits_param(_picker_auto_out_a_bits_param),.auto_out_a_bits_size(_picker_auto_out_a_bits_size),.auto_out_a_bits_source(_picker_auto_out_a_bits_source),.auto_out_a_bits_address(_picker_auto_out_a_bits_address),.auto_out_a_bits_mask(_picker_auto_out_a_bits_mask),.auto_out_a_bits_data(_picker_auto_out_a_bits_data),.auto_out_d_ready(_picker_auto_out_d_ready),.auto_out_d_valid(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid),.auto_out_d_bits_opcode(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode),.auto_out_d_bits_size(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size),.auto_out_d_bits_source(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source),.auto_out_d_bits_denied(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied),.auto_out_d_bits_data(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data),.auto_out_d_bits_corrupt(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt)); 
  TLInterconnectCoupler_12 coupler_to_memory_controller_port_named_axi4(.clock(auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock),.reset(auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset),.auto_widget_in_a_ready(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_ready),.auto_widget_in_a_valid(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_valid),.auto_widget_in_a_bits_opcode(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_opcode),.auto_widget_in_a_bits_param(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_param),.auto_widget_in_a_bits_size(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_size),.auto_widget_in_a_bits_source(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_source),.auto_widget_in_a_bits_address(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_address),.auto_widget_in_a_bits_mask(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_mask),.auto_widget_in_a_bits_data(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_data),.auto_widget_in_d_ready(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_ready),.auto_widget_in_d_valid(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_valid),.auto_widget_in_d_bits_opcode(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_opcode),.auto_widget_in_d_bits_size(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_size),.auto_widget_in_d_bits_source(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_source),.auto_widget_in_d_bits_denied(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_denied),.auto_widget_in_d_bits_data(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_data),.auto_widget_in_d_bits_corrupt(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_corrupt),.auto_axi4yank_out_aw_ready(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready),.auto_axi4yank_out_aw_valid(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid),.auto_axi4yank_out_aw_bits_id(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id),.auto_axi4yank_out_aw_bits_addr(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr),.auto_axi4yank_out_aw_bits_len(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len),.auto_axi4yank_out_aw_bits_size(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size),.auto_axi4yank_out_w_ready(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready),.auto_axi4yank_out_w_valid(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid),.auto_axi4yank_out_w_bits_data(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data),.auto_axi4yank_out_w_bits_strb(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb),.auto_axi4yank_out_w_bits_last(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last),.auto_axi4yank_out_b_ready(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready),.auto_axi4yank_out_b_valid(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid),.auto_axi4yank_out_b_bits_id(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id),.auto_axi4yank_out_b_bits_resp(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp),.auto_axi4yank_out_ar_ready(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready),.auto_axi4yank_out_ar_valid(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid),.auto_axi4yank_out_ar_bits_id(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id),.auto_axi4yank_out_ar_bits_addr(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr),.auto_axi4yank_out_ar_bits_len(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len),.auto_axi4yank_out_ar_bits_size(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size),.auto_axi4yank_out_r_ready(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready),.auto_axi4yank_out_r_valid(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid),.auto_axi4yank_out_r_bits_id(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id),.auto_axi4yank_out_r_bits_data(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data),.auto_axi4yank_out_r_bits_resp(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp),.auto_axi4yank_out_r_bits_last(auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last),.auto_tl_in_a_ready(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_a_ready),.auto_tl_in_a_valid(_picker_auto_out_a_valid),.auto_tl_in_a_bits_opcode(_picker_auto_out_a_bits_opcode),.auto_tl_in_a_bits_param(_picker_auto_out_a_bits_param),.auto_tl_in_a_bits_size(_picker_auto_out_a_bits_size),.auto_tl_in_a_bits_source(_picker_auto_out_a_bits_source),.auto_tl_in_a_bits_address(_picker_auto_out_a_bits_address),.auto_tl_in_a_bits_mask(_picker_auto_out_a_bits_mask),.auto_tl_in_a_bits_data(_picker_auto_out_a_bits_data),.auto_tl_in_d_ready(_picker_auto_out_d_ready),.auto_tl_in_d_valid(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_valid),.auto_tl_in_d_bits_opcode(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_opcode),.auto_tl_in_d_bits_size(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_size),.auto_tl_in_d_bits_source(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_source),.auto_tl_in_d_bits_denied(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_denied),.auto_tl_in_d_bits_data(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_data),.auto_tl_in_d_bits_corrupt(_coupler_to_memory_controller_port_named_axi4_auto_tl_in_d_bits_corrupt),.auto_tl_out_a_ready(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_a_ready),.auto_tl_out_a_valid(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_valid),.auto_tl_out_a_bits_opcode(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_opcode),.auto_tl_out_a_bits_param(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_param),.auto_tl_out_a_bits_size(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_size),.auto_tl_out_a_bits_source(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_source),.auto_tl_out_a_bits_address(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_address),.auto_tl_out_a_bits_mask(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_mask),.auto_tl_out_a_bits_data(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_a_bits_data),.auto_tl_out_d_ready(_coupler_to_memory_controller_port_named_axi4_auto_tl_out_d_ready),.auto_tl_out_d_valid(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_valid),.auto_tl_out_d_bits_opcode(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_opcode),.auto_tl_out_d_bits_size(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_size),.auto_tl_out_d_bits_source(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_source),.auto_tl_out_d_bits_denied(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_denied),.auto_tl_out_d_bits_data(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_data),.auto_tl_out_d_bits_corrupt(_coupler_to_memory_controller_port_named_axi4_auto_widget_in_d_bits_corrupt)); 
endmodule
 
module TLMonitor_21 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_b_ready,
  input io_in_b_valid,
  input [1:0] io_in_b_bits_param,
  input [31:0] io_in_b_bits_address,
  input io_in_c_ready,
  input io_in_c_valid,
  input [2:0] io_in_c_bits_opcode,
  input [2:0] io_in_c_bits_param,
  input [2:0] io_in_c_bits_size,
  input [4:0] io_in_c_bits_source,
  input [31:0] io_in_c_bits_address,
  input io_in_c_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [2:0] io_in_d_bits_size,
  input [4:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt,
  input io_in_e_valid,
  input [1:0] io_in_e_bits_sink) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire [12:0] _GEN_0={10'h0,io_in_c_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [31:0] address ;  
   wire _d_first_T_3=io_in_d_ready&io_in_d_valid ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [2:0] size_1 ;  
   reg [4:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [2:0] b_first_counter ;  
   reg [1:0] param_2 ;  
   reg [31:0] address_1 ;  
   wire _c_first_T_1=io_in_c_ready&io_in_c_valid ;  
   reg [2:0] c_first_counter ;  
   reg [2:0] opcode_3 ;  
   reg [2:0] param_3 ;  
   reg [2:0] size_3 ;  
   reg [4:0] source_3 ;  
   reg [31:0] address_2 ;  
   reg [18:0] inflight ;  
   reg [75:0] inflight_opcodes ;  
   reg [75:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [75:0] _GEN_1={69'h0,io_in_d_bits_source,2'h0} ;  
   wire [75:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_1 ;  
   wire [31:0] _GEN_2={27'h0,io_in_a_bits_source} ;  
   wire _GEN_3=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [31:0] _GEN_4={27'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [18:0] inflight_1 ;  
   reg [75:0] inflight_sizes_1 ;  
   reg [2:0] c_first_counter_1 ;  
   wire c_first_1=c_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   wire _GEN_5=io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1] ;  
   wire [31:0] _GEN_6={27'h0,io_in_c_bits_source} ;  
   wire _GEN_7=_c_first_T_1&c_first_1&_GEN_5 ;  
   reg [31:0] watchdog_1 ;  
   reg [3:0] inflight_2 ;  
   reg [2:0] d_first_counter_3 ;  
   wire d_first_3=d_first_counter_3==3'h0 ;  
   wire _GEN_8=_d_first_T_3&d_first_3&io_in_d_bits_opcode[2]&~(io_in_d_bits_opcode[1]) ;  
   wire [3:0] _GEN_9={2'h0,io_in_d_bits_sink} ;  
   wire [3:0] d_set=_GEN_8 ? 4'h1<<_GEN_9:4'h0 ;  
   wire [3:0] _GEN_10={2'h0,io_in_e_bits_sink} ;  
   wire _source_ok_T_12=io_in_a_bits_source==5'h10 ;  
   wire _source_ok_T_13=io_in_a_bits_source==5'h11 ;  
   wire _source_ok_T_14=io_in_a_bits_source==5'h12 ;  
   wire source_ok=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_11=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_12=~(|(io_in_a_bits_source[4:3]))|io_in_a_bits_source[4:3]==2'h1|_source_ok_T_12|_source_ok_T_13|_source_ok_T_14 ;  
   wire _GEN_13=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_14=io_in_a_bits_size!=3'h7&_GEN_13 ;  
   wire _GEN_15=_GEN_12&_GEN_14 ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_17=_source_ok_T_12&io_in_a_bits_size==3'h6&_GEN_13 ;  
   wire _GEN_18=io_in_a_bits_param>3'h2 ;  
   wire _GEN_19=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_20=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_21=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_22=io_in_a_bits_mask!=mask ;  
   wire _GEN_23=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_24=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_25=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_26=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_27=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source[4:3]==2'h0|io_in_d_bits_source[4:3]==2'h1|io_in_d_bits_source==5'h10|io_in_d_bits_source==5'h11|io_in_d_bits_source==5'h12 ;  
   wire _GEN_28=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_29=io_in_d_bits_size<3'h3 ;  
   wire _GEN_30=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_31=io_in_d_bits_param==2'h2 ;  
   wire _GEN_32=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_33=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_34=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_35=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_36=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_37=io_in_b_valid&~reset ;  
   wire _source_ok_T_48=io_in_c_bits_source==5'h10 ;  
   wire _source_ok_T_49=io_in_c_bits_source==5'h11 ;  
   wire _source_ok_T_50=io_in_c_bits_source==5'h12 ;  
   wire source_ok_2=~(|(io_in_c_bits_source[4:3]))|io_in_c_bits_source[4:3]==2'h1|_source_ok_T_48|_source_ok_T_49|_source_ok_T_50 ;  
   wire [12:0] _is_aligned_mask_T_7=13'h3F<<_GEN_0 ;  
   wire [5:0] _GEN_38=io_in_c_bits_address[5:0]&~(_is_aligned_mask_T_7[5:0]) ;  
   wire _GEN_39=io_in_c_bits_address[31:28]!=4'h8 ;  
   wire _GEN_40=io_in_c_valid&io_in_c_bits_opcode==3'h4&~reset ;  
   wire _GEN_41=io_in_c_bits_size<3'h3 ;  
   wire _GEN_42=io_in_c_valid&io_in_c_bits_opcode==3'h5&~reset ;  
   wire _GEN_43=(~(|(io_in_c_bits_source[4:3]))|io_in_c_bits_source[4:3]==2'h1|_source_ok_T_48|_source_ok_T_49|_source_ok_T_50)&io_in_c_bits_size!=3'h7&~_GEN_39 ;  
   wire _GEN_44=io_in_c_valid&io_in_c_bits_opcode==3'h6&~reset ;  
   wire _GEN_45=_source_ok_T_48&io_in_c_bits_size==3'h6&~_GEN_39 ;  
   wire _GEN_46=io_in_c_valid&(&io_in_c_bits_opcode)&~reset ;  
   wire _GEN_47=io_in_c_valid&io_in_c_bits_opcode==3'h0&~reset ;  
   wire _GEN_48=io_in_c_valid&io_in_c_bits_opcode==3'h1&~reset ;  
   wire _GEN_49=io_in_c_valid&io_in_c_bits_opcode==3'h2&~reset ;  
   wire _GEN_50=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_51=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_52=io_in_b_valid&(|b_first_counter)&~reset ;  
   wire _GEN_53=io_in_c_valid&(|c_first_counter)&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [31:0] _a_set_wo_ready_T=32'h1<<_GEN_2 ;  
   wire [18:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_54=io_in_d_valid&d_first_1 ;  
   wire _GEN_55=_GEN_54&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_56={14'h0,io_in_d_bits_source} ;  
   wire _GEN_57=_GEN_55&same_cycle_resp&~reset ;  
   wire _GEN_58=_GEN_55&~same_cycle_resp&~reset ;  
   wire _same_cycle_resp_T_3=io_in_c_valid&c_first_1 ;  
   wire [31:0] _c_set_wo_ready_T=32'h1<<_GEN_6 ;  
   wire [18:0] c_set_wo_ready=_same_cycle_resp_T_3&_GEN_5 ? _c_set_wo_ready_T[18:0]:19'h0 ;  
   wire _GEN_59=io_in_d_valid&d_first_2 ;  
   wire _GEN_60=_GEN_59&d_release_ack ;  
   wire same_cycle_resp_1=_same_cycle_resp_T_3&io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1]&io_in_c_bits_source==io_in_d_bits_source ;  
   wire [18:0] _GEN_61=inflight>>io_in_a_bits_source ;  
   wire [18:0] _GEN_62=inflight>>_GEN_56 ;  
   wire [75:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_1 ;  
   wire [31:0] _d_clr_wo_ready_T=32'h1<<_GEN_4 ;  
   wire [18:0] _GEN_63=inflight_1>>io_in_c_bits_source ;  
   wire [18:0] _GEN_64=inflight_1>>_GEN_56 ;  
   wire [75:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_1 ;  
   wire [31:0] _d_clr_wo_ready_T_1=32'h1<<_GEN_4 ;  
   wire [3:0] _GEN_65=inflight_2>>_GEN_9 ;  
   wire [3:0] _GEN_66=(d_set|inflight_2)>>_GEN_10 ;  
  always @( posedge clock)
       begin 
         if (_GEN_16&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&_GEN_29)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~_GEN_33)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~_GEN_33)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_b_bits_address[31:28]!=4'h8)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|(io_in_b_bits_address[5:0])))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(&io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&(|_GEN_38))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&(|_GEN_38))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~_GEN_45)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&(|_GEN_38))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid report param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&~_GEN_45)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&(|_GEN_38))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&(|_GEN_38))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_48&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_48&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_48&(|_GEN_38))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_48&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_49&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_49&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_49&(|_GEN_38))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_49&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_49&io_in_c_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_50&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_50&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_50&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_50&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_50&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_51&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_51&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_51&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_51&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_51&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_51&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_52&io_in_b_bits_param!=param_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel param changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_52&io_in_b_bits_address!=address_1)
            begin 
              if (1)$display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&io_in_c_bits_opcode!=opcode_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&io_in_c_bits_param!=param_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel param changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&io_in_c_bits_size!=size_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel size changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&io_in_c_bits_source!=source_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel source changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_53&io_in_c_bits_address!=address_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel address changed with multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~reset&_GEN_61[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&~reset&~(_GEN_62[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_57&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_57&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_54&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_55 ? _d_clr_wo_ready_T[18:0]:19'h0)|a_set_wo_ready==19'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==19'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~reset&_GEN_63[0])
            begin 
              if (1)$display("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&~reset&~(_GEN_64[0]|same_cycle_resp_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&same_cycle_resp_1&~reset&io_in_d_bits_size!=io_in_c_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&~same_cycle_resp_1&~reset&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&c_first_1&io_in_c_valid&io_in_c_bits_source==io_in_d_bits_source&d_release_ack&~(io_in_c_bits_opcode==3'h4|io_in_c_bits_opcode==3'h5)&~reset&~(~io_in_d_ready|io_in_c_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if ((|c_set_wo_ready)&~reset&c_set_wo_ready==(_GEN_60 ? _d_clr_wo_ready_T_1[18:0]:19'h0))
            begin 
              if (1)$display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==19'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~reset&_GEN_65[0])
            begin 
              if (1)$display("Assertion failed: 'D' channel re-used a sink ID (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_e_valid&~reset&~(_GEN_66[0]))
            begin 
              if (1)$display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/BankedL2Params.scala:60:27)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_67={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_67 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_67 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_67 ;  
   wire [12:0] _d_first_beats1_decode_T_13=13'h3F<<_GEN_67 ;  
   wire [12:0] _c_first_beats1_decode_T_1=13'h3F<<_GEN_0 ;  
   wire [12:0] _c_first_beats1_decode_T_5=13'h3F<<_GEN_0 ;  
   wire [258:0] _GEN_68={252'h0,io_in_a_bits_source,2'h0} ;  
   wire _GEN_69=_d_first_T_3&d_first_1&~d_release_ack ;  
   wire [270:0] _GEN_70={264'h0,io_in_d_bits_source,2'h0} ;  
   wire _GEN_71=_d_first_T_3&d_first_2&d_release_ack ;  
   wire [31:0] _d_clr_T=32'h1<<_GEN_4 ;  
   wire [31:0] _a_set_T=32'h1<<_GEN_2 ;  
   wire [270:0] _d_opcodes_clr_T_5=271'hF<<_GEN_70 ;  
   wire [258:0] _a_opcodes_set_T_1={255'h0,_GEN_3 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_68 ;  
   wire [270:0] _d_sizes_clr_T_5=271'hF<<_GEN_70 ;  
   wire [258:0] _a_sizes_set_T_1={255'h0,_GEN_3 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_68 ;  
   wire [31:0] _d_clr_T_1=32'h1<<_GEN_4 ;  
   wire [31:0] _c_set_T=32'h1<<_GEN_6 ;  
   wire [270:0] _d_sizes_clr_T_11=271'hF<<_GEN_70 ;  
   wire [258:0] _c_sizes_set_T_1={255'h0,_GEN_7 ? {io_in_c_bits_size,1'h1}:4'h0}<<{252'h0,io_in_c_bits_source,2'h0} ;  
   wire b_first_done=io_in_b_ready&io_in_b_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              b_first_counter <=3'h0;
              c_first_counter <=3'h0;
              inflight <=19'h0;
              inflight_opcodes <=76'h0;
              inflight_sizes <=76'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=19'h0;
              inflight_sizes_1 <=76'h0;
              c_first_counter_1 <=3'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
              inflight_2 <=4'h0;
              d_first_counter_3 <=3'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_3)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   if (d_first_3)
                      d_first_counter_3 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_13[5:3]):3'h0;
                    else 
                      d_first_counter_3 <=d_first_counter_3-3'h1;
                 end 
              if (b_first_done)
                 begin 
                   if (|b_first_counter)
                      b_first_counter <=b_first_counter-3'h1;
                    else 
                      b_first_counter <=3'h0;
                 end 
              if (_c_first_T_1)
                 begin 
                   if (|c_first_counter)
                      c_first_counter <=c_first_counter-3'h1;
                    else 
                      c_first_counter <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_1[5:3]):3'h0;
                   if (c_first_1)
                      c_first_counter_1 <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      c_first_counter_1 <=c_first_counter_1-3'h1;
                 end 
              inflight <=(inflight|(_GEN_3 ? _a_set_T[18:0]:19'h0))&~(_GEN_69 ? _d_clr_T[18:0]:19'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_3 ? _a_opcodes_set_T_1[75:0]:76'h0))&~(_GEN_69 ? _d_opcodes_clr_T_5[75:0]:76'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_3 ? _a_sizes_set_T_1[75:0]:76'h0))&~(_GEN_69 ? _d_sizes_clr_T_5[75:0]:76'h0);
              if (_a_first_T_1|_d_first_T_3)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=(inflight_1|(_GEN_7 ? _c_set_T[18:0]:19'h0))&~(_GEN_71 ? _d_clr_T_1[18:0]:19'h0);
              inflight_sizes_1 <=(inflight_sizes_1|(_GEN_7 ? _c_sizes_set_T_1[75:0]:76'h0))&~(_GEN_71 ? _d_sizes_clr_T_11[75:0]:76'h0);
              if (_c_first_T_1|_d_first_T_3)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight_2 <=(inflight_2|d_set)&~(io_in_e_valid ? 4'h1<<_GEN_10:4'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_3&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
         if (b_first_done&~(|b_first_counter))
            begin 
              param_2 <=io_in_b_bits_param;
              address_1 <=io_in_b_bits_address;
            end 
         if (_c_first_T_1&~(|c_first_counter))
            begin 
              opcode_3 <=io_in_c_bits_opcode;
              param_3 <=io_in_c_bits_param;
              size_3 <=io_in_c_bits_size;
              source_3 <=io_in_c_bits_source;
              address_2 <=io_in_c_bits_address;
            end 
       end
  
endmodule
 
module BroadcastFilter (
  output io_request_ready,
  input io_request_valid,
  input [1:0] io_request_bits_mshr,
  input [31:0] io_request_bits_address,
  input io_request_bits_allocOH,
  input io_request_bits_needT,
  input io_response_ready,
  output io_response_valid,
  output [1:0] io_response_bits_mshr,
  output [31:0] io_response_bits_address,
  output io_response_bits_allocOH,
  output io_response_bits_needT) ; 
  assign io_request_ready=io_response_ready; 
  assign io_response_valid=io_request_valid; 
  assign io_response_bits_mshr=io_request_bits_mshr; 
  assign io_response_bits_address=io_request_bits_address; 
  assign io_response_bits_allocOH=io_request_bits_allocOH; 
  assign io_response_bits_needT=io_request_bits_needT; 
endmodule
 
module ram_8x72 (
  input [2:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [71:0] R0_data,
  input [2:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [71:0] W0_data) ; 
   reg [71:0] Memory[0:7] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:72'bx; 
endmodule
 
module Queue_74 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [7:0] io_enq_bits_mask,
  input [63:0] io_enq_bits_data,
  input io_deq_ready,
  output io_deq_valid,
  output [7:0] io_deq_bits_mask,
  output [63:0] io_deq_bits_data) ; 
   wire [71:0] _ram_ext_R0_data ;  
   reg [2:0] enq_ptr_value ;  
   reg [2:0] deq_ptr_value ;  
   reg maybe_full ;  
   wire ptr_match=enq_ptr_value==deq_ptr_value ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              enq_ptr_value <=3'h0;
              deq_ptr_value <=3'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 enq_ptr_value <=enq_ptr_value+3'h1;
              if (do_deq)
                 deq_ptr_value <=deq_ptr_value+3'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_8x72 ram_ext(.R0_addr(deq_ptr_value),.R0_en(1'h1),.R0_clk(clock),.R0_data(_ram_ext_R0_data),.W0_addr(enq_ptr_value),.W0_en(do_enq),.W0_clk(clock),.W0_data({io_enq_bits_data,io_enq_bits_mask})); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
  assign io_deq_bits_mask=_ram_ext_R0_data[7:0]; 
  assign io_deq_bits_data=_ram_ext_R0_data[71:8]; 
endmodule
 
module TLBroadcastTracker (
  input clock,
  input reset,
  input io_in_a_first,
  output io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input [63:0] io_in_a_bits_data,
  input io_out_a_ready,
  output io_out_a_valid,
  output [2:0] io_out_a_bits_opcode,
  output [2:0] io_out_a_bits_param,
  output [2:0] io_out_a_bits_size,
  output [6:0] io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output [7:0] io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input io_probe_valid,
  input io_probe_bits_count,
  input io_probenack,
  input io_probedack,
  input io_probesack,
  input io_d_last,
  input io_e_last,
  output [4:0] io_source,
  output [25:0] io_line,
  output io_idle,
  output io_need_d) ; 
   wire io_in_a_ready_0 ;  
   wire _o_data_q_io_enq_ready ;  
   wire _o_data_q_io_deq_valid ;  
   reg got_e ;  
   reg sent_d ;  
   reg shared ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [31:0] address ;  
   reg count ;  
   wire idle=got_e&sent_d ;  
   wire _GEN=io_in_a_ready_0&io_in_a_valid&io_in_a_first ;  
   wire _GEN_0=io_probenack|io_probedack ;  
  always @( posedge clock)
       begin 
         if (_GEN&~reset&~idle)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:439 assert (idle)\n");
              if (1)$display("");
            end 
         if (io_d_last&~reset&sent_d)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n");
              if (1)$display("");
            end 
         if (io_e_last&~reset&got_e)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&~count)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n");
              if (1)$display("");
            end 
       end
  
  assign io_in_a_ready_0=(idle|~io_in_a_first)&_o_data_q_io_enq_ready; 
   wire acquire=opcode==3'h6|(&opcode) ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              got_e <=1'h1;
              sent_d <=1'h1;
              address <=32'h0;
            end 
          else 
            begin 
              got_e <=io_e_last|(_GEN ? io_in_a_bits_opcode!=3'h6&io_in_a_bits_opcode!=3'h7:got_e);
              sent_d <=io_d_last|~_GEN&sent_d;
              if (_GEN)
                 address <=io_in_a_bits_address;
            end 
         if (io_probesack)
            shared <=1'h1;
          else 
            shared <=~_GEN&shared;
         if (_GEN)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
            end 
         if (_GEN_0)
            count <=count-~(io_probenack&io_probedack);
          else 
            if (io_probe_valid)
               count <=io_probe_bits_count;
             else 
               count <=_GEN|count;
       end
  
  Queue_74 o_data_q(.clock(clock),.reset(reset),.io_enq_ready(_o_data_q_io_enq_ready),.io_enq_valid((idle|~io_in_a_first)&io_in_a_valid),.io_enq_bits_mask(io_in_a_bits_mask),.io_enq_bits_data(io_in_a_bits_data),.io_deq_ready(io_out_a_ready&~count),.io_deq_valid(_o_data_q_io_deq_valid),.io_deq_bits_mask(io_out_a_bits_mask),.io_deq_bits_data(io_out_a_bits_data)); 
  assign io_in_a_ready=io_in_a_ready_0; 
  assign io_out_a_valid=_o_data_q_io_deq_valid&~count; 
  assign io_out_a_bits_opcode=acquire ? 3'h4:opcode; 
  assign io_out_a_bits_param=acquire ? 3'h0:param; 
  assign io_out_a_bits_size=size; 
  assign io_out_a_bits_source={acquire ? {1'h1,~shared}:2'h0,source}; 
  assign io_out_a_bits_address=address; 
  assign io_source=source; 
  assign io_line=address[31:6]; 
  assign io_idle=idle; 
  assign io_need_d=~sent_d; 
endmodule
 
module TLBroadcastTracker_1 (
  input clock,
  input reset,
  input io_in_a_first,
  output io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input [63:0] io_in_a_bits_data,
  input io_out_a_ready,
  output io_out_a_valid,
  output [2:0] io_out_a_bits_opcode,
  output [2:0] io_out_a_bits_param,
  output [2:0] io_out_a_bits_size,
  output [6:0] io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output [7:0] io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input io_probe_valid,
  input io_probe_bits_count,
  input io_probenack,
  input io_probedack,
  input io_probesack,
  input io_d_last,
  input io_e_last,
  output [4:0] io_source,
  output [25:0] io_line,
  output io_idle,
  output io_need_d) ; 
   wire io_in_a_ready_0 ;  
   wire _o_data_q_io_enq_ready ;  
   wire _o_data_q_io_deq_valid ;  
   reg got_e ;  
   reg sent_d ;  
   reg shared ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [31:0] address ;  
   reg count ;  
   wire idle=got_e&sent_d ;  
   wire _GEN=io_in_a_ready_0&io_in_a_valid&io_in_a_first ;  
   wire _GEN_0=io_probenack|io_probedack ;  
  always @( posedge clock)
       begin 
         if (_GEN&~reset&~idle)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:439 assert (idle)\n");
              if (1)$display("");
            end 
         if (io_d_last&~reset&sent_d)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n");
              if (1)$display("");
            end 
         if (io_e_last&~reset&got_e)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&~count)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n");
              if (1)$display("");
            end 
       end
  
  assign io_in_a_ready_0=(idle|~io_in_a_first)&_o_data_q_io_enq_ready; 
   wire acquire=opcode==3'h6|(&opcode) ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              got_e <=1'h1;
              sent_d <=1'h1;
              address <=32'h40;
            end 
          else 
            begin 
              got_e <=io_e_last|(_GEN ? io_in_a_bits_opcode!=3'h6&io_in_a_bits_opcode!=3'h7:got_e);
              sent_d <=io_d_last|~_GEN&sent_d;
              if (_GEN)
                 address <=io_in_a_bits_address;
            end 
         if (io_probesack)
            shared <=1'h1;
          else 
            shared <=~_GEN&shared;
         if (_GEN)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
            end 
         if (_GEN_0)
            count <=count-~(io_probenack&io_probedack);
          else 
            if (io_probe_valid)
               count <=io_probe_bits_count;
             else 
               count <=_GEN|count;
       end
  
  Queue_74 o_data_q(.clock(clock),.reset(reset),.io_enq_ready(_o_data_q_io_enq_ready),.io_enq_valid((idle|~io_in_a_first)&io_in_a_valid),.io_enq_bits_mask(io_in_a_bits_mask),.io_enq_bits_data(io_in_a_bits_data),.io_deq_ready(io_out_a_ready&~count),.io_deq_valid(_o_data_q_io_deq_valid),.io_deq_bits_mask(io_out_a_bits_mask),.io_deq_bits_data(io_out_a_bits_data)); 
  assign io_in_a_ready=io_in_a_ready_0; 
  assign io_out_a_valid=_o_data_q_io_deq_valid&~count; 
  assign io_out_a_bits_opcode=acquire ? 3'h4:opcode; 
  assign io_out_a_bits_param=acquire ? 3'h0:param; 
  assign io_out_a_bits_size=size; 
  assign io_out_a_bits_source={acquire ? {1'h1,~shared}:2'h0,source}; 
  assign io_out_a_bits_address=address; 
  assign io_source=source; 
  assign io_line=address[31:6]; 
  assign io_idle=idle; 
  assign io_need_d=~sent_d; 
endmodule
 
module TLBroadcastTracker_2 (
  input clock,
  input reset,
  input io_in_a_first,
  output io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input [63:0] io_in_a_bits_data,
  input io_out_a_ready,
  output io_out_a_valid,
  output [2:0] io_out_a_bits_opcode,
  output [2:0] io_out_a_bits_param,
  output [2:0] io_out_a_bits_size,
  output [6:0] io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output [7:0] io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input io_probe_valid,
  input io_probe_bits_count,
  input io_probenack,
  input io_probedack,
  input io_probesack,
  input io_d_last,
  input io_e_last,
  output [4:0] io_source,
  output [25:0] io_line,
  output io_idle,
  output io_need_d) ; 
   wire io_in_a_ready_0 ;  
   wire _o_data_q_io_enq_ready ;  
   wire _o_data_q_io_deq_valid ;  
   reg got_e ;  
   reg sent_d ;  
   reg shared ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [31:0] address ;  
   reg count ;  
   wire idle=got_e&sent_d ;  
   wire _GEN=io_in_a_ready_0&io_in_a_valid&io_in_a_first ;  
   wire _GEN_0=io_probenack|io_probedack ;  
  always @( posedge clock)
       begin 
         if (_GEN&~reset&~idle)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:439 assert (idle)\n");
              if (1)$display("");
            end 
         if (io_d_last&~reset&sent_d)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n");
              if (1)$display("");
            end 
         if (io_e_last&~reset&got_e)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&~count)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n");
              if (1)$display("");
            end 
       end
  
  assign io_in_a_ready_0=(idle|~io_in_a_first)&_o_data_q_io_enq_ready; 
   wire acquire=opcode==3'h6|(&opcode) ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              got_e <=1'h1;
              sent_d <=1'h1;
              address <=32'h80;
            end 
          else 
            begin 
              got_e <=io_e_last|(_GEN ? io_in_a_bits_opcode!=3'h6&io_in_a_bits_opcode!=3'h7:got_e);
              sent_d <=io_d_last|~_GEN&sent_d;
              if (_GEN)
                 address <=io_in_a_bits_address;
            end 
         if (io_probesack)
            shared <=1'h1;
          else 
            shared <=~_GEN&shared;
         if (_GEN)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
            end 
         if (_GEN_0)
            count <=count-~(io_probenack&io_probedack);
          else 
            if (io_probe_valid)
               count <=io_probe_bits_count;
             else 
               count <=_GEN|count;
       end
  
  Queue_74 o_data_q(.clock(clock),.reset(reset),.io_enq_ready(_o_data_q_io_enq_ready),.io_enq_valid((idle|~io_in_a_first)&io_in_a_valid),.io_enq_bits_mask(io_in_a_bits_mask),.io_enq_bits_data(io_in_a_bits_data),.io_deq_ready(io_out_a_ready&~count),.io_deq_valid(_o_data_q_io_deq_valid),.io_deq_bits_mask(io_out_a_bits_mask),.io_deq_bits_data(io_out_a_bits_data)); 
  assign io_in_a_ready=io_in_a_ready_0; 
  assign io_out_a_valid=_o_data_q_io_deq_valid&~count; 
  assign io_out_a_bits_opcode=acquire ? 3'h4:opcode; 
  assign io_out_a_bits_param=acquire ? 3'h0:param; 
  assign io_out_a_bits_size=size; 
  assign io_out_a_bits_source={acquire ? {1'h1,~shared}:2'h0,source}; 
  assign io_out_a_bits_address=address; 
  assign io_source=source; 
  assign io_line=address[31:6]; 
  assign io_idle=idle; 
  assign io_need_d=~sent_d; 
endmodule
 
module TLBroadcastTracker_3 (
  input clock,
  input reset,
  input io_in_a_first,
  output io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [4:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input [63:0] io_in_a_bits_data,
  input io_out_a_ready,
  output io_out_a_valid,
  output [2:0] io_out_a_bits_opcode,
  output [2:0] io_out_a_bits_param,
  output [2:0] io_out_a_bits_size,
  output [6:0] io_out_a_bits_source,
  output [31:0] io_out_a_bits_address,
  output [7:0] io_out_a_bits_mask,
  output [63:0] io_out_a_bits_data,
  input io_probe_valid,
  input io_probe_bits_count,
  input io_probenack,
  input io_probedack,
  input io_probesack,
  input io_d_last,
  input io_e_last,
  output [4:0] io_source,
  output [25:0] io_line,
  output io_idle,
  output io_need_d) ; 
   wire io_in_a_ready_0 ;  
   wire _o_data_q_io_enq_ready ;  
   wire _o_data_q_io_deq_valid ;  
   reg got_e ;  
   reg sent_d ;  
   reg shared ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [4:0] source ;  
   reg [31:0] address ;  
   reg count ;  
   wire idle=got_e&sent_d ;  
   wire _GEN=io_in_a_ready_0&io_in_a_valid&io_in_a_first ;  
   wire _GEN_0=io_probenack|io_probedack ;  
  always @( posedge clock)
       begin 
         if (_GEN&~reset&~idle)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:439 assert (idle)\n");
              if (1)$display("");
            end 
         if (io_d_last&~reset&sent_d)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:460 assert (!sent_d)\n");
              if (1)$display("");
            end 
         if (io_e_last&~reset&got_e)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:464 assert (!got_e)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&~count)
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:469 assert (count > 0.U)\n");
              if (1)$display("");
            end 
       end
  
  assign io_in_a_ready_0=(idle|~io_in_a_first)&_o_data_q_io_enq_ready; 
   wire acquire=opcode==3'h6|(&opcode) ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              got_e <=1'h1;
              sent_d <=1'h1;
              address <=32'hC0;
            end 
          else 
            begin 
              got_e <=io_e_last|(_GEN ? io_in_a_bits_opcode!=3'h6&io_in_a_bits_opcode!=3'h7:got_e);
              sent_d <=io_d_last|~_GEN&sent_d;
              if (_GEN)
                 address <=io_in_a_bits_address;
            end 
         if (io_probesack)
            shared <=1'h1;
          else 
            shared <=~_GEN&shared;
         if (_GEN)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
            end 
         if (_GEN_0)
            count <=count-~(io_probenack&io_probedack);
          else 
            if (io_probe_valid)
               count <=io_probe_bits_count;
             else 
               count <=_GEN|count;
       end
  
  Queue_74 o_data_q(.clock(clock),.reset(reset),.io_enq_ready(_o_data_q_io_enq_ready),.io_enq_valid((idle|~io_in_a_first)&io_in_a_valid),.io_enq_bits_mask(io_in_a_bits_mask),.io_enq_bits_data(io_in_a_bits_data),.io_deq_ready(io_out_a_ready&~count),.io_deq_valid(_o_data_q_io_deq_valid),.io_deq_bits_mask(io_out_a_bits_mask),.io_deq_bits_data(io_out_a_bits_data)); 
  assign io_in_a_ready=io_in_a_ready_0; 
  assign io_out_a_valid=_o_data_q_io_deq_valid&~count; 
  assign io_out_a_bits_opcode=acquire ? 3'h4:opcode; 
  assign io_out_a_bits_param=acquire ? 3'h0:param; 
  assign io_out_a_bits_size=size; 
  assign io_out_a_bits_source={acquire ? {1'h1,~shared}:2'h0,source}; 
  assign io_out_a_bits_address=address; 
  assign io_source=source; 
  assign io_line=address[31:6]; 
  assign io_idle=idle; 
  assign io_need_d=~sent_d; 
endmodule
 
module TLBroadcast (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [4:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [1:0] auto_in_b_bits_param,
  output [31:0] auto_in_b_bits_address,
  output auto_in_c_ready,
  input auto_in_c_valid,
  input [2:0] auto_in_c_bits_opcode,
  input [2:0] auto_in_c_bits_param,
  input [2:0] auto_in_c_bits_size,
  input [4:0] auto_in_c_bits_source,
  input [31:0] auto_in_c_bits_address,
  input [63:0] auto_in_c_bits_data,
  input auto_in_c_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [2:0] auto_in_d_bits_size,
  output [4:0] auto_in_d_bits_source,
  output [1:0] auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_in_e_valid,
  input [1:0] auto_in_e_bits_sink,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [2:0] auto_out_a_bits_size,
  output [6:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [2:0] auto_out_d_bits_size,
  input [6:0] auto_out_d_bits_source,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
   reg [2:0] a_first_counter ;  
   reg probe_todo ;  
   wire putfull_ready ;  
   wire d_normal_ready ;  
   wire releaseack_ready ;  
   wire nodeIn_c_ready ;  
   wire [2:0] d_normal_bits_opcode ;  
   wire [4:0] d_normal_bits_source ;  
   wire d_normal_valid ;  
   wire _TLBroadcastTracker_3_io_in_a_ready ;  
   wire _TLBroadcastTracker_3_io_out_a_valid ;  
   wire [2:0] _TLBroadcastTracker_3_io_out_a_bits_opcode ;  
   wire [2:0] _TLBroadcastTracker_3_io_out_a_bits_param ;  
   wire [2:0] _TLBroadcastTracker_3_io_out_a_bits_size ;  
   wire [6:0] _TLBroadcastTracker_3_io_out_a_bits_source ;  
   wire [31:0] _TLBroadcastTracker_3_io_out_a_bits_address ;  
   wire [7:0] _TLBroadcastTracker_3_io_out_a_bits_mask ;  
   wire [63:0] _TLBroadcastTracker_3_io_out_a_bits_data ;  
   wire [4:0] _TLBroadcastTracker_3_io_source ;  
   wire [25:0] _TLBroadcastTracker_3_io_line ;  
   wire _TLBroadcastTracker_3_io_idle ;  
   wire _TLBroadcastTracker_3_io_need_d ;  
   wire _TLBroadcastTracker_2_io_in_a_ready ;  
   wire _TLBroadcastTracker_2_io_out_a_valid ;  
   wire [2:0] _TLBroadcastTracker_2_io_out_a_bits_opcode ;  
   wire [2:0] _TLBroadcastTracker_2_io_out_a_bits_param ;  
   wire [2:0] _TLBroadcastTracker_2_io_out_a_bits_size ;  
   wire [6:0] _TLBroadcastTracker_2_io_out_a_bits_source ;  
   wire [31:0] _TLBroadcastTracker_2_io_out_a_bits_address ;  
   wire [7:0] _TLBroadcastTracker_2_io_out_a_bits_mask ;  
   wire [63:0] _TLBroadcastTracker_2_io_out_a_bits_data ;  
   wire [4:0] _TLBroadcastTracker_2_io_source ;  
   wire [25:0] _TLBroadcastTracker_2_io_line ;  
   wire _TLBroadcastTracker_2_io_idle ;  
   wire _TLBroadcastTracker_2_io_need_d ;  
   wire _TLBroadcastTracker_1_io_in_a_ready ;  
   wire _TLBroadcastTracker_1_io_out_a_valid ;  
   wire [2:0] _TLBroadcastTracker_1_io_out_a_bits_opcode ;  
   wire [2:0] _TLBroadcastTracker_1_io_out_a_bits_param ;  
   wire [2:0] _TLBroadcastTracker_1_io_out_a_bits_size ;  
   wire [6:0] _TLBroadcastTracker_1_io_out_a_bits_source ;  
   wire [31:0] _TLBroadcastTracker_1_io_out_a_bits_address ;  
   wire [7:0] _TLBroadcastTracker_1_io_out_a_bits_mask ;  
   wire [63:0] _TLBroadcastTracker_1_io_out_a_bits_data ;  
   wire [4:0] _TLBroadcastTracker_1_io_source ;  
   wire [25:0] _TLBroadcastTracker_1_io_line ;  
   wire _TLBroadcastTracker_1_io_idle ;  
   wire _TLBroadcastTracker_1_io_need_d ;  
   wire _TLBroadcastTracker_io_in_a_ready ;  
   wire _TLBroadcastTracker_io_out_a_valid ;  
   wire [2:0] _TLBroadcastTracker_io_out_a_bits_opcode ;  
   wire [2:0] _TLBroadcastTracker_io_out_a_bits_param ;  
   wire [2:0] _TLBroadcastTracker_io_out_a_bits_size ;  
   wire [6:0] _TLBroadcastTracker_io_out_a_bits_source ;  
   wire [31:0] _TLBroadcastTracker_io_out_a_bits_address ;  
   wire [7:0] _TLBroadcastTracker_io_out_a_bits_mask ;  
   wire [63:0] _TLBroadcastTracker_io_out_a_bits_data ;  
   wire [4:0] _TLBroadcastTracker_io_source ;  
   wire [25:0] _TLBroadcastTracker_io_line ;  
   wire _TLBroadcastTracker_io_idle ;  
   wire _TLBroadcastTracker_io_need_d ;  
   wire _filter_io_request_ready ;  
   wire _filter_io_response_valid ;  
   wire [1:0] _filter_io_response_bits_mshr ;  
   wire [31:0] _filter_io_response_bits_address ;  
   wire _filter_io_response_bits_allocOH ;  
   wire _filter_io_response_bits_needT ;  
   wire d_drop=auto_out_d_bits_source[6:5]==2'h1 ;  
   wire _GEN=d_normal_ready&d_normal_valid ;  
   wire [12:0] _GEN_0={10'h0,auto_out_d_bits_size} ;  
   wire [12:0] _beats1_decode_T_1=13'h3F<<_GEN_0 ;  
   wire [2:0] beats1=d_normal_bits_opcode[0] ? ~(_beats1_decode_T_1[5:3]):3'h0 ;  
   reg [2:0] counter ;  
   wire d_first=counter==3'h0 ;  
   wire d_last=counter==3'h1|beats1==3'h0 ;  
   wire [3:0] _d_trackerOH_T_8={_TLBroadcastTracker_3_io_need_d&_TLBroadcastTracker_3_io_source==d_normal_bits_source,_TLBroadcastTracker_2_io_need_d&_TLBroadcastTracker_2_io_source==d_normal_bits_source,_TLBroadcastTracker_1_io_need_d&_TLBroadcastTracker_1_io_source==d_normal_bits_source,_TLBroadcastTracker_io_need_d&_TLBroadcastTracker_io_source==d_normal_bits_source} ;  
   reg [3:0] d_trackerOH_r ;  
   wire [3:0] d_trackerOH=d_first ? _d_trackerOH_T_8:d_trackerOH_r ;  
   wire nodeOut_d_ready=d_normal_ready|d_drop ;  
  assign d_normal_valid=auto_out_d_valid&~d_drop; 
  assign d_normal_bits_source=auto_out_d_bits_source[4:0]; 
  assign d_normal_bits_opcode=auto_out_d_bits_source[6] ? (auto_out_d_bits_opcode[0] ? 3'h5:3'h6):auto_out_d_bits_opcode; 
   wire d_response=auto_out_d_bits_opcode[0]|~(auto_out_d_bits_source[6]) ;  
   wire _GEN_1=nodeOut_d_ready&auto_out_d_valid ;  
   wire c_probeack=auto_in_c_bits_opcode==3'h4 ;  
   wire c_probeackdata=auto_in_c_bits_opcode==3'h5 ;  
   wire c_release=auto_in_c_bits_opcode==3'h6 ;  
   wire c_trackerOH_0=_TLBroadcastTracker_io_line==auto_in_c_bits_address[31:6] ;  
   wire c_trackerOH_1=_TLBroadcastTracker_1_io_line==auto_in_c_bits_address[31:6] ;  
   wire c_trackerOH_2=_TLBroadcastTracker_2_io_line==auto_in_c_bits_address[31:6] ;  
   wire c_trackerOH_3=_TLBroadcastTracker_3_io_line==auto_in_c_bits_address[31:6] ;  
   wire _c_first_T=nodeIn_c_ready&auto_in_c_valid ;  
   wire _clearOH_T_1=c_probeack|c_probeackdata ;  
   wire _GEN_2=_c_first_T&c_probeack ;  
   wire _GEN_3=auto_in_c_bits_param==3'h0|auto_in_c_bits_param==3'h4 ;  
  assign nodeIn_c_ready=c_probeack|(c_release ? releaseack_ready:putfull_ready); 
   wire winner_0=auto_in_c_valid&c_release ;  
   wire putfull_valid=auto_in_c_valid&(c_probeackdata|(&auto_in_c_bits_opcode)) ;  
   wire _putfull_bits_a_mask_T=auto_in_c_bits_size>3'h2 ;  
   wire putfull_bits_a_mask_size=auto_in_c_bits_size[1:0]==2'h2 ;  
   wire putfull_bits_a_mask_acc=_putfull_bits_a_mask_T|putfull_bits_a_mask_size&~(auto_in_c_bits_address[2]) ;  
   wire putfull_bits_a_mask_acc_1=_putfull_bits_a_mask_T|putfull_bits_a_mask_size&auto_in_c_bits_address[2] ;  
   wire putfull_bits_a_mask_size_1=auto_in_c_bits_size[1:0]==2'h1 ;  
   wire putfull_bits_a_mask_eq_2=~(auto_in_c_bits_address[2])&~(auto_in_c_bits_address[1]) ;  
   wire putfull_bits_a_mask_acc_2=putfull_bits_a_mask_acc|putfull_bits_a_mask_size_1&putfull_bits_a_mask_eq_2 ;  
   wire putfull_bits_a_mask_eq_3=~(auto_in_c_bits_address[2])&auto_in_c_bits_address[1] ;  
   wire putfull_bits_a_mask_acc_3=putfull_bits_a_mask_acc|putfull_bits_a_mask_size_1&putfull_bits_a_mask_eq_3 ;  
   wire putfull_bits_a_mask_eq_4=auto_in_c_bits_address[2]&~(auto_in_c_bits_address[1]) ;  
   wire putfull_bits_a_mask_acc_4=putfull_bits_a_mask_acc_1|putfull_bits_a_mask_size_1&putfull_bits_a_mask_eq_4 ;  
   wire putfull_bits_a_mask_eq_5=auto_in_c_bits_address[2]&auto_in_c_bits_address[1] ;  
   wire putfull_bits_a_mask_acc_5=putfull_bits_a_mask_acc_1|putfull_bits_a_mask_size_1&putfull_bits_a_mask_eq_5 ;  
   reg [2:0] beatsLeft ;  
   wire idle=beatsLeft==3'h0 ;  
   wire winner_1=~winner_0&d_normal_valid ;  
   wire _nodeIn_d_valid_T=winner_0|d_normal_valid ;  
   reg state_0 ;  
   reg state_1 ;  
   wire muxState_0=idle ? winner_0:state_0 ;  
   wire muxState_1=idle ? winner_1:state_1 ;  
  assign releaseack_ready=auto_in_d_ready&(idle|state_0); 
  assign d_normal_ready=auto_in_d_ready&(idle ? ~winner_0:state_1); 
   wire nodeIn_d_valid=idle ? _nodeIn_d_valid_T:state_0&winner_0|state_1&d_normal_valid ;  
   wire _nodeIn_d_bits_T_2=muxState_1&auto_out_d_bits_corrupt ;  
   wire _nodeIn_d_bits_T_8=muxState_1&auto_out_d_bits_denied ;  
   wire [1:0] _nodeIn_d_bits_T_11=muxState_1 ? {|(d_trackerOH[3:2]),d_trackerOH[3]|d_trackerOH[1]}:2'h0 ;  
   wire [4:0] _nodeIn_d_bits_T_14=(muxState_0 ? auto_in_c_bits_source:5'h0)|(muxState_1 ? d_normal_bits_source:5'h0) ;  
   wire [2:0] _nodeIn_d_bits_T_17=(muxState_0 ? auto_in_c_bits_size:3'h0)|(muxState_1 ? auto_out_d_bits_size:3'h0) ;  
   wire [1:0] _nodeIn_d_bits_T_20=muxState_1&auto_out_d_bits_source[6]&auto_out_d_bits_opcode[0] ? {1'h0,~(auto_out_d_bits_source[5])}:2'h0 ;  
   wire [2:0] _nodeIn_d_bits_T_23=(muxState_0 ? 3'h6:3'h0)|(muxState_1 ? d_normal_bits_opcode:3'h0) ;  
   reg [2:0] beatsLeft_1 ;  
   wire idle_1=beatsLeft_1==3'h0 ;  
   wire _GEN_4=_TLBroadcastTracker_io_out_a_valid|putfull_valid ;  
   wire _GEN_5=_TLBroadcastTracker_2_io_out_a_valid|_TLBroadcastTracker_1_io_out_a_valid|_GEN_4 ;  
   wire _GEN_6=_TLBroadcastTracker_1_io_out_a_valid|_TLBroadcastTracker_io_out_a_valid|putfull_valid ;  
   wire winner_1_1=~putfull_valid&_TLBroadcastTracker_io_out_a_valid ;  
   wire winner_1_2=~_GEN_4&_TLBroadcastTracker_1_io_out_a_valid ;  
   wire winner_1_3=~_GEN_6&_TLBroadcastTracker_2_io_out_a_valid ;  
   wire winner_1_4=~_GEN_5&_TLBroadcastTracker_3_io_out_a_valid ;  
   wire _nodeOut_a_valid_T=putfull_valid|_TLBroadcastTracker_io_out_a_valid ;  
   wire prefixOR_2=putfull_valid|winner_1_1 ;  
   wire prefixOR_3=prefixOR_2|winner_1_2 ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~auto_out_d_valid|~d_drop|auto_out_d_bits_opcode==3'h0))
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:125 assert (!out.d.valid || !d_drop || out.d.bits.opcode === TLMessages.AccessAck)\n");
              if (1)$display("");
            end 
         if (~reset&~(~d_normal_valid|(|d_trackerOH)|d_normal_bits_opcode==3'h6))
            begin 
              if (1)$display("Assertion failed\n    at Broadcast.scala:137 assert (!d_normal.valid || (d_trackerOH.orR || d_normal.bits.opcode === TLMessages.ReleaseAck))\n");
              if (1)$display("");
            end 
         if (~reset&~(~winner_0|~winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_nodeIn_d_valid_T|winner_0|winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
         if (~reset&~((~putfull_valid|~winner_1_1)&(~prefixOR_2|~winner_1_2)&(~prefixOR_3|~winner_1_3)&(~(prefixOR_3|winner_1_3)|~winner_1_4)))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~(_nodeOut_a_valid_T|_TLBroadcastTracker_1_io_out_a_valid|_TLBroadcastTracker_2_io_out_a_valid|_TLBroadcastTracker_3_io_out_a_valid)|putfull_valid|winner_1_1|winner_1_2|winner_1_3|winner_1_4))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg state_1_0 ;  
   reg state_1_1 ;  
   reg state_1_2 ;  
   reg state_1_3 ;  
   reg state_1_4 ;  
   wire muxState_1_0=idle_1 ? putfull_valid:state_1_0 ;  
   wire muxState_1_1=idle_1 ? winner_1_1:state_1_1 ;  
   wire muxState_1_2=idle_1 ? winner_1_2:state_1_2 ;  
   wire muxState_1_3=idle_1 ? winner_1_3:state_1_3 ;  
   wire muxState_1_4=idle_1 ? winner_1_4:state_1_4 ;  
  assign putfull_ready=auto_out_a_ready&(idle_1|state_1_0); 
   wire nodeOut_a_valid=idle_1 ? _nodeOut_a_valid_T|_TLBroadcastTracker_1_io_out_a_valid|_TLBroadcastTracker_2_io_out_a_valid|_TLBroadcastTracker_3_io_out_a_valid:state_1_0&putfull_valid|state_1_1&_TLBroadcastTracker_io_out_a_valid|state_1_2&_TLBroadcastTracker_1_io_out_a_valid|state_1_3&_TLBroadcastTracker_2_io_out_a_valid|state_1_4&_TLBroadcastTracker_3_io_out_a_valid ;  
   reg [25:0] probe_line ;  
   reg [1:0] probe_perms ;  
   wire [31:0] nodeIn_b_bits_b_address={probe_line,6'h0} ;  
   wire _matchTrackers_T_1=_TLBroadcastTracker_io_line==auto_in_a_bits_address[31:6] ;  
   wire _matchTrackers_T_3=_TLBroadcastTracker_1_io_line==auto_in_a_bits_address[31:6] ;  
   wire _matchTrackers_T_5=_TLBroadcastTracker_2_io_line==auto_in_a_bits_address[31:6] ;  
   wire _matchTrackers_T_7=_TLBroadcastTracker_3_io_line==auto_in_a_bits_address[31:6] ;  
   wire [3:0] filter_io_request_bits_mshr_lo=(|{_matchTrackers_T_7,_matchTrackers_T_5,_matchTrackers_T_3,_matchTrackers_T_1}) ? {_matchTrackers_T_7,_matchTrackers_T_5,_matchTrackers_T_3,_matchTrackers_T_1}:{~(_TLBroadcastTracker_2_io_idle|_TLBroadcastTracker_1_io_idle|_TLBroadcastTracker_io_idle),~(_TLBroadcastTracker_1_io_idle|_TLBroadcastTracker_io_idle),~_TLBroadcastTracker_io_idle,1'h1}&{_TLBroadcastTracker_3_io_idle,_TLBroadcastTracker_2_io_idle,_TLBroadcastTracker_1_io_idle,_TLBroadcastTracker_io_idle} ;  
   wire [3:0] _GEN_7=filter_io_request_bits_mshr_lo&{_TLBroadcastTracker_3_io_in_a_ready,_TLBroadcastTracker_2_io_in_a_ready,_TLBroadcastTracker_1_io_in_a_ready,_TLBroadcastTracker_io_in_a_ready} ;  
   wire nodeIn_a_ready=((|a_first_counter)|_filter_io_request_ready)&(|_GEN_7) ;  
   wire _GEN_8=(|a_first_counter)|_filter_io_request_ready ;  
   wire _sack_T=~probe_todo&_filter_io_response_valid ;  
   wire [12:0] _decode_T_5=13'h3F<<_GEN_0 ;  
   wire [12:0] _decode_T_25=13'h3F<<_TLBroadcastTracker_3_io_out_a_bits_size ;  
   wire [12:0] _decode_T_21=13'h3F<<_TLBroadcastTracker_2_io_out_a_bits_size ;  
   wire [12:0] _decode_T_17=13'h3F<<_TLBroadcastTracker_1_io_out_a_bits_size ;  
   wire [12:0] _decode_T_13=13'h3F<<_TLBroadcastTracker_io_out_a_bits_size ;  
   wire [12:0] _decode_T_9=13'h3F<<auto_in_c_bits_size ;  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<auto_in_a_bits_size ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              counter <=3'h0;
              beatsLeft <=3'h0;
              state_0 <=1'h0;
              state_1 <=1'h0;
              beatsLeft_1 <=3'h0;
              state_1_0 <=1'h0;
              state_1_1 <=1'h0;
              state_1_2 <=1'h0;
              state_1_3 <=1'h0;
              state_1_4 <=1'h0;
              probe_todo <=1'h0;
              a_first_counter <=3'h0;
            end 
          else 
            begin 
              if (_GEN)
                 begin 
                   if (d_first)
                      counter <=beats1;
                    else 
                      counter <=counter-3'h1;
                 end 
              if (idle&auto_in_d_ready)
                 beatsLeft <=winner_1&d_normal_bits_opcode[0] ? ~(_decode_T_5[5:3]):3'h0;
               else 
                 beatsLeft <=beatsLeft-{2'h0,auto_in_d_ready&nodeIn_d_valid};
              if (idle)
                 begin 
                   state_0 <=winner_0;
                   state_1 <=winner_1;
                 end 
              if (idle_1&auto_out_a_ready)
                 beatsLeft_1 <=(putfull_valid ? ~(_decode_T_9[5:3]):3'h0)|(winner_1_1&~(_TLBroadcastTracker_io_out_a_bits_opcode[2]) ? ~(_decode_T_13[5:3]):3'h0)|(winner_1_2&~(_TLBroadcastTracker_1_io_out_a_bits_opcode[2]) ? ~(_decode_T_17[5:3]):3'h0)|(winner_1_3&~(_TLBroadcastTracker_2_io_out_a_bits_opcode[2]) ? ~(_decode_T_21[5:3]):3'h0)|(winner_1_4&~(_TLBroadcastTracker_3_io_out_a_bits_opcode[2]) ? ~(_decode_T_25[5:3]):3'h0);
               else 
                 beatsLeft_1 <=beatsLeft_1-{2'h0,auto_out_a_ready&nodeOut_a_valid};
              if (idle_1)
                 begin 
                   state_1_0 <=putfull_valid;
                   state_1_1 <=winner_1_1;
                   state_1_2 <=winner_1_2;
                   state_1_3 <=winner_1_3;
                   state_1_4 <=winner_1_4;
                 end 
              if (_sack_T)
                 probe_todo <=~_filter_io_response_bits_allocOH;
               else 
                 probe_todo <=~(auto_in_b_ready&probe_todo)&probe_todo;
              if (nodeIn_a_ready&auto_in_a_valid)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=auto_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                 end 
            end 
         if (d_first)
            d_trackerOH_r <=_d_trackerOH_T_8;
         if (_sack_T)
            begin 
              probe_line <=_filter_io_response_bits_address[31:6];
              probe_perms <=_filter_io_response_bits_needT ? 2'h2:2'h1;
            end 
       end
  
  TLMonitor_21 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_b_ready(auto_in_b_ready),.io_in_b_valid(probe_todo),.io_in_b_bits_param(probe_perms),.io_in_b_bits_address(nodeIn_b_bits_b_address),.io_in_c_ready(nodeIn_c_ready),.io_in_c_valid(auto_in_c_valid),.io_in_c_bits_opcode(auto_in_c_bits_opcode),.io_in_c_bits_param(auto_in_c_bits_param),.io_in_c_bits_size(auto_in_c_bits_size),.io_in_c_bits_source(auto_in_c_bits_source),.io_in_c_bits_address(auto_in_c_bits_address),.io_in_c_bits_corrupt(auto_in_c_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(_nodeIn_d_bits_T_23),.io_in_d_bits_param(_nodeIn_d_bits_T_20),.io_in_d_bits_size(_nodeIn_d_bits_T_17),.io_in_d_bits_source(_nodeIn_d_bits_T_14),.io_in_d_bits_sink(_nodeIn_d_bits_T_11),.io_in_d_bits_denied(_nodeIn_d_bits_T_8),.io_in_d_bits_corrupt(_nodeIn_d_bits_T_2),.io_in_e_valid(auto_in_e_valid),.io_in_e_bits_sink(auto_in_e_bits_sink)); 
  BroadcastFilter filter(.io_request_ready(_filter_io_request_ready),.io_request_valid(auto_in_a_valid&~(|a_first_counter)&(|_GEN_7)),.io_request_bits_mshr({|(filter_io_request_bits_mshr_lo[3:2]),filter_io_request_bits_mshr_lo[3]|filter_io_request_bits_mshr_lo[1]}),.io_request_bits_address(auto_in_a_bits_address),.io_request_bits_allocOH(auto_in_a_bits_source==5'h10),.io_request_bits_needT((&auto_in_a_bits_opcode)|auto_in_a_bits_opcode==3'h6 ? auto_in_a_bits_param==3'h2|auto_in_a_bits_param==3'h1:auto_in_a_bits_opcode==3'h5 ? auto_in_a_bits_param==3'h1:auto_in_a_bits_opcode!=3'h4),.io_response_ready(~probe_todo),.io_response_valid(_filter_io_response_valid),.io_response_bits_mshr(_filter_io_response_bits_mshr),.io_response_bits_address(_filter_io_response_bits_address),.io_response_bits_allocOH(_filter_io_response_bits_allocOH),.io_response_bits_needT(_filter_io_response_bits_needT)); 
  TLBroadcastTracker TLBroadcastTracker(.clock(clock),.reset(reset),.io_in_a_first(~(|a_first_counter)),.io_in_a_ready(_TLBroadcastTracker_io_in_a_ready),.io_in_a_valid(auto_in_a_valid&filter_io_request_bits_mshr_lo[0]&_GEN_8),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_data(auto_in_a_bits_data),.io_out_a_ready(auto_out_a_ready&(idle_1 ? ~putfull_valid:state_1_1)),.io_out_a_valid(_TLBroadcastTracker_io_out_a_valid),.io_out_a_bits_opcode(_TLBroadcastTracker_io_out_a_bits_opcode),.io_out_a_bits_param(_TLBroadcastTracker_io_out_a_bits_param),.io_out_a_bits_size(_TLBroadcastTracker_io_out_a_bits_size),.io_out_a_bits_source(_TLBroadcastTracker_io_out_a_bits_source),.io_out_a_bits_address(_TLBroadcastTracker_io_out_a_bits_address),.io_out_a_bits_mask(_TLBroadcastTracker_io_out_a_bits_mask),.io_out_a_bits_data(_TLBroadcastTracker_io_out_a_bits_data),.io_probe_valid(_sack_T&_filter_io_response_bits_mshr==2'h0),.io_probe_bits_count(~_filter_io_response_bits_allocOH),.io_probenack(_GEN_2&c_trackerOH_0),.io_probedack(d_trackerOH[0]&_GEN_1&d_drop),.io_probesack(_c_first_T&c_trackerOH_0&_clearOH_T_1&_GEN_3),.io_d_last(d_trackerOH[0]&_GEN&d_response&d_last),.io_e_last(auto_in_e_bits_sink==2'h0&auto_in_e_valid),.io_source(_TLBroadcastTracker_io_source),.io_line(_TLBroadcastTracker_io_line),.io_idle(_TLBroadcastTracker_io_idle),.io_need_d(_TLBroadcastTracker_io_need_d)); 
  TLBroadcastTracker_1 TLBroadcastTracker_1(.clock(clock),.reset(reset),.io_in_a_first(~(|a_first_counter)),.io_in_a_ready(_TLBroadcastTracker_1_io_in_a_ready),.io_in_a_valid(auto_in_a_valid&filter_io_request_bits_mshr_lo[1]&_GEN_8),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_data(auto_in_a_bits_data),.io_out_a_ready(auto_out_a_ready&(idle_1 ? ~_GEN_4:state_1_2)),.io_out_a_valid(_TLBroadcastTracker_1_io_out_a_valid),.io_out_a_bits_opcode(_TLBroadcastTracker_1_io_out_a_bits_opcode),.io_out_a_bits_param(_TLBroadcastTracker_1_io_out_a_bits_param),.io_out_a_bits_size(_TLBroadcastTracker_1_io_out_a_bits_size),.io_out_a_bits_source(_TLBroadcastTracker_1_io_out_a_bits_source),.io_out_a_bits_address(_TLBroadcastTracker_1_io_out_a_bits_address),.io_out_a_bits_mask(_TLBroadcastTracker_1_io_out_a_bits_mask),.io_out_a_bits_data(_TLBroadcastTracker_1_io_out_a_bits_data),.io_probe_valid(_sack_T&_filter_io_response_bits_mshr==2'h1),.io_probe_bits_count(~_filter_io_response_bits_allocOH),.io_probenack(_GEN_2&c_trackerOH_1),.io_probedack(d_trackerOH[1]&_GEN_1&d_drop),.io_probesack(_c_first_T&c_trackerOH_1&_clearOH_T_1&_GEN_3),.io_d_last(d_trackerOH[1]&_GEN&d_response&d_last),.io_e_last(auto_in_e_bits_sink==2'h1&auto_in_e_valid),.io_source(_TLBroadcastTracker_1_io_source),.io_line(_TLBroadcastTracker_1_io_line),.io_idle(_TLBroadcastTracker_1_io_idle),.io_need_d(_TLBroadcastTracker_1_io_need_d)); 
  TLBroadcastTracker_2 TLBroadcastTracker_2(.clock(clock),.reset(reset),.io_in_a_first(~(|a_first_counter)),.io_in_a_ready(_TLBroadcastTracker_2_io_in_a_ready),.io_in_a_valid(auto_in_a_valid&filter_io_request_bits_mshr_lo[2]&_GEN_8),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_data(auto_in_a_bits_data),.io_out_a_ready(auto_out_a_ready&(idle_1 ? ~_GEN_6:state_1_3)),.io_out_a_valid(_TLBroadcastTracker_2_io_out_a_valid),.io_out_a_bits_opcode(_TLBroadcastTracker_2_io_out_a_bits_opcode),.io_out_a_bits_param(_TLBroadcastTracker_2_io_out_a_bits_param),.io_out_a_bits_size(_TLBroadcastTracker_2_io_out_a_bits_size),.io_out_a_bits_source(_TLBroadcastTracker_2_io_out_a_bits_source),.io_out_a_bits_address(_TLBroadcastTracker_2_io_out_a_bits_address),.io_out_a_bits_mask(_TLBroadcastTracker_2_io_out_a_bits_mask),.io_out_a_bits_data(_TLBroadcastTracker_2_io_out_a_bits_data),.io_probe_valid(_sack_T&_filter_io_response_bits_mshr==2'h2),.io_probe_bits_count(~_filter_io_response_bits_allocOH),.io_probenack(_GEN_2&c_trackerOH_2),.io_probedack(d_trackerOH[2]&_GEN_1&d_drop),.io_probesack(_c_first_T&c_trackerOH_2&_clearOH_T_1&_GEN_3),.io_d_last(d_trackerOH[2]&_GEN&d_response&d_last),.io_e_last(auto_in_e_bits_sink==2'h2&auto_in_e_valid),.io_source(_TLBroadcastTracker_2_io_source),.io_line(_TLBroadcastTracker_2_io_line),.io_idle(_TLBroadcastTracker_2_io_idle),.io_need_d(_TLBroadcastTracker_2_io_need_d)); 
  TLBroadcastTracker_3 TLBroadcastTracker_3(.clock(clock),.reset(reset),.io_in_a_first(~(|a_first_counter)),.io_in_a_ready(_TLBroadcastTracker_3_io_in_a_ready),.io_in_a_valid(auto_in_a_valid&filter_io_request_bits_mshr_lo[3]&_GEN_8),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_data(auto_in_a_bits_data),.io_out_a_ready(auto_out_a_ready&(idle_1 ? ~_GEN_5:state_1_4)),.io_out_a_valid(_TLBroadcastTracker_3_io_out_a_valid),.io_out_a_bits_opcode(_TLBroadcastTracker_3_io_out_a_bits_opcode),.io_out_a_bits_param(_TLBroadcastTracker_3_io_out_a_bits_param),.io_out_a_bits_size(_TLBroadcastTracker_3_io_out_a_bits_size),.io_out_a_bits_source(_TLBroadcastTracker_3_io_out_a_bits_source),.io_out_a_bits_address(_TLBroadcastTracker_3_io_out_a_bits_address),.io_out_a_bits_mask(_TLBroadcastTracker_3_io_out_a_bits_mask),.io_out_a_bits_data(_TLBroadcastTracker_3_io_out_a_bits_data),.io_probe_valid(_sack_T&(&_filter_io_response_bits_mshr)),.io_probe_bits_count(~_filter_io_response_bits_allocOH),.io_probenack(_GEN_2&c_trackerOH_3),.io_probedack(d_trackerOH[3]&_GEN_1&d_drop),.io_probesack(_c_first_T&c_trackerOH_3&_clearOH_T_1&_GEN_3),.io_d_last(d_trackerOH[3]&_GEN&d_response&d_last),.io_e_last((&auto_in_e_bits_sink)&auto_in_e_valid),.io_source(_TLBroadcastTracker_3_io_source),.io_line(_TLBroadcastTracker_3_io_line),.io_idle(_TLBroadcastTracker_3_io_idle),.io_need_d(_TLBroadcastTracker_3_io_need_d)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_b_valid=probe_todo; 
  assign auto_in_b_bits_param=probe_perms; 
  assign auto_in_b_bits_address=nodeIn_b_bits_b_address; 
  assign auto_in_c_ready=nodeIn_c_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_bits_T_23; 
  assign auto_in_d_bits_param=_nodeIn_d_bits_T_20; 
  assign auto_in_d_bits_size=_nodeIn_d_bits_T_17; 
  assign auto_in_d_bits_source=_nodeIn_d_bits_T_14; 
  assign auto_in_d_bits_sink=_nodeIn_d_bits_T_11; 
  assign auto_in_d_bits_denied=_nodeIn_d_bits_T_8; 
  assign auto_in_d_bits_data=muxState_1 ? auto_out_d_bits_data:64'h0; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_bits_T_2; 
  assign auto_out_a_valid=nodeOut_a_valid; 
  assign auto_out_a_bits_opcode=(muxState_1_1 ? _TLBroadcastTracker_io_out_a_bits_opcode:3'h0)|(muxState_1_2 ? _TLBroadcastTracker_1_io_out_a_bits_opcode:3'h0)|(muxState_1_3 ? _TLBroadcastTracker_2_io_out_a_bits_opcode:3'h0)|(muxState_1_4 ? _TLBroadcastTracker_3_io_out_a_bits_opcode:3'h0); 
  assign auto_out_a_bits_param=(muxState_1_1 ? _TLBroadcastTracker_io_out_a_bits_param:3'h0)|(muxState_1_2 ? _TLBroadcastTracker_1_io_out_a_bits_param:3'h0)|(muxState_1_3 ? _TLBroadcastTracker_2_io_out_a_bits_param:3'h0)|(muxState_1_4 ? _TLBroadcastTracker_3_io_out_a_bits_param:3'h0); 
  assign auto_out_a_bits_size=(muxState_1_0 ? auto_in_c_bits_size:3'h0)|(muxState_1_1 ? _TLBroadcastTracker_io_out_a_bits_size:3'h0)|(muxState_1_2 ? _TLBroadcastTracker_1_io_out_a_bits_size:3'h0)|(muxState_1_3 ? _TLBroadcastTracker_2_io_out_a_bits_size:3'h0)|(muxState_1_4 ? _TLBroadcastTracker_3_io_out_a_bits_size:3'h0); 
  assign auto_out_a_bits_source=(muxState_1_0 ? {(&auto_in_c_bits_opcode) ? 2'h2:2'h1,(&auto_in_c_bits_opcode) ? auto_in_c_bits_source:(c_trackerOH_0 ? _TLBroadcastTracker_io_source:5'h0)|(c_trackerOH_1 ? _TLBroadcastTracker_1_io_source:5'h0)|(c_trackerOH_2 ? _TLBroadcastTracker_2_io_source:5'h0)|(c_trackerOH_3 ? _TLBroadcastTracker_3_io_source:5'h0)}:7'h0)|(muxState_1_1 ? _TLBroadcastTracker_io_out_a_bits_source:7'h0)|(muxState_1_2 ? _TLBroadcastTracker_1_io_out_a_bits_source:7'h0)|(muxState_1_3 ? _TLBroadcastTracker_2_io_out_a_bits_source:7'h0)|(muxState_1_4 ? _TLBroadcastTracker_3_io_out_a_bits_source:7'h0); 
  assign auto_out_a_bits_address=(muxState_1_0 ? auto_in_c_bits_address:32'h0)|(muxState_1_1 ? _TLBroadcastTracker_io_out_a_bits_address:32'h0)|(muxState_1_2 ? _TLBroadcastTracker_1_io_out_a_bits_address:32'h0)|(muxState_1_3 ? _TLBroadcastTracker_2_io_out_a_bits_address:32'h0)|(muxState_1_4 ? _TLBroadcastTracker_3_io_out_a_bits_address:32'h0); 
  assign auto_out_a_bits_mask=(muxState_1_0 ? {putfull_bits_a_mask_acc_5|putfull_bits_a_mask_eq_5&auto_in_c_bits_address[0],putfull_bits_a_mask_acc_5|putfull_bits_a_mask_eq_5&~(auto_in_c_bits_address[0]),putfull_bits_a_mask_acc_4|putfull_bits_a_mask_eq_4&auto_in_c_bits_address[0],putfull_bits_a_mask_acc_4|putfull_bits_a_mask_eq_4&~(auto_in_c_bits_address[0]),putfull_bits_a_mask_acc_3|putfull_bits_a_mask_eq_3&auto_in_c_bits_address[0],putfull_bits_a_mask_acc_3|putfull_bits_a_mask_eq_3&~(auto_in_c_bits_address[0]),putfull_bits_a_mask_acc_2|putfull_bits_a_mask_eq_2&auto_in_c_bits_address[0],putfull_bits_a_mask_acc_2|putfull_bits_a_mask_eq_2&~(auto_in_c_bits_address[0])}:8'h0)|(muxState_1_1 ? _TLBroadcastTracker_io_out_a_bits_mask:8'h0)|(muxState_1_2 ? _TLBroadcastTracker_1_io_out_a_bits_mask:8'h0)|(muxState_1_3 ? _TLBroadcastTracker_2_io_out_a_bits_mask:8'h0)|(muxState_1_4 ? _TLBroadcastTracker_3_io_out_a_bits_mask:8'h0); 
  assign auto_out_a_bits_data=(muxState_1_0 ? auto_in_c_bits_data:64'h0)|(muxState_1_1 ? _TLBroadcastTracker_io_out_a_bits_data:64'h0)|(muxState_1_2 ? _TLBroadcastTracker_1_io_out_a_bits_data:64'h0)|(muxState_1_3 ? _TLBroadcastTracker_2_io_out_a_bits_data:64'h0)|(muxState_1_4 ? _TLBroadcastTracker_3_io_out_a_bits_data:64'h0); 
  assign auto_out_d_ready=nodeOut_d_ready; 
endmodule
 
module TLMonitor_22 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [2:0] io_in_a_bits_size,
  input [6:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [2:0] io_in_d_bits_size,
  input [6:0] io_in_d_bits_source,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [12:0] _GEN={10'h0,io_in_a_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [2:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [2:0] size ;  
   reg [6:0] source ;  
   reg [31:0] address ;  
   reg [2:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [2:0] size_1 ;  
   reg [6:0] source_1 ;  
   reg denied ;  
   reg [127:0] inflight ;  
   reg [511:0] inflight_opcodes ;  
   reg [511:0] inflight_sizes ;  
   reg [2:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==3'h0 ;  
   reg [2:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==3'h0 ;  
   wire [511:0] _GEN_0={503'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN_0 ;  
   wire [127:0] _GEN_1={121'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [127:0] _GEN_3={121'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [127:0] inflight_1 ;  
   reg [511:0] inflight_sizes_1 ;  
   reg [2:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==3'h0 ;  
   reg [31:0] watchdog_1 ;  
   wire [12:0] _is_aligned_mask_T_1=13'h3F<<_GEN ;  
   wire [5:0] _GEN_4=io_in_a_bits_address[5:0]&~(_is_aligned_mask_T_1[5:0]) ;  
   wire _mask_T=io_in_a_bits_size>3'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_a_bits_param>3'h2 ;  
   wire _GEN_7=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_8=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_9=io_in_a_bits_size!=3'h7&io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_11=io_in_a_bits_mask!=mask ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_18=io_in_d_bits_size<3'h3 ;  
   wire _GEN_19=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_20=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_21=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_22=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_23=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [127:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 128'h1<<_GEN_1:128'h0 ;  
   wire _GEN_24=io_in_d_valid&d_first_1 ;  
   wire _GEN_25=_GEN_24&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_26=_GEN_25&same_cycle_resp&~reset ;  
   wire _GEN_27=_GEN_25&~same_cycle_resp&~reset ;  
   wire _GEN_28=io_in_d_valid&d_first_2&d_release_ack&~reset ;  
   wire [127:0] _GEN_29=inflight>>_GEN_1 ;  
   wire [127:0] _GEN_30=inflight>>_GEN_3 ;  
   wire [511:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_0 ;  
   wire [127:0] _GEN_31=inflight_1>>_GEN_3 ;  
   wire [511:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_0 ;  
  always @( posedge clock)
       begin 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_4))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_29[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~reset&~(_GEN_30[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_d_bits_size!=_a_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_25 ? 128'h1<<_GEN_3:128'h0)|a_set_wo_ready==128'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==128'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(_GEN_31[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&io_in_d_bits_size!=_c_size_lookup_T_1[3:1])
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==128'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/subsystem/BankedL2Params.scala:65:103)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [12:0] _a_first_beats1_decode_T_1=13'h3F<<_GEN ;  
   wire [12:0] _a_first_beats1_decode_T_5=13'h3F<<_GEN ;  
   wire [12:0] _GEN_32={10'h0,io_in_d_bits_size} ;  
   wire [12:0] _d_first_beats1_decode_T_1=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_5=13'h3F<<_GEN_32 ;  
   wire [12:0] _d_first_beats1_decode_T_9=13'h3F<<_GEN_32 ;  
   wire [1026:0] _GEN_33={1018'h0,io_in_a_bits_source,2'h0} ;  
   wire [1038:0] _GEN_34={1030'h0,io_in_d_bits_source,2'h0} ;  
   wire [1038:0] _d_opcodes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_opcodes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_5=1039'hF<<_GEN_34 ;  
   wire [1026:0] _a_sizes_set_T_1={1023'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:4'h0}<<_GEN_33 ;  
   wire [1038:0] _d_sizes_clr_T_11=1039'hF<<_GEN_34 ;  
   wire _d_first_T_2=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_35=_d_first_T_2&d_first_1&~d_release_ack ;  
   wire _GEN_36=_d_first_T_2&d_first_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=3'h0;
              d_first_counter <=3'h0;
              inflight <=128'h0;
              inflight_opcodes <=512'h0;
              inflight_sizes <=512'h0;
              a_first_counter_1 <=3'h0;
              d_first_counter_1 <=3'h0;
              watchdog <=32'h0;
              inflight_1 <=128'h0;
              inflight_sizes_1 <=512'h0;
              d_first_counter_2 <=3'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-3'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_1[5:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 3'h0:~(_a_first_beats1_decode_T_5[5:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-3'h1;
                 end 
              if (_d_first_T_2)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-3'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[5:3]):3'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[5:3]):3'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-3'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[5:3]):3'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-3'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|(_GEN_2 ? 128'h1<<_GEN_1:128'h0))&~(_GEN_35 ? 128'h1<<_GEN_3:128'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_opcodes_clr_T_5[511:0]:512'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[511:0]:512'h0))&~(_GEN_35 ? _d_sizes_clr_T_5[511:0]:512'h0);
              if (_a_first_T_1|_d_first_T_2)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_36 ? 128'h1<<_GEN_3:128'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_36 ? _d_sizes_clr_T_11[511:0]:512'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_2&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module BankBinder (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [2:0] auto_in_a_bits_size,
  input [6:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [2:0] auto_in_d_bits_size,
  output [6:0] auto_in_d_bits_source,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [2:0] auto_out_a_bits_size,
  output [6:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [2:0] auto_out_d_bits_size,
  input [6:0] auto_out_d_bits_source,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt) ; 
  TLMonitor_22 monitor(.clock(clock),.reset(reset),.io_in_a_ready(auto_out_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_out_d_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source),.io_in_d_bits_denied(auto_out_d_bits_denied),.io_in_d_bits_corrupt(auto_out_d_bits_corrupt)); 
  assign auto_in_a_ready=auto_out_a_ready; 
  assign auto_in_d_valid=auto_out_d_valid; 
  assign auto_in_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_d_bits_source=auto_out_d_bits_source; 
  assign auto_in_d_bits_denied=auto_out_d_bits_denied; 
  assign auto_in_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign auto_out_a_valid=auto_in_a_valid; 
  assign auto_out_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_a_bits_param=auto_in_a_bits_param; 
  assign auto_out_a_bits_size=auto_in_a_bits_size; 
  assign auto_out_a_bits_source=auto_in_a_bits_source; 
  assign auto_out_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_a_bits_mask=auto_in_a_bits_mask; 
  assign auto_out_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_d_ready=auto_in_d_ready; 
endmodule
 
module CoherenceManagerWrapper (
  input auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready,
  output auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid,
  output [2:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode,
  output [2:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_param,
  output [2:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size,
  output [6:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source,
  output [31:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address,
  output [7:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask,
  output [63:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data,
  output auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready,
  input auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid,
  input [2:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode,
  input [2:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size,
  input [6:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source,
  input auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied,
  input [63:0] auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data,
  input auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt,
  output auto_coherent_jbar_in_a_ready,
  input auto_coherent_jbar_in_a_valid,
  input [2:0] auto_coherent_jbar_in_a_bits_opcode,
  input [2:0] auto_coherent_jbar_in_a_bits_param,
  input [2:0] auto_coherent_jbar_in_a_bits_size,
  input [4:0] auto_coherent_jbar_in_a_bits_source,
  input [31:0] auto_coherent_jbar_in_a_bits_address,
  input [7:0] auto_coherent_jbar_in_a_bits_mask,
  input [63:0] auto_coherent_jbar_in_a_bits_data,
  input auto_coherent_jbar_in_a_bits_corrupt,
  input auto_coherent_jbar_in_b_ready,
  output auto_coherent_jbar_in_b_valid,
  output [1:0] auto_coherent_jbar_in_b_bits_param,
  output [31:0] auto_coherent_jbar_in_b_bits_address,
  output auto_coherent_jbar_in_c_ready,
  input auto_coherent_jbar_in_c_valid,
  input [2:0] auto_coherent_jbar_in_c_bits_opcode,
  input [2:0] auto_coherent_jbar_in_c_bits_param,
  input [2:0] auto_coherent_jbar_in_c_bits_size,
  input [4:0] auto_coherent_jbar_in_c_bits_source,
  input [31:0] auto_coherent_jbar_in_c_bits_address,
  input [63:0] auto_coherent_jbar_in_c_bits_data,
  input auto_coherent_jbar_in_c_bits_corrupt,
  input auto_coherent_jbar_in_d_ready,
  output auto_coherent_jbar_in_d_valid,
  output [2:0] auto_coherent_jbar_in_d_bits_opcode,
  output [1:0] auto_coherent_jbar_in_d_bits_param,
  output [2:0] auto_coherent_jbar_in_d_bits_size,
  output [4:0] auto_coherent_jbar_in_d_bits_source,
  output [1:0] auto_coherent_jbar_in_d_bits_sink,
  output auto_coherent_jbar_in_d_bits_denied,
  output [63:0] auto_coherent_jbar_in_d_bits_data,
  output auto_coherent_jbar_in_d_bits_corrupt,
  input auto_coherent_jbar_in_e_valid,
  input [1:0] auto_coherent_jbar_in_e_bits_sink,
  input auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock,
  input auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset,
  input auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock,
  input auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset,
  output auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock,
  output auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset) ; 
   wire _binder_auto_in_a_ready ;  
   wire _binder_auto_in_d_valid ;  
   wire [2:0] _binder_auto_in_d_bits_opcode ;  
   wire [2:0] _binder_auto_in_d_bits_size ;  
   wire [6:0] _binder_auto_in_d_bits_source ;  
   wire _binder_auto_in_d_bits_denied ;  
   wire [63:0] _binder_auto_in_d_bits_data ;  
   wire _binder_auto_in_d_bits_corrupt ;  
   wire _broadcast_1_auto_out_a_valid ;  
   wire [2:0] _broadcast_1_auto_out_a_bits_opcode ;  
   wire [2:0] _broadcast_1_auto_out_a_bits_param ;  
   wire [2:0] _broadcast_1_auto_out_a_bits_size ;  
   wire [6:0] _broadcast_1_auto_out_a_bits_source ;  
   wire [31:0] _broadcast_1_auto_out_a_bits_address ;  
   wire [7:0] _broadcast_1_auto_out_a_bits_mask ;  
   wire [63:0] _broadcast_1_auto_out_a_bits_data ;  
   wire _broadcast_1_auto_out_d_ready ;  
  TLBroadcast broadcast_1(.clock(auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock),.reset(auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset),.auto_in_a_ready(auto_coherent_jbar_in_a_ready),.auto_in_a_valid(auto_coherent_jbar_in_a_valid),.auto_in_a_bits_opcode(auto_coherent_jbar_in_a_bits_opcode),.auto_in_a_bits_param(auto_coherent_jbar_in_a_bits_param),.auto_in_a_bits_size(auto_coherent_jbar_in_a_bits_size),.auto_in_a_bits_source(auto_coherent_jbar_in_a_bits_source),.auto_in_a_bits_address(auto_coherent_jbar_in_a_bits_address),.auto_in_a_bits_mask(auto_coherent_jbar_in_a_bits_mask),.auto_in_a_bits_data(auto_coherent_jbar_in_a_bits_data),.auto_in_a_bits_corrupt(auto_coherent_jbar_in_a_bits_corrupt),.auto_in_b_ready(auto_coherent_jbar_in_b_ready),.auto_in_b_valid(auto_coherent_jbar_in_b_valid),.auto_in_b_bits_param(auto_coherent_jbar_in_b_bits_param),.auto_in_b_bits_address(auto_coherent_jbar_in_b_bits_address),.auto_in_c_ready(auto_coherent_jbar_in_c_ready),.auto_in_c_valid(auto_coherent_jbar_in_c_valid),.auto_in_c_bits_opcode(auto_coherent_jbar_in_c_bits_opcode),.auto_in_c_bits_param(auto_coherent_jbar_in_c_bits_param),.auto_in_c_bits_size(auto_coherent_jbar_in_c_bits_size),.auto_in_c_bits_source(auto_coherent_jbar_in_c_bits_source),.auto_in_c_bits_address(auto_coherent_jbar_in_c_bits_address),.auto_in_c_bits_data(auto_coherent_jbar_in_c_bits_data),.auto_in_c_bits_corrupt(auto_coherent_jbar_in_c_bits_corrupt),.auto_in_d_ready(auto_coherent_jbar_in_d_ready),.auto_in_d_valid(auto_coherent_jbar_in_d_valid),.auto_in_d_bits_opcode(auto_coherent_jbar_in_d_bits_opcode),.auto_in_d_bits_param(auto_coherent_jbar_in_d_bits_param),.auto_in_d_bits_size(auto_coherent_jbar_in_d_bits_size),.auto_in_d_bits_source(auto_coherent_jbar_in_d_bits_source),.auto_in_d_bits_sink(auto_coherent_jbar_in_d_bits_sink),.auto_in_d_bits_denied(auto_coherent_jbar_in_d_bits_denied),.auto_in_d_bits_data(auto_coherent_jbar_in_d_bits_data),.auto_in_d_bits_corrupt(auto_coherent_jbar_in_d_bits_corrupt),.auto_in_e_valid(auto_coherent_jbar_in_e_valid),.auto_in_e_bits_sink(auto_coherent_jbar_in_e_bits_sink),.auto_out_a_ready(_binder_auto_in_a_ready),.auto_out_a_valid(_broadcast_1_auto_out_a_valid),.auto_out_a_bits_opcode(_broadcast_1_auto_out_a_bits_opcode),.auto_out_a_bits_param(_broadcast_1_auto_out_a_bits_param),.auto_out_a_bits_size(_broadcast_1_auto_out_a_bits_size),.auto_out_a_bits_source(_broadcast_1_auto_out_a_bits_source),.auto_out_a_bits_address(_broadcast_1_auto_out_a_bits_address),.auto_out_a_bits_mask(_broadcast_1_auto_out_a_bits_mask),.auto_out_a_bits_data(_broadcast_1_auto_out_a_bits_data),.auto_out_d_ready(_broadcast_1_auto_out_d_ready),.auto_out_d_valid(_binder_auto_in_d_valid),.auto_out_d_bits_opcode(_binder_auto_in_d_bits_opcode),.auto_out_d_bits_size(_binder_auto_in_d_bits_size),.auto_out_d_bits_source(_binder_auto_in_d_bits_source),.auto_out_d_bits_denied(_binder_auto_in_d_bits_denied),.auto_out_d_bits_data(_binder_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_binder_auto_in_d_bits_corrupt)); 
  BankBinder binder(.clock(auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock),.reset(auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset),.auto_in_a_ready(_binder_auto_in_a_ready),.auto_in_a_valid(_broadcast_1_auto_out_a_valid),.auto_in_a_bits_opcode(_broadcast_1_auto_out_a_bits_opcode),.auto_in_a_bits_param(_broadcast_1_auto_out_a_bits_param),.auto_in_a_bits_size(_broadcast_1_auto_out_a_bits_size),.auto_in_a_bits_source(_broadcast_1_auto_out_a_bits_source),.auto_in_a_bits_address(_broadcast_1_auto_out_a_bits_address),.auto_in_a_bits_mask(_broadcast_1_auto_out_a_bits_mask),.auto_in_a_bits_data(_broadcast_1_auto_out_a_bits_data),.auto_in_d_ready(_broadcast_1_auto_out_d_ready),.auto_in_d_valid(_binder_auto_in_d_valid),.auto_in_d_bits_opcode(_binder_auto_in_d_bits_opcode),.auto_in_d_bits_size(_binder_auto_in_d_bits_size),.auto_in_d_bits_source(_binder_auto_in_d_bits_source),.auto_in_d_bits_denied(_binder_auto_in_d_bits_denied),.auto_in_d_bits_data(_binder_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_binder_auto_in_d_bits_corrupt),.auto_out_a_ready(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready),.auto_out_a_valid(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid),.auto_out_a_bits_opcode(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode),.auto_out_a_bits_param(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_param),.auto_out_a_bits_size(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size),.auto_out_a_bits_source(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source),.auto_out_a_bits_address(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address),.auto_out_a_bits_mask(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask),.auto_out_a_bits_data(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data),.auto_out_d_ready(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready),.auto_out_d_valid(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid),.auto_out_d_bits_opcode(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode),.auto_out_d_bits_size(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size),.auto_out_d_bits_source(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source),.auto_out_d_bits_denied(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied),.auto_out_d_bits_data(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data),.auto_out_d_bits_corrupt(auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt)); 
  assign auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock=auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock; 
  assign auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset=auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset; 
endmodule
 
module TLMonitor_23 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_b_ready,
  input io_in_b_valid,
  input [2:0] io_in_b_bits_opcode,
  input [1:0] io_in_b_bits_param,
  input [3:0] io_in_b_bits_size,
  input io_in_b_bits_source,
  input [31:0] io_in_b_bits_address,
  input [7:0] io_in_b_bits_mask,
  input io_in_b_bits_corrupt,
  input io_in_c_ready,
  input io_in_c_valid,
  input [2:0] io_in_c_bits_opcode,
  input [2:0] io_in_c_bits_param,
  input [3:0] io_in_c_bits_size,
  input io_in_c_bits_source,
  input [31:0] io_in_c_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt,
  input io_in_e_ready,
  input io_in_e_valid,
  input [1:0] io_in_e_bits_sink) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire [26:0] _GEN_0={23'h0,io_in_c_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg source ;  
   reg [31:0] address ;  
   wire _d_first_T_3=io_in_d_ready&io_in_d_valid ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [8:0] b_first_counter ;  
   reg [2:0] opcode_2 ;  
   reg [1:0] param_2 ;  
   reg [3:0] size_2 ;  
   reg source_2 ;  
   reg [31:0] address_1 ;  
   wire _c_first_T_1=io_in_c_ready&io_in_c_valid ;  
   reg [8:0] c_first_counter ;  
   reg [2:0] opcode_3 ;  
   reg [2:0] param_3 ;  
   reg [3:0] size_3 ;  
   reg source_3 ;  
   reg [31:0] address_2 ;  
   reg [1:0] inflight ;  
   reg [7:0] inflight_opcodes ;  
   reg [15:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [7:0] _a_opcode_lookup_T_1=inflight_opcodes>>{5'h0,io_in_d_bits_source,2'h0} ;  
   wire [1:0] _GEN_1={1'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [1:0] _GEN_3={1'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [1:0] inflight_1 ;  
   reg [15:0] inflight_sizes_1 ;  
   reg [8:0] c_first_counter_1 ;  
   wire c_first_1=c_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   wire _GEN_4=io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1] ;  
   wire [1:0] _GEN_5={1'h0,io_in_c_bits_source} ;  
   wire _GEN_6=_c_first_T_1&c_first_1&_GEN_4 ;  
   reg [31:0] watchdog_1 ;  
   reg [3:0] inflight_2 ;  
   reg [8:0] d_first_counter_3 ;  
   wire d_first_3=d_first_counter_3==9'h0 ;  
   wire _GEN_7=_d_first_T_3&d_first_3&io_in_d_bits_opcode[2]&~(io_in_d_bits_opcode[1]) ;  
   wire [3:0] _GEN_8={2'h0,io_in_d_bits_sink} ;  
   wire [3:0] d_set=_GEN_7 ? 4'h1<<_GEN_8:4'h0 ;  
   wire _GEN_9=io_in_e_ready&io_in_e_valid ;  
   wire [3:0] _GEN_10={2'h0,io_in_e_bits_sink} ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_11=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_12=io_in_a_bits_size<4'hD ;  
   wire _GEN_13=io_in_a_bits_size<4'h7 ;  
   wire _GEN_14=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_15=_GEN_12&_GEN_13&_GEN_14 ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_17=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_18={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_19={io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0 ;  
   wire _GEN_20={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_21={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_22={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_23=_GEN_17|_GEN_18 ;  
   wire _GEN_24=~io_in_a_bits_source&io_in_a_bits_size==4'h6&_GEN_12&(_GEN_23|_GEN_19|_GEN_20|_GEN_21|_GEN_22|_GEN_14) ;  
   wire _GEN_25=io_in_a_bits_param>3'h2 ;  
   wire _GEN_26=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_27=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_28=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_29=_GEN_12&_GEN_18 ;  
   wire _GEN_30=io_in_a_bits_mask!=mask ;  
   wire _GEN_31=_GEN_12&(_GEN_29|_GEN_13&(_GEN_17|_GEN_20|_GEN_21|_GEN_14)|io_in_a_bits_size<4'h9&_GEN_22) ;  
   wire _GEN_32=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_33=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_34=_GEN_12&io_in_a_bits_size<4'h4&(_GEN_23|_GEN_20|_GEN_21) ;  
   wire _GEN_35=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_36=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_37=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_38=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_39=io_in_d_bits_size<4'h3 ;  
   wire _GEN_40=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_41=io_in_d_bits_param==2'h2 ;  
   wire _GEN_42=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_43=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_44=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_45=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_46=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire [19:0] _GEN_47={io_in_b_bits_address[31:14],~(io_in_b_bits_address[13:12])} ;  
   wire [5:0] _GEN_48={io_in_b_bits_address[31:28],~(io_in_b_bits_address[27:26])} ;  
   wire [15:0] _GEN_49={io_in_b_bits_address[31:26],io_in_b_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_50={io_in_b_bits_address[31:17],~(io_in_b_bits_address[16])} ;  
   wire _GEN_51=io_in_b_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_52={io_in_b_bits_address[31],~(io_in_b_bits_address[30:29])} ;  
   wire address_ok=~(|_GEN_47)|~(|_GEN_48)|~(|_GEN_49)|~(|(io_in_b_bits_address[31:12]))|~(|_GEN_50)|~_GEN_51|~(|_GEN_52) ;  
   wire [26:0] _is_aligned_mask_T_4=27'hFFF<<io_in_b_bits_size ;  
   wire [11:0] _GEN_53=io_in_b_bits_address[11:0]&~(_is_aligned_mask_T_4[11:0]) ;  
   wire _mask_T_1=io_in_b_bits_size>4'h2 ;  
   wire mask_size_3=io_in_b_bits_size[1:0]==2'h2 ;  
   wire mask_acc_14=_mask_T_1|mask_size_3&~(io_in_b_bits_address[2]) ;  
   wire mask_acc_15=_mask_T_1|mask_size_3&io_in_b_bits_address[2] ;  
   wire mask_size_4=io_in_b_bits_size[1:0]==2'h1 ;  
   wire mask_eq_16=~(io_in_b_bits_address[2])&~(io_in_b_bits_address[1]) ;  
   wire mask_acc_16=mask_acc_14|mask_size_4&mask_eq_16 ;  
   wire mask_eq_17=~(io_in_b_bits_address[2])&io_in_b_bits_address[1] ;  
   wire mask_acc_17=mask_acc_14|mask_size_4&mask_eq_17 ;  
   wire mask_eq_18=io_in_b_bits_address[2]&~(io_in_b_bits_address[1]) ;  
   wire mask_acc_18=mask_acc_15|mask_size_4&mask_eq_18 ;  
   wire mask_eq_19=io_in_b_bits_address[2]&io_in_b_bits_address[1] ;  
   wire mask_acc_19=mask_acc_15|mask_size_4&mask_eq_19 ;  
   wire [7:0] mask_1={mask_acc_19|mask_eq_19&io_in_b_bits_address[0],mask_acc_19|mask_eq_19&~(io_in_b_bits_address[0]),mask_acc_18|mask_eq_18&io_in_b_bits_address[0],mask_acc_18|mask_eq_18&~(io_in_b_bits_address[0]),mask_acc_17|mask_eq_17&io_in_b_bits_address[0],mask_acc_17|mask_eq_17&~(io_in_b_bits_address[0]),mask_acc_16|mask_eq_16&io_in_b_bits_address[0],mask_acc_16|mask_eq_16&~(io_in_b_bits_address[0])} ;  
   wire _GEN_54=io_in_b_valid&io_in_b_bits_opcode==3'h6&~reset ;  
   wire _GEN_55=io_in_b_bits_mask!=mask_1 ;  
   wire _GEN_56=io_in_b_valid&io_in_b_bits_opcode==3'h4&~reset ;  
   wire _GEN_57=io_in_b_valid&io_in_b_bits_opcode==3'h0&~reset ;  
   wire _GEN_58=io_in_b_valid&io_in_b_bits_opcode==3'h1&~reset ;  
   wire _GEN_59=io_in_b_valid&io_in_b_bits_opcode==3'h2&~reset ;  
   wire _GEN_60=io_in_b_valid&io_in_b_bits_opcode==3'h3&~reset ;  
   wire _GEN_61=io_in_b_valid&io_in_b_bits_opcode==3'h5&~reset ;  
   wire [26:0] _is_aligned_mask_T_7=27'hFFF<<_GEN_0 ;  
   wire [11:0] _GEN_62=io_in_c_bits_address[11:0]&~(_is_aligned_mask_T_7[11:0]) ;  
   wire [19:0] _GEN_63={io_in_c_bits_address[31:14],~(io_in_c_bits_address[13:12])} ;  
   wire [5:0] _GEN_64={io_in_c_bits_address[31:28],~(io_in_c_bits_address[27:26])} ;  
   wire [15:0] _GEN_65={io_in_c_bits_address[31:26],io_in_c_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_66={io_in_c_bits_address[31:17],~(io_in_c_bits_address[16])} ;  
   wire _GEN_67=io_in_c_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_68={io_in_c_bits_address[31],~(io_in_c_bits_address[30:29])} ;  
   wire address_ok_1=~(|_GEN_63)|~(|_GEN_64)|~(|_GEN_65)|~(|(io_in_c_bits_address[31:12]))|~(|_GEN_66)|~_GEN_67|~(|_GEN_68) ;  
   wire _GEN_69=io_in_c_valid&io_in_c_bits_opcode==3'h4&~reset ;  
   wire _GEN_70=io_in_c_bits_size<4'h3 ;  
   wire _GEN_71=io_in_c_valid&io_in_c_bits_opcode==3'h5&~reset ;  
   wire _GEN_72=io_in_c_bits_size<4'hD ;  
   wire _GEN_73=_GEN_72&io_in_c_bits_size<4'h7&~_GEN_67 ;  
   wire _GEN_74=io_in_c_valid&io_in_c_bits_opcode==3'h6&~reset ;  
   wire _GEN_75=~io_in_c_bits_source&io_in_c_bits_size==4'h6&_GEN_72&(~(|(io_in_c_bits_address[31:12]))|~(|_GEN_63)|~(|_GEN_66)|~(|_GEN_65)|~(|_GEN_64)|~(|_GEN_68)|~_GEN_67) ;  
   wire _GEN_76=io_in_c_valid&(&io_in_c_bits_opcode)&~reset ;  
   wire _GEN_77=io_in_c_valid&io_in_c_bits_opcode==3'h0&~reset ;  
   wire _GEN_78=io_in_c_valid&io_in_c_bits_opcode==3'h1&~reset ;  
   wire _GEN_79=io_in_c_valid&io_in_c_bits_opcode==3'h2&~reset ;  
   wire _GEN_80=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_81=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_82=io_in_b_valid&(|b_first_counter)&~reset ;  
   wire _GEN_83=io_in_c_valid&(|c_first_counter)&~reset ;  
   wire [15:0] _GEN_84={12'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [1:0] a_set_wo_ready=_same_cycle_resp_T_1 ? 2'h1<<_GEN_1:2'h0 ;  
   wire _GEN_85=io_in_d_valid&d_first_1 ;  
   wire _GEN_86=_GEN_85&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_87=_GEN_86&same_cycle_resp&~reset ;  
   wire _GEN_88=_GEN_86&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_89={4'h0,io_in_d_bits_size} ;  
   wire _same_cycle_resp_T_3=io_in_c_valid&c_first_1 ;  
   wire [1:0] c_set_wo_ready=_same_cycle_resp_T_3&_GEN_4 ? 2'h1<<_GEN_5:2'h0 ;  
   wire _GEN_90=io_in_d_valid&d_first_2 ;  
   wire _GEN_91=_GEN_90&d_release_ack ;  
   wire same_cycle_resp_1=_same_cycle_resp_T_3&io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1]&io_in_c_bits_source==io_in_d_bits_source ;  
   wire [1:0] _GEN_92=inflight>>_GEN_1 ;  
   wire [1:0] _GEN_93=inflight>>_GEN_3 ;  
   wire [15:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_84 ;  
   wire [1:0] _GEN_94=inflight_1>>_GEN_5 ;  
   wire [1:0] _GEN_95=inflight_1>>_GEN_3 ;  
   wire [15:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_84 ;  
   wire [3:0] _GEN_96=inflight_2>>_GEN_8 ;  
   wire [3:0] _GEN_97=(d_set|inflight_2)>>_GEN_10 ;  
  always @( posedge clock)
       begin 
         if (_GEN_16&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_GEN_24)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(_GEN_29|_GEN_13&(_GEN_17|_GEN_19|_GEN_20|_GEN_21|_GEN_22|_GEN_14)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&~_GEN_34)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_35&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~_GEN_34)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~(_GEN_12&_GEN_29))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&_GEN_30)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_40&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_39)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&_GEN_41)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_42&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_44&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&~_GEN_43)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_b_valid&~reset&(&io_in_b_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'B' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_54&~(~io_in_b_bits_source&io_in_b_bits_size==4'h6&io_in_b_bits_size<4'hD&(~(|(io_in_b_bits_address[31:12]))|~(|_GEN_47)|~(|_GEN_50)|~(|_GEN_49)|~(|_GEN_48)|~(|_GEN_52)|~_GEN_51)))
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_54&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_54&(|_GEN_53))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_54&(&io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_54&_GEN_55)
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_54&io_in_b_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_56&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Get carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_56&(|_GEN_53))
            begin 
              if (1)$display("Assertion failed: 'B' channel Get address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_56&(|io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel Get carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_56&_GEN_55)
            begin 
              if (1)$display("Assertion failed: 'B' channel Get contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_56&io_in_b_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'B' channel Get is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_57)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_57&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_57&(|_GEN_53))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_57&(|io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_57&_GEN_55)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&(|_GEN_53))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&(|io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&(|(io_in_b_bits_mask&~mask_1)))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&(|_GEN_53))
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&_GEN_55)
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Logical type unsupported by client (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&(|_GEN_53))
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&_GEN_55)
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Hint type unsupported by client (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&(|_GEN_53))
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&_GEN_55)
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&io_in_b_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&_GEN_70)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&(|_GEN_62))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_69&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&_GEN_70)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(|_GEN_62))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&~_GEN_73)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&~_GEN_75)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&_GEN_70)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&(|_GEN_62))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_74&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&~_GEN_73)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&~_GEN_75)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&_GEN_70)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&(|_GEN_62))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_77&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_77&(|_GEN_62))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_77&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&(|_GEN_62))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_79&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_79&(|_GEN_62))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_79&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_b_bits_opcode!=opcode_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_b_bits_param!=param_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_b_bits_size!=size_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_b_bits_source!=source_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_b_bits_address!=address_1)
            begin 
              if (1)$display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_c_bits_opcode!=opcode_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_c_bits_param!=param_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_c_bits_size!=size_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_c_bits_source!=source_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_c_bits_address!=address_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel address changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_92[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_86&~reset&~(_GEN_93[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_87&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_87&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_88&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_88&_GEN_89!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_85&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_86 ? 2'h1<<_GEN_3:2'h0)|a_set_wo_ready==2'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==2'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~reset&_GEN_94[0])
            begin 
              if (1)$display("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_91&~reset&~(_GEN_95[0]|same_cycle_resp_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_91&same_cycle_resp_1&~reset&io_in_d_bits_size!=io_in_c_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_91&~same_cycle_resp_1&~reset&_GEN_89!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_90&c_first_1&io_in_c_valid&io_in_c_bits_source==io_in_d_bits_source&d_release_ack&~(io_in_c_bits_opcode==3'h4|io_in_c_bits_opcode==3'h5)&~reset&~(~io_in_d_ready|io_in_c_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if ((|c_set_wo_ready)&~reset&c_set_wo_ready==(_GEN_91 ? 2'h1<<_GEN_3:2'h0))
            begin 
              if (1)$display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==2'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~reset&_GEN_96[0])
            begin 
              if (1)$display("Assertion failed: 'D' channel re-used a sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~reset&~(_GEN_97[0]))
            begin 
              if (1)$display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_98={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_98 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_98 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_98 ;  
   wire [26:0] _d_first_beats1_decode_T_13=27'hFFF<<_GEN_98 ;  
   wire [26:0] _c_first_beats1_decode_T_1=27'hFFF<<_GEN_0 ;  
   wire [26:0] _c_first_beats1_decode_T_5=27'hFFF<<_GEN_0 ;  
   wire _GEN_99=_d_first_T_3&d_first_1&~d_release_ack ;  
   wire [30:0] _GEN_100={27'h0,io_in_d_bits_source,3'h0} ;  
   wire _GEN_101=_d_first_T_3&d_first_2&d_release_ack ;  
   wire [30:0] _d_opcodes_clr_T_5=31'hF<<{28'h0,io_in_d_bits_source,2'h0} ;  
   wire [18:0] _a_opcodes_set_T_1={15'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{16'h0,io_in_a_bits_source,2'h0} ;  
   wire [30:0] _d_sizes_clr_T_5=31'hFF<<_GEN_100 ;  
   wire [19:0] _a_sizes_set_T_1={15'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:5'h0}<<{16'h0,io_in_a_bits_source,3'h0} ;  
   wire [30:0] _d_sizes_clr_T_11=31'hFF<<_GEN_100 ;  
   wire [19:0] _c_sizes_set_T_1={15'h0,_GEN_6 ? {io_in_c_bits_size,1'h1}:5'h0}<<{16'h0,io_in_c_bits_source,3'h0} ;  
   wire b_first_done=io_in_b_ready&io_in_b_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              b_first_counter <=9'h0;
              c_first_counter <=9'h0;
              inflight <=2'h0;
              inflight_opcodes <=8'h0;
              inflight_sizes <=16'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=2'h0;
              inflight_sizes_1 <=16'h0;
              c_first_counter_1 <=9'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
              inflight_2 <=4'h0;
              d_first_counter_3 <=9'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_3)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   if (d_first_3)
                      d_first_counter_3 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_13[11:3]):9'h0;
                    else 
                      d_first_counter_3 <=d_first_counter_3-9'h1;
                 end 
              if (b_first_done)
                 begin 
                   if (|b_first_counter)
                      b_first_counter <=b_first_counter-9'h1;
                    else 
                      b_first_counter <=9'h0;
                 end 
              if (_c_first_T_1)
                 begin 
                   if (|c_first_counter)
                      c_first_counter <=c_first_counter-9'h1;
                    else 
                      c_first_counter <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_1[11:3]):9'h0;
                   if (c_first_1)
                      c_first_counter_1 <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      c_first_counter_1 <=c_first_counter_1-9'h1;
                 end 
              inflight <=(inflight|(_GEN_2 ? 2'h1<<_GEN_1:2'h0))&~(_GEN_99 ? 2'h1<<_GEN_3:2'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[7:0]:8'h0))&~(_GEN_99 ? _d_opcodes_clr_T_5[7:0]:8'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[15:0]:16'h0))&~(_GEN_99 ? _d_sizes_clr_T_5[15:0]:16'h0);
              if (_a_first_T_1|_d_first_T_3)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=(inflight_1|(_GEN_6 ? 2'h1<<_GEN_5:2'h0))&~(_GEN_101 ? 2'h1<<_GEN_3:2'h0);
              inflight_sizes_1 <=(inflight_sizes_1|(_GEN_6 ? _c_sizes_set_T_1[15:0]:16'h0))&~(_GEN_101 ? _d_sizes_clr_T_11[15:0]:16'h0);
              if (_c_first_T_1|_d_first_T_3)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight_2 <=(inflight_2|d_set)&~(_GEN_9 ? 4'h1<<_GEN_10:4'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_3&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
         if (b_first_done&~(|b_first_counter))
            begin 
              opcode_2 <=io_in_b_bits_opcode;
              param_2 <=io_in_b_bits_param;
              size_2 <=io_in_b_bits_size;
              source_2 <=io_in_b_bits_source;
              address_1 <=io_in_b_bits_address;
            end 
         if (_c_first_T_1&~(|c_first_counter))
            begin 
              opcode_3 <=io_in_c_bits_opcode;
              param_3 <=io_in_c_bits_param;
              size_3 <=io_in_c_bits_size;
              source_3 <=io_in_c_bits_source;
              address_2 <=io_in_c_bits_address;
            end 
       end
  
endmodule
 
module TLMonitor_24 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [31:0] io_in_a_bits_address,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [31:0] address ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg inflight ;  
   reg [3:0] inflight_opcodes ;  
   reg [7:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire a_set=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire _GEN=io_in_d_valid&d_first_1 ;  
   wire d_clr=_GEN&~d_release_ack ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg inflight_1 ;  
   reg [7:0] inflight_sizes_1 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   wire d_clr_1=io_in_d_valid&d_first_2&d_release_ack ;  
   reg [31:0] watchdog_1 ;  
   wire _GEN_0=io_in_a_valid&~reset ;  
   wire _GEN_1=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_2=io_in_d_bits_size<4'h3 ;  
   wire _GEN_3=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_4=io_in_d_bits_param==2'h2 ;  
   wire _GEN_5=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_6=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_7=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_8=io_in_d_bits_opcode==3'h1 ;  
   wire _GEN_9=io_in_d_valid&_GEN_8&~reset ;  
   wire _GEN_10=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_11=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire a_set_wo_ready=io_in_a_valid&a_first_1 ;  
   wire _GEN_12=d_clr&a_set_wo_ready&~reset ;  
   wire _GEN_13=d_clr&~a_set_wo_ready&~reset ;  
   wire [7:0] _GEN_14={4'h0,io_in_d_bits_size} ;  
   wire _GEN_15=d_clr_1&~reset ;  
  always @( posedge clock)
       begin 
         if (_GEN_0&~({io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0|io_in_a_bits_address[31:12]==20'h0|{io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0|{io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0|{io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0|{io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0|io_in_a_bits_address[31:28]==4'h8))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&(|(io_in_a_bits_address[5:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_a_valid&(|a_first_counter)&~reset&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (a_set&~reset&inflight)
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (d_clr&~reset&~(inflight|a_set_wo_ready))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_d_bits_size!=4'h6)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_14!={1'h0,inflight_sizes[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN&a_first_1&io_in_a_valid&~d_release_ack&~reset&~io_in_a_ready)
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=d_clr|~a_set_wo_ready))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~inflight_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_14!={1'h0,inflight_sizes_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight_1|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _GEN_16={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_16 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_16 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_16 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              inflight <=1'h0;
              inflight_opcodes <=4'h0;
              inflight_sizes <=8'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=1'h0;
              inflight_sizes_1 <=8'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=9'h0;
                   if (a_first_1)
                      a_first_counter_1 <=9'h0;
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (io_in_d_valid)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   watchdog_1 <=32'h0;
                 end 
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight <=(inflight|a_set)&~d_clr;
              inflight_opcodes <=(inflight_opcodes|(a_set ? 4'h9:4'h0))&~{4{d_clr}};
              inflight_sizes <=(inflight_sizes|(a_set ? {3'h0,a_set ? 5'hD:5'h0}:8'h0))&~{8{d_clr}};
              if (_a_first_T_1|io_in_d_valid)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~d_clr_1;
              inflight_sizes_1 <=inflight_sizes_1&~{8{d_clr_1}};
            end 
         if (_a_first_T_1&~(|a_first_counter))
            address <=io_in_a_bits_address;
         if (io_in_d_valid&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLXbar_8 (
  input clock,
  input reset,
  output auto_in_1_a_ready,
  input auto_in_1_a_valid,
  input [31:0] auto_in_1_a_bits_address,
  output auto_in_1_d_valid,
  output [2:0] auto_in_1_d_bits_opcode,
  output [3:0] auto_in_1_d_bits_size,
  output [63:0] auto_in_1_d_bits_data,
  output auto_in_1_d_bits_corrupt,
  output auto_in_0_a_ready,
  input auto_in_0_a_valid,
  input [2:0] auto_in_0_a_bits_opcode,
  input [2:0] auto_in_0_a_bits_param,
  input [3:0] auto_in_0_a_bits_size,
  input auto_in_0_a_bits_source,
  input [31:0] auto_in_0_a_bits_address,
  input [7:0] auto_in_0_a_bits_mask,
  input [63:0] auto_in_0_a_bits_data,
  input auto_in_0_b_ready,
  output auto_in_0_b_valid,
  output [1:0] auto_in_0_b_bits_param,
  output [3:0] auto_in_0_b_bits_size,
  output auto_in_0_b_bits_source,
  output [31:0] auto_in_0_b_bits_address,
  output auto_in_0_c_ready,
  input auto_in_0_c_valid,
  input [2:0] auto_in_0_c_bits_opcode,
  input [2:0] auto_in_0_c_bits_param,
  input [3:0] auto_in_0_c_bits_size,
  input auto_in_0_c_bits_source,
  input [31:0] auto_in_0_c_bits_address,
  input [63:0] auto_in_0_c_bits_data,
  input auto_in_0_d_ready,
  output auto_in_0_d_valid,
  output [2:0] auto_in_0_d_bits_opcode,
  output [1:0] auto_in_0_d_bits_param,
  output [3:0] auto_in_0_d_bits_size,
  output auto_in_0_d_bits_source,
  output [1:0] auto_in_0_d_bits_sink,
  output auto_in_0_d_bits_denied,
  output [63:0] auto_in_0_d_bits_data,
  output auto_in_0_e_ready,
  input auto_in_0_e_valid,
  input [1:0] auto_in_0_e_bits_sink,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [1:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [2:0] auto_out_b_bits_opcode,
  input [1:0] auto_out_b_bits_param,
  input [3:0] auto_out_b_bits_size,
  input [1:0] auto_out_b_bits_source,
  input [31:0] auto_out_b_bits_address,
  input [7:0] auto_out_b_bits_mask,
  input auto_out_b_bits_corrupt,
  input auto_out_c_ready,
  output auto_out_c_valid,
  output [2:0] auto_out_c_bits_opcode,
  output [2:0] auto_out_c_bits_param,
  output [3:0] auto_out_c_bits_size,
  output [1:0] auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [1:0] auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt,
  input auto_out_e_ready,
  output auto_out_e_valid,
  output [1:0] auto_out_e_bits_sink) ; 
   wire requestDOI_0_1=auto_out_d_bits_source==2'h2 ;  
   wire portsBIO_filtered_valid_0=auto_out_b_valid&~(auto_out_b_bits_source[1]) ;  
   wire portsDIO_filtered_0_valid=auto_out_d_valid&~(auto_out_d_bits_source[1]) ;  
   wire portsDIO_filtered_1_valid=auto_out_d_valid&requestDOI_0_1 ;  
   reg [8:0] beatsLeft ;  
   wire idle=beatsLeft==9'h0 ;  
   wire [1:0] readys_valid={auto_in_1_a_valid,auto_in_0_a_valid} ;  
   reg [1:0] readys_mask ;  
   wire [1:0] _readys_filter_T_1=readys_valid&~readys_mask ;  
   wire [1:0] readys_readys=~({readys_mask[1],_readys_filter_T_1[1]|readys_mask[0]}&({_readys_filter_T_1[0],auto_in_1_a_valid}|_readys_filter_T_1)) ;  
   wire winner_0=readys_readys[0]&auto_in_0_a_valid ;  
   wire winner_1=readys_readys[1]&auto_in_1_a_valid ;  
   wire _out_0_a_valid_T=auto_in_0_a_valid|auto_in_1_a_valid ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~winner_0|~winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_out_0_a_valid_T|winner_0|winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg state_0 ;  
   reg state_1 ;  
   wire muxState_0=idle ? winner_0:state_0 ;  
   wire muxState_1=idle ? winner_1:state_1 ;  
   wire portsAOI_filtered_0_ready=auto_out_a_ready&(idle ? readys_readys[0]:state_0) ;  
   wire portsAOI_filtered_1_0_ready=auto_out_a_ready&(idle ? readys_readys[1]:state_1) ;  
   wire out_0_a_valid=idle ? _out_0_a_valid_T:state_0&auto_in_0_a_valid|state_1&auto_in_1_a_valid ;  
   wire [26:0] _beatsAI_decode_T_1=27'hFFF<<auto_in_0_a_bits_size ;  
   wire [1:0] _readys_mask_T=readys_readys&readys_valid ;  
   wire latch=idle&auto_out_a_ready ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              beatsLeft <=9'h0;
              readys_mask <=2'h3;
              state_0 <=1'h0;
              state_1 <=1'h0;
            end 
          else 
            begin 
              if (latch)
                 beatsLeft <=winner_0&~(auto_in_0_a_bits_opcode[2]) ? ~(_beatsAI_decode_T_1[11:3]):9'h0;
               else 
                 beatsLeft <=beatsLeft-{8'h0,auto_out_a_ready&out_0_a_valid};
              if (latch&(|readys_valid))
                 readys_mask <=_readys_mask_T|{_readys_mask_T[0],1'h0};
              if (idle)
                 begin 
                   state_0 <=winner_0;
                   state_1 <=winner_1;
                 end 
            end 
       end
  
  TLMonitor_23 monitor(.clock(clock),.reset(reset),.io_in_a_ready(portsAOI_filtered_0_ready),.io_in_a_valid(auto_in_0_a_valid),.io_in_a_bits_opcode(auto_in_0_a_bits_opcode),.io_in_a_bits_param(auto_in_0_a_bits_param),.io_in_a_bits_size(auto_in_0_a_bits_size),.io_in_a_bits_source(auto_in_0_a_bits_source),.io_in_a_bits_address(auto_in_0_a_bits_address),.io_in_a_bits_mask(auto_in_0_a_bits_mask),.io_in_b_ready(auto_in_0_b_ready),.io_in_b_valid(portsBIO_filtered_valid_0),.io_in_b_bits_opcode(auto_out_b_bits_opcode),.io_in_b_bits_param(auto_out_b_bits_param),.io_in_b_bits_size(auto_out_b_bits_size),.io_in_b_bits_source(auto_out_b_bits_source[0]),.io_in_b_bits_address(auto_out_b_bits_address),.io_in_b_bits_mask(auto_out_b_bits_mask),.io_in_b_bits_corrupt(auto_out_b_bits_corrupt),.io_in_c_ready(auto_out_c_ready),.io_in_c_valid(auto_in_0_c_valid),.io_in_c_bits_opcode(auto_in_0_c_bits_opcode),.io_in_c_bits_param(auto_in_0_c_bits_param),.io_in_c_bits_size(auto_in_0_c_bits_size),.io_in_c_bits_source(auto_in_0_c_bits_source),.io_in_c_bits_address(auto_in_0_c_bits_address),.io_in_d_ready(auto_in_0_d_ready),.io_in_d_valid(portsDIO_filtered_0_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_param(auto_out_d_bits_param),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_source(auto_out_d_bits_source[0]),.io_in_d_bits_sink(auto_out_d_bits_sink),.io_in_d_bits_denied(auto_out_d_bits_denied),.io_in_d_bits_corrupt(auto_out_d_bits_corrupt),.io_in_e_ready(auto_out_e_ready),.io_in_e_valid(auto_in_0_e_valid),.io_in_e_bits_sink(auto_in_0_e_bits_sink)); 
  TLMonitor_24 monitor_1(.clock(clock),.reset(reset),.io_in_a_ready(portsAOI_filtered_1_0_ready),.io_in_a_valid(auto_in_1_a_valid),.io_in_a_bits_address(auto_in_1_a_bits_address),.io_in_d_valid(portsDIO_filtered_1_valid),.io_in_d_bits_opcode(auto_out_d_bits_opcode),.io_in_d_bits_param(auto_out_d_bits_param),.io_in_d_bits_size(auto_out_d_bits_size),.io_in_d_bits_sink(auto_out_d_bits_sink),.io_in_d_bits_denied(auto_out_d_bits_denied),.io_in_d_bits_corrupt(auto_out_d_bits_corrupt)); 
  assign auto_in_1_a_ready=portsAOI_filtered_1_0_ready; 
  assign auto_in_1_d_valid=portsDIO_filtered_1_valid; 
  assign auto_in_1_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_1_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_1_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_1_d_bits_corrupt=auto_out_d_bits_corrupt; 
  assign auto_in_0_a_ready=portsAOI_filtered_0_ready; 
  assign auto_in_0_b_valid=portsBIO_filtered_valid_0; 
  assign auto_in_0_b_bits_param=auto_out_b_bits_param; 
  assign auto_in_0_b_bits_size=auto_out_b_bits_size; 
  assign auto_in_0_b_bits_source=auto_out_b_bits_source[0]; 
  assign auto_in_0_b_bits_address=auto_out_b_bits_address; 
  assign auto_in_0_c_ready=auto_out_c_ready; 
  assign auto_in_0_d_valid=portsDIO_filtered_0_valid; 
  assign auto_in_0_d_bits_opcode=auto_out_d_bits_opcode; 
  assign auto_in_0_d_bits_param=auto_out_d_bits_param; 
  assign auto_in_0_d_bits_size=auto_out_d_bits_size; 
  assign auto_in_0_d_bits_source=auto_out_d_bits_source[0]; 
  assign auto_in_0_d_bits_sink=auto_out_d_bits_sink; 
  assign auto_in_0_d_bits_denied=auto_out_d_bits_denied; 
  assign auto_in_0_d_bits_data=auto_out_d_bits_data; 
  assign auto_in_0_e_ready=auto_out_e_ready; 
  assign auto_out_a_valid=out_0_a_valid; 
  assign auto_out_a_bits_opcode=(muxState_0 ? auto_in_0_a_bits_opcode:3'h0)|{muxState_1,2'h0}; 
  assign auto_out_a_bits_param=muxState_0 ? auto_in_0_a_bits_param:3'h0; 
  assign auto_out_a_bits_size=(muxState_0 ? auto_in_0_a_bits_size:4'h0)|(muxState_1 ? 4'h6:4'h0); 
  assign auto_out_a_bits_source=(muxState_0 ? {1'h0,auto_in_0_a_bits_source}:2'h0)|{muxState_1,1'h0}; 
  assign auto_out_a_bits_address=(muxState_0 ? auto_in_0_a_bits_address:32'h0)|(muxState_1 ? auto_in_1_a_bits_address:32'h0); 
  assign auto_out_a_bits_mask=(muxState_0 ? auto_in_0_a_bits_mask:8'h0)|{8{muxState_1}}; 
  assign auto_out_a_bits_data=muxState_0 ? auto_in_0_a_bits_data:64'h0; 
  assign auto_out_b_ready=~(auto_out_b_bits_source[1])&auto_in_0_b_ready; 
  assign auto_out_c_valid=auto_in_0_c_valid; 
  assign auto_out_c_bits_opcode=auto_in_0_c_bits_opcode; 
  assign auto_out_c_bits_param=auto_in_0_c_bits_param; 
  assign auto_out_c_bits_size=auto_in_0_c_bits_size; 
  assign auto_out_c_bits_source={1'h0,auto_in_0_c_bits_source}; 
  assign auto_out_c_bits_address=auto_in_0_c_bits_address; 
  assign auto_out_c_bits_data=auto_in_0_c_bits_data; 
  assign auto_out_d_ready=~(auto_out_d_bits_source[1])&auto_in_0_d_ready|requestDOI_0_1; 
  assign auto_out_e_valid=auto_in_0_e_valid; 
  assign auto_out_e_bits_sink=auto_in_0_e_bits_sink; 
endmodule
 
module IntXbar_1 (
  input auto_int_in_2_0,
  input auto_int_in_1_0,
  input auto_int_in_1_1,
  input auto_int_in_0_0,
  output auto_int_out_0,
  output auto_int_out_1,
  output auto_int_out_2,
  output auto_int_out_3) ; 
  assign auto_int_out_0=auto_int_in_0_0; 
  assign auto_int_out_1=auto_int_in_1_0; 
  assign auto_int_out_2=auto_int_in_1_1; 
  assign auto_int_out_3=auto_int_in_2_0; 
endmodule
 
module OptimizationBarrier (
  input io_x_u,
  input io_x_ae_ptw,
  input io_x_ae_final,
  input io_x_pf,
  input io_x_gf,
  input io_x_sw,
  input io_x_sx,
  input io_x_sr,
  input io_x_pw,
  input io_x_px,
  input io_x_pr,
  input io_x_ppp,
  input io_x_pal,
  input io_x_paa,
  input io_x_eff,
  input io_x_c,
  output io_y_u,
  output io_y_ae_ptw,
  output io_y_ae_final,
  output io_y_pf,
  output io_y_gf,
  output io_y_sw,
  output io_y_sx,
  output io_y_sr,
  output io_y_pw,
  output io_y_px,
  output io_y_pr,
  output io_y_ppp,
  output io_y_pal,
  output io_y_paa,
  output io_y_eff,
  output io_y_c) ; 
  assign io_y_u=io_x_u; 
  assign io_y_ae_ptw=io_x_ae_ptw; 
  assign io_y_ae_final=io_x_ae_final; 
  assign io_y_pf=io_x_pf; 
  assign io_y_gf=io_x_gf; 
  assign io_y_sw=io_x_sw; 
  assign io_y_sx=io_x_sx; 
  assign io_y_sr=io_x_sr; 
  assign io_y_pw=io_x_pw; 
  assign io_y_px=io_x_px; 
  assign io_y_pr=io_x_pr; 
  assign io_y_ppp=io_x_ppp; 
  assign io_y_pal=io_x_pal; 
  assign io_y_paa=io_x_paa; 
  assign io_y_eff=io_x_eff; 
  assign io_y_c=io_x_c; 
endmodule
 
module PMPChecker (
  input [1:0] io_prv,
  input io_pmp_cfg_l_0,
  input io_pmp_cfg_l_1,
  input io_pmp_cfg_l_2,
  input io_pmp_cfg_l_3,
  input io_pmp_cfg_l_4,
  input io_pmp_cfg_l_5,
  input io_pmp_cfg_l_6,
  input io_pmp_cfg_l_7,
  input [1:0] io_pmp_cfg_a_0,
  input [1:0] io_pmp_cfg_a_1,
  input [1:0] io_pmp_cfg_a_2,
  input [1:0] io_pmp_cfg_a_3,
  input [1:0] io_pmp_cfg_a_4,
  input [1:0] io_pmp_cfg_a_5,
  input [1:0] io_pmp_cfg_a_6,
  input [1:0] io_pmp_cfg_a_7,
  input io_pmp_cfg_w_0,
  input io_pmp_cfg_w_1,
  input io_pmp_cfg_w_2,
  input io_pmp_cfg_w_3,
  input io_pmp_cfg_w_4,
  input io_pmp_cfg_w_5,
  input io_pmp_cfg_w_6,
  input io_pmp_cfg_w_7,
  input io_pmp_cfg_r_0,
  input io_pmp_cfg_r_1,
  input io_pmp_cfg_r_2,
  input io_pmp_cfg_r_3,
  input io_pmp_cfg_r_4,
  input io_pmp_cfg_r_5,
  input io_pmp_cfg_r_6,
  input io_pmp_cfg_r_7,
  input [29:0] io_pmp_addr_0,
  input [29:0] io_pmp_addr_1,
  input [29:0] io_pmp_addr_2,
  input [29:0] io_pmp_addr_3,
  input [29:0] io_pmp_addr_4,
  input [29:0] io_pmp_addr_5,
  input [29:0] io_pmp_addr_6,
  input [29:0] io_pmp_addr_7,
  input [31:0] io_pmp_mask_0,
  input [31:0] io_pmp_mask_1,
  input [31:0] io_pmp_mask_2,
  input [31:0] io_pmp_mask_3,
  input [31:0] io_pmp_mask_4,
  input [31:0] io_pmp_mask_5,
  input [31:0] io_pmp_mask_6,
  input [31:0] io_pmp_mask_7,
  input [31:0] io_addr,
  input [1:0] io_size,
  output io_r,
  output io_w) ; 
   wire [5:0] _GEN={4'h0,io_size} ;  
   wire [5:0] _res_hit_lsbMask_T_1=6'h7<<_GEN ;  
   wire [5:0] _res_hit_T_4=6'h7<<_GEN ;  
   wire res_hit=io_pmp_cfg_a_7[1] ? ((io_addr[31:3]^io_pmp_addr_7[29:1])&~(io_pmp_mask_7[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_7[0],2'h0})&~(io_pmp_mask_7[2:0]|~(_res_hit_lsbMask_T_1[2:0])))==3'h0:io_pmp_cfg_a_7[0]&~(io_addr[31:3]<io_pmp_addr_6[29:1]|(io_addr[31:3]^io_pmp_addr_6[29:1])==29'h0&(io_addr[2:0]|~(_res_hit_T_4[2:0]))<{io_pmp_addr_6[0],2'h0})&(io_addr[31:3]<io_pmp_addr_7[29:1]|(io_addr[31:3]^io_pmp_addr_7[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_7[0],2'h0}) ;  
   wire res_ignore=io_prv[1]&~io_pmp_cfg_l_7 ;  
   wire [5:0] _res_aligned_lsbMask_T_1=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask=~(_res_aligned_lsbMask_T_1[2:0]) ;  
   wire res_aligned=io_pmp_cfg_a_7[1] ? (res_aligned_lsbMask&~(io_pmp_mask_7[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_6[29:1])==29'h0&io_pmp_addr_6[0]&~(io_addr[2])|(io_addr[31:3]^io_pmp_addr_7[29:1])==29'h0&io_pmp_addr_7[0]&(io_addr[2]|res_aligned_lsbMask[2])) ;  
   wire [5:0] _res_hit_lsbMask_T_5=6'h7<<_GEN ;  
   wire [5:0] _res_hit_T_18=6'h7<<_GEN ;  
   wire res_hit_1=io_pmp_cfg_a_6[1] ? ((io_addr[31:3]^io_pmp_addr_6[29:1])&~(io_pmp_mask_6[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_6[0],2'h0})&~(io_pmp_mask_6[2:0]|~(_res_hit_lsbMask_T_5[2:0])))==3'h0:io_pmp_cfg_a_6[0]&~(io_addr[31:3]<io_pmp_addr_5[29:1]|(io_addr[31:3]^io_pmp_addr_5[29:1])==29'h0&(io_addr[2:0]|~(_res_hit_T_18[2:0]))<{io_pmp_addr_5[0],2'h0})&(io_addr[31:3]<io_pmp_addr_6[29:1]|(io_addr[31:3]^io_pmp_addr_6[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_6[0],2'h0}) ;  
   wire res_ignore_1=io_prv[1]&~io_pmp_cfg_l_6 ;  
   wire [5:0] _res_aligned_lsbMask_T_4=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask_1=~(_res_aligned_lsbMask_T_4[2:0]) ;  
   wire res_aligned_1=io_pmp_cfg_a_6[1] ? (res_aligned_lsbMask_1&~(io_pmp_mask_6[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_5[29:1])==29'h0&io_pmp_addr_5[0]&~(io_addr[2])|(io_addr[31:3]^io_pmp_addr_6[29:1])==29'h0&io_pmp_addr_6[0]&(io_addr[2]|res_aligned_lsbMask_1[2])) ;  
   wire [5:0] _res_hit_lsbMask_T_9=6'h7<<_GEN ;  
   wire [5:0] _res_hit_T_32=6'h7<<_GEN ;  
   wire res_hit_2=io_pmp_cfg_a_5[1] ? ((io_addr[31:3]^io_pmp_addr_5[29:1])&~(io_pmp_mask_5[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_5[0],2'h0})&~(io_pmp_mask_5[2:0]|~(_res_hit_lsbMask_T_9[2:0])))==3'h0:io_pmp_cfg_a_5[0]&~(io_addr[31:3]<io_pmp_addr_4[29:1]|(io_addr[31:3]^io_pmp_addr_4[29:1])==29'h0&(io_addr[2:0]|~(_res_hit_T_32[2:0]))<{io_pmp_addr_4[0],2'h0})&(io_addr[31:3]<io_pmp_addr_5[29:1]|(io_addr[31:3]^io_pmp_addr_5[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_5[0],2'h0}) ;  
   wire res_ignore_2=io_prv[1]&~io_pmp_cfg_l_5 ;  
   wire [5:0] _res_aligned_lsbMask_T_7=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask_2=~(_res_aligned_lsbMask_T_7[2:0]) ;  
   wire res_aligned_2=io_pmp_cfg_a_5[1] ? (res_aligned_lsbMask_2&~(io_pmp_mask_5[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_4[29:1])==29'h0&io_pmp_addr_4[0]&~(io_addr[2])|(io_addr[31:3]^io_pmp_addr_5[29:1])==29'h0&io_pmp_addr_5[0]&(io_addr[2]|res_aligned_lsbMask_2[2])) ;  
   wire [5:0] _res_hit_lsbMask_T_13=6'h7<<_GEN ;  
   wire [5:0] _res_hit_T_46=6'h7<<_GEN ;  
   wire res_hit_3=io_pmp_cfg_a_4[1] ? ((io_addr[31:3]^io_pmp_addr_4[29:1])&~(io_pmp_mask_4[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_4[0],2'h0})&~(io_pmp_mask_4[2:0]|~(_res_hit_lsbMask_T_13[2:0])))==3'h0:io_pmp_cfg_a_4[0]&~(io_addr[31:3]<io_pmp_addr_3[29:1]|(io_addr[31:3]^io_pmp_addr_3[29:1])==29'h0&(io_addr[2:0]|~(_res_hit_T_46[2:0]))<{io_pmp_addr_3[0],2'h0})&(io_addr[31:3]<io_pmp_addr_4[29:1]|(io_addr[31:3]^io_pmp_addr_4[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_4[0],2'h0}) ;  
   wire res_ignore_3=io_prv[1]&~io_pmp_cfg_l_4 ;  
   wire [5:0] _res_aligned_lsbMask_T_10=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask_3=~(_res_aligned_lsbMask_T_10[2:0]) ;  
   wire res_aligned_3=io_pmp_cfg_a_4[1] ? (res_aligned_lsbMask_3&~(io_pmp_mask_4[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_3[29:1])==29'h0&io_pmp_addr_3[0]&~(io_addr[2])|(io_addr[31:3]^io_pmp_addr_4[29:1])==29'h0&io_pmp_addr_4[0]&(io_addr[2]|res_aligned_lsbMask_3[2])) ;  
   wire [5:0] _res_hit_lsbMask_T_17=6'h7<<_GEN ;  
   wire [5:0] _res_hit_T_60=6'h7<<_GEN ;  
   wire res_hit_4=io_pmp_cfg_a_3[1] ? ((io_addr[31:3]^io_pmp_addr_3[29:1])&~(io_pmp_mask_3[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_3[0],2'h0})&~(io_pmp_mask_3[2:0]|~(_res_hit_lsbMask_T_17[2:0])))==3'h0:io_pmp_cfg_a_3[0]&~(io_addr[31:3]<io_pmp_addr_2[29:1]|(io_addr[31:3]^io_pmp_addr_2[29:1])==29'h0&(io_addr[2:0]|~(_res_hit_T_60[2:0]))<{io_pmp_addr_2[0],2'h0})&(io_addr[31:3]<io_pmp_addr_3[29:1]|(io_addr[31:3]^io_pmp_addr_3[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_3[0],2'h0}) ;  
   wire res_ignore_4=io_prv[1]&~io_pmp_cfg_l_3 ;  
   wire [5:0] _res_aligned_lsbMask_T_13=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask_4=~(_res_aligned_lsbMask_T_13[2:0]) ;  
   wire res_aligned_4=io_pmp_cfg_a_3[1] ? (res_aligned_lsbMask_4&~(io_pmp_mask_3[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_2[29:1])==29'h0&io_pmp_addr_2[0]&~(io_addr[2])|(io_addr[31:3]^io_pmp_addr_3[29:1])==29'h0&io_pmp_addr_3[0]&(io_addr[2]|res_aligned_lsbMask_4[2])) ;  
   wire [5:0] _res_hit_lsbMask_T_21=6'h7<<_GEN ;  
   wire [5:0] _res_hit_T_74=6'h7<<_GEN ;  
   wire res_hit_5=io_pmp_cfg_a_2[1] ? ((io_addr[31:3]^io_pmp_addr_2[29:1])&~(io_pmp_mask_2[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_2[0],2'h0})&~(io_pmp_mask_2[2:0]|~(_res_hit_lsbMask_T_21[2:0])))==3'h0:io_pmp_cfg_a_2[0]&~(io_addr[31:3]<io_pmp_addr_1[29:1]|(io_addr[31:3]^io_pmp_addr_1[29:1])==29'h0&(io_addr[2:0]|~(_res_hit_T_74[2:0]))<{io_pmp_addr_1[0],2'h0})&(io_addr[31:3]<io_pmp_addr_2[29:1]|(io_addr[31:3]^io_pmp_addr_2[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_2[0],2'h0}) ;  
   wire res_ignore_5=io_prv[1]&~io_pmp_cfg_l_2 ;  
   wire [5:0] _res_aligned_lsbMask_T_16=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask_5=~(_res_aligned_lsbMask_T_16[2:0]) ;  
   wire res_aligned_5=io_pmp_cfg_a_2[1] ? (res_aligned_lsbMask_5&~(io_pmp_mask_2[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_1[29:1])==29'h0&io_pmp_addr_1[0]&~(io_addr[2])|(io_addr[31:3]^io_pmp_addr_2[29:1])==29'h0&io_pmp_addr_2[0]&(io_addr[2]|res_aligned_lsbMask_5[2])) ;  
   wire [5:0] _res_hit_lsbMask_T_25=6'h7<<_GEN ;  
   wire [5:0] _res_hit_T_88=6'h7<<_GEN ;  
   wire res_hit_6=io_pmp_cfg_a_1[1] ? ((io_addr[31:3]^io_pmp_addr_1[29:1])&~(io_pmp_mask_1[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_1[0],2'h0})&~(io_pmp_mask_1[2:0]|~(_res_hit_lsbMask_T_25[2:0])))==3'h0:io_pmp_cfg_a_1[0]&~(io_addr[31:3]<io_pmp_addr_0[29:1]|(io_addr[31:3]^io_pmp_addr_0[29:1])==29'h0&(io_addr[2:0]|~(_res_hit_T_88[2:0]))<{io_pmp_addr_0[0],2'h0})&(io_addr[31:3]<io_pmp_addr_1[29:1]|(io_addr[31:3]^io_pmp_addr_1[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_1[0],2'h0}) ;  
   wire res_ignore_6=io_prv[1]&~io_pmp_cfg_l_1 ;  
   wire [5:0] _res_aligned_lsbMask_T_19=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask_6=~(_res_aligned_lsbMask_T_19[2:0]) ;  
   wire res_aligned_6=io_pmp_cfg_a_1[1] ? (res_aligned_lsbMask_6&~(io_pmp_mask_1[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_0[29:1])==29'h0&io_pmp_addr_0[0]&~(io_addr[2])|(io_addr[31:3]^io_pmp_addr_1[29:1])==29'h0&io_pmp_addr_1[0]&(io_addr[2]|res_aligned_lsbMask_6[2])) ;  
   wire [5:0] _res_hit_lsbMask_T_29=6'h7<<_GEN ;  
   wire res_hit_7=io_pmp_cfg_a_0[1] ? ((io_addr[31:3]^io_pmp_addr_0[29:1])&~(io_pmp_mask_0[31:3]))==29'h0&((io_addr[2:0]^{io_pmp_addr_0[0],2'h0})&~(io_pmp_mask_0[2:0]|~(_res_hit_lsbMask_T_29[2:0])))==3'h0:io_pmp_cfg_a_0[0]&(io_addr[31:3]<io_pmp_addr_0[29:1]|(io_addr[31:3]^io_pmp_addr_0[29:1])==29'h0&io_addr[2:0]<{io_pmp_addr_0[0],2'h0}) ;  
   wire res_ignore_7=io_prv[1]&~io_pmp_cfg_l_0 ;  
   wire [5:0] _res_aligned_lsbMask_T_22=6'h7<<_GEN ;  
   wire [2:0] res_aligned_lsbMask_7=~(_res_aligned_lsbMask_T_22[2:0]) ;  
   wire res_aligned_7=io_pmp_cfg_a_0[1] ? (res_aligned_lsbMask_7&~(io_pmp_mask_0[2:0]))==3'h0:~((io_addr[31:3]^io_pmp_addr_0[29:1])==29'h0&io_pmp_addr_0[0]&(io_addr[2]|res_aligned_lsbMask_7[2])) ;  
  assign io_r=res_hit_7 ? res_aligned_7&(io_pmp_cfg_r_0|res_ignore_7):res_hit_6 ? res_aligned_6&(io_pmp_cfg_r_1|res_ignore_6):res_hit_5 ? res_aligned_5&(io_pmp_cfg_r_2|res_ignore_5):res_hit_4 ? res_aligned_4&(io_pmp_cfg_r_3|res_ignore_4):res_hit_3 ? res_aligned_3&(io_pmp_cfg_r_4|res_ignore_3):res_hit_2 ? res_aligned_2&(io_pmp_cfg_r_5|res_ignore_2):res_hit_1 ? res_aligned_1&(io_pmp_cfg_r_6|res_ignore_1):res_hit ? res_aligned&(io_pmp_cfg_r_7|res_ignore):io_prv[1]; 
  assign io_w=res_hit_7 ? res_aligned_7&(io_pmp_cfg_w_0|res_ignore_7):res_hit_6 ? res_aligned_6&(io_pmp_cfg_w_1|res_ignore_6):res_hit_5 ? res_aligned_5&(io_pmp_cfg_w_2|res_ignore_5):res_hit_4 ? res_aligned_4&(io_pmp_cfg_w_3|res_ignore_4):res_hit_3 ? res_aligned_3&(io_pmp_cfg_w_4|res_ignore_3):res_hit_2 ? res_aligned_2&(io_pmp_cfg_w_5|res_ignore_2):res_hit_1 ? res_aligned_1&(io_pmp_cfg_w_6|res_ignore_1):res_hit ? res_aligned&(io_pmp_cfg_w_7|res_ignore):io_prv[1]; 
endmodule
 
module data_arrays_0_512x64 (
  input [8:0] RW0_addr,
  input RW0_en,
  input RW0_clk,
  input RW0_wmode,
  input [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input [7:0] RW0_wmask) ; 
   reg [63:0] Memory[0:511] ;  
   reg [8:0] _RW0_raddr_d0 ;  
   reg _RW0_ren_d0 ;  
   reg _RW0_rmode_d0 ;  
  always @( posedge RW0_clk)
       begin 
         _RW0_raddr_d0 <=RW0_addr;
         _RW0_ren_d0 <=RW0_en;
         _RW0_rmode_d0 <=RW0_wmode;
         if (RW0_en&RW0_wmask[0]&RW0_wmode)
            Memory [RW0_addr][32'h0+:8]<=RW0_wdata[7:0];
         if (RW0_en&RW0_wmask[1]&RW0_wmode)
            Memory [RW0_addr][32'h8+:8]<=RW0_wdata[15:8];
         if (RW0_en&RW0_wmask[2]&RW0_wmode)
            Memory [RW0_addr][32'h10+:8]<=RW0_wdata[23:16];
         if (RW0_en&RW0_wmask[3]&RW0_wmode)
            Memory [RW0_addr][32'h18+:8]<=RW0_wdata[31:24];
         if (RW0_en&RW0_wmask[4]&RW0_wmode)
            Memory [RW0_addr][32'h20+:8]<=RW0_wdata[39:32];
         if (RW0_en&RW0_wmask[5]&RW0_wmode)
            Memory [RW0_addr][32'h28+:8]<=RW0_wdata[47:40];
         if (RW0_en&RW0_wmask[6]&RW0_wmode)
            Memory [RW0_addr][32'h30+:8]<=RW0_wdata[55:48];
         if (RW0_en&RW0_wmask[7]&RW0_wmode)
            Memory [RW0_addr][32'h38+:8]<=RW0_wdata[63:56];
       end
  
  assign RW0_rdata=_RW0_ren_d0&~_RW0_rmode_d0 ? Memory[_RW0_raddr_d0]:64'bx; 
endmodule
 
module DCacheDataArray (
  input clock,
  input io_req_valid,
  input [11:0] io_req_bits_addr,
  input io_req_bits_write,
  input [63:0] io_req_bits_wdata,
  input [7:0] io_req_bits_eccMask,
  output [63:0] io_resp_0) ; 
   wire data_arrays_0_rdata_data_en ;  
   wire data_arrays_0_rdata_MPORT_en ;  
  assign data_arrays_0_rdata_MPORT_en=io_req_valid&io_req_bits_write; 
  assign data_arrays_0_rdata_data_en=io_req_valid&~io_req_bits_write; 
  data_arrays_0_512x64 data_arrays_0_ext(.RW0_addr(io_req_bits_addr[11:3]),.RW0_en(data_arrays_0_rdata_data_en|data_arrays_0_rdata_MPORT_en),.RW0_clk(clock),.RW0_wmode(io_req_bits_write),.RW0_wdata(io_req_bits_wdata),.RW0_rdata(io_resp_0),.RW0_wmask(io_req_bits_eccMask)); 
endmodule
 
module AMOALU (
  input [7:0] io_mask,
  input [4:0] io_cmd,
  input [63:0] io_lhs,
  input [63:0] io_rhs,
  output [63:0] io_out) ; 
   wire _logic_xor_T_1=io_cmd==5'hA ;  
   wire logic_and=_logic_xor_T_1|io_cmd==5'hB ;  
   wire logic_xor=io_cmd==5'h9|_logic_xor_T_1 ;  
   wire [63:0] adder_out_mask={32'hFFFFFFFF,io_mask[3],31'h7FFFFFFF} ;  
   wire [63:0] wmask={{8{io_mask[7]}},{8{io_mask[6]}},{8{io_mask[5]}},{8{io_mask[4]}},{8{io_mask[3]}},{8{io_mask[2]}},{8{io_mask[1]}},{8{io_mask[0]}}} ;  
  assign io_out=wmask&(io_cmd==5'h8 ? (io_lhs&adder_out_mask)+(io_rhs&adder_out_mask):logic_and|logic_xor ? (logic_and ? io_lhs&io_rhs:64'h0)|(logic_xor ? io_lhs^io_rhs:64'h0):((io_mask[4] ? (io_lhs[63]==io_rhs[63] ? io_lhs[63:32]<io_rhs[63:32]|io_lhs[63:32]==io_rhs[63:32]&io_lhs[31:0]<io_rhs[31:0]:io_cmd[1] ? io_rhs[63]:io_lhs[63]):io_lhs[31]==io_rhs[31] ? io_lhs[31:0]<io_rhs[31:0]:io_cmd[1] ? io_rhs[31]:io_lhs[31]) ? io_cmd==5'hC|io_cmd==5'hE:io_cmd==5'hD|io_cmd==5'hF) ? io_lhs:io_rhs)|~wmask&io_lhs; 
endmodule
 
module tag_array_0_64x22 (
  input [5:0] RW0_addr,
  input RW0_en,
  input RW0_clk,
  input RW0_wmode,
  input [21:0] RW0_wdata,
  output [21:0] RW0_rdata) ; 
   reg [21:0] Memory[0:63] ;  
   reg [5:0] _RW0_raddr_d0 ;  
   reg _RW0_ren_d0 ;  
   reg _RW0_rmode_d0 ;  
  always @( posedge RW0_clk)
       begin 
         _RW0_raddr_d0 <=RW0_addr;
         _RW0_ren_d0 <=RW0_en;
         _RW0_rmode_d0 <=RW0_wmode;
         if (RW0_en&RW0_wmode&1'h1)
            Memory [RW0_addr]<=RW0_wdata;
       end
  
  assign RW0_rdata=_RW0_ren_d0&~_RW0_rmode_d0 ? Memory[_RW0_raddr_d0]:22'bx; 
endmodule
 
module DCache (
  input clock,
  input reset,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [1:0] auto_out_b_bits_param,
  input [3:0] auto_out_b_bits_size,
  input auto_out_b_bits_source,
  input [31:0] auto_out_b_bits_address,
  input auto_out_c_ready,
  output auto_out_c_valid,
  output [2:0] auto_out_c_bits_opcode,
  output [2:0] auto_out_c_bits_param,
  output [3:0] auto_out_c_bits_size,
  output auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_e_ready,
  output auto_out_e_valid,
  output [1:0] auto_out_e_bits_sink,
  output io_cpu_req_ready,
  input io_cpu_req_valid,
  input [33:0] io_cpu_req_bits_addr,
  input [5:0] io_cpu_req_bits_tag,
  input [4:0] io_cpu_req_bits_cmd,
  input [1:0] io_cpu_req_bits_size,
  input io_cpu_req_bits_signed,
  input io_cpu_req_bits_dv,
  input io_cpu_s1_kill,
  input [63:0] io_cpu_s1_data_data,
  input [7:0] io_cpu_s1_data_mask,
  output io_cpu_s2_nack,
  output io_cpu_resp_valid,
  output [33:0] io_cpu_resp_bits_addr,
  output [5:0] io_cpu_resp_bits_tag,
  output [4:0] io_cpu_resp_bits_cmd,
  output [1:0] io_cpu_resp_bits_size,
  output io_cpu_resp_bits_signed,
  output [1:0] io_cpu_resp_bits_dprv,
  output io_cpu_resp_bits_dv,
  output [63:0] io_cpu_resp_bits_data,
  output [7:0] io_cpu_resp_bits_mask,
  output io_cpu_resp_bits_replay,
  output io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output [63:0] io_cpu_resp_bits_data_raw,
  output [63:0] io_cpu_resp_bits_store_data,
  output io_cpu_replay_next,
  output io_cpu_s2_xcpt_ma_ld,
  output io_cpu_s2_xcpt_ma_st,
  output io_cpu_s2_xcpt_pf_ld,
  output io_cpu_s2_xcpt_pf_st,
  output io_cpu_s2_xcpt_ae_ld,
  output io_cpu_s2_xcpt_ae_st,
  output io_cpu_ordered,
  output io_cpu_perf_release,
  output io_cpu_perf_grant,
  output io_ptw_req_bits_bits_need_gpa,
  output io_ptw_req_bits_bits_stage2,
  input io_ptw_status_debug,
  input io_ptw_pmp_cfg_l_0,
  input io_ptw_pmp_cfg_l_1,
  input io_ptw_pmp_cfg_l_2,
  input io_ptw_pmp_cfg_l_3,
  input io_ptw_pmp_cfg_l_4,
  input io_ptw_pmp_cfg_l_5,
  input io_ptw_pmp_cfg_l_6,
  input io_ptw_pmp_cfg_l_7,
  input [1:0] io_ptw_pmp_cfg_a_0,
  input [1:0] io_ptw_pmp_cfg_a_1,
  input [1:0] io_ptw_pmp_cfg_a_2,
  input [1:0] io_ptw_pmp_cfg_a_3,
  input [1:0] io_ptw_pmp_cfg_a_4,
  input [1:0] io_ptw_pmp_cfg_a_5,
  input [1:0] io_ptw_pmp_cfg_a_6,
  input [1:0] io_ptw_pmp_cfg_a_7,
  input io_ptw_pmp_cfg_w_0,
  input io_ptw_pmp_cfg_w_1,
  input io_ptw_pmp_cfg_w_2,
  input io_ptw_pmp_cfg_w_3,
  input io_ptw_pmp_cfg_w_4,
  input io_ptw_pmp_cfg_w_5,
  input io_ptw_pmp_cfg_w_6,
  input io_ptw_pmp_cfg_w_7,
  input io_ptw_pmp_cfg_r_0,
  input io_ptw_pmp_cfg_r_1,
  input io_ptw_pmp_cfg_r_2,
  input io_ptw_pmp_cfg_r_3,
  input io_ptw_pmp_cfg_r_4,
  input io_ptw_pmp_cfg_r_5,
  input io_ptw_pmp_cfg_r_6,
  input io_ptw_pmp_cfg_r_7,
  input [29:0] io_ptw_pmp_addr_0,
  input [29:0] io_ptw_pmp_addr_1,
  input [29:0] io_ptw_pmp_addr_2,
  input [29:0] io_ptw_pmp_addr_3,
  input [29:0] io_ptw_pmp_addr_4,
  input [29:0] io_ptw_pmp_addr_5,
  input [29:0] io_ptw_pmp_addr_6,
  input [29:0] io_ptw_pmp_addr_7,
  input [31:0] io_ptw_pmp_mask_0,
  input [31:0] io_ptw_pmp_mask_1,
  input [31:0] io_ptw_pmp_mask_2,
  input [31:0] io_ptw_pmp_mask_3,
  input [31:0] io_ptw_pmp_mask_4,
  input [31:0] io_ptw_pmp_mask_5,
  input [31:0] io_ptw_pmp_mask_6,
  input [31:0] io_ptw_pmp_mask_7) ; 
   wire io_cpu_s2_xcpt_ma_st_0 ;  
   wire io_cpu_s2_xcpt_ma_ld_0 ;  
   wire io_cpu_s2_xcpt_ae_st_0 ;  
   wire io_cpu_s2_xcpt_ae_ld_0 ;  
   wire io_cpu_s2_xcpt_pf_st_0 ;  
   wire io_cpu_s2_xcpt_pf_ld_0 ;  
   wire [21:0] metaArb_io_in_bits_data_7 ;  
   wire metaArb_io_in_valid_4 ;  
   wire [11:0] dataArb_io_in_bits_addr_2 ;  
   wire dataArb_io_in_valid_2 ;  
   wire [3:0] nodeOut_c_bits_size ;  
   wire [2:0] nodeOut_c_bits_opcode ;  
   wire nodeOut_c_valid ;  
   wire [5:0] metaArb_io_in_bits_idx_6 ;  
   wire metaArb_io_in_valid_6 ;  
   wire s1_nack ;  
   wire dataArb_io_in_bits_write_1 ;  
   wire dataArb_io_in_valid_1 ;  
   wire nodeOut_d_ready ;  
   wire [21:0] metaArb_io_in_bits_data_3 ;  
   wire metaArb_io_in_valid_3 ;  
   wire [11:0] dataArb_io_in_bits_addr_1 ;  
   wire [7:0] dataArb_io_in_bits_eccMask_0 ;  
   wire [63:0] dataArb_io_in_bits_wdata_0 ;  
   wire [11:0] _dataArb_io_in_0_bits_wordMask_wordMask_T ;  
   wire dataArb_io_in_valid_0 ;  
   wire pstore_drain ;  
   wire [21:0] metaArb_io_in_bits_data_2 ;  
   wire [5:0] metaArb_io_in_bits_idx_3 ;  
   wire [5:0] metaArb_io_in_bits_idx_4 ;  
   wire metaArb_io_in_valid_2 ;  
   reg [33:0] s2_req_addr ;  
   wire readEnable ;  
   wire writeEnable ;  
   wire [5:0] metaArb_io_in_bits_idx_7 ;  
   wire [11:0] dataArb_io_in_bits_addr_3 ;  
   wire dataArb_io_in_valid_3 ;  
   reg [5:0] flushCounter ;  
   reg resetting ;  
   reg [33:0] s1_tlb_req_vaddr ;  
   wire [63:0] _amoalus_0_io_out ;  
   wire [63:0] _data_io_resp_0 ;  
   wire [21:0] _tag_array_0_ext_RW0_rdata ;  
   wire _tlb_pmp_io_r ;  
   wire _tlb_pmp_io_w ;  
   wire _GEN=metaArb_io_in_valid_2|metaArb_io_in_valid_3 ;  
   wire metaArb_io_out_bits_write=resetting|metaArb_io_in_valid_2|metaArb_io_in_valid_3|metaArb_io_in_valid_4 ;  
   wire metaArb__grant_T_2=resetting|metaArb_io_in_valid_2|metaArb_io_in_valid_3 ;  
   wire metaArb__grant_T_3=metaArb__grant_T_2|metaArb_io_in_valid_4 ;  
   wire metaArb__grant_T_5=metaArb__grant_T_3|metaArb_io_in_valid_6 ;  
   wire metaArb_io_out_valid=metaArb__grant_T_5|io_cpu_req_valid ;  
   wire dataArb__grant_T=dataArb_io_in_valid_0|dataArb_io_in_valid_1 ;  
   wire dataArb__grant_T_1=dataArb__grant_T|dataArb_io_in_valid_2 ;  
   wire dataArb_io_out_valid=dataArb__grant_T_1|dataArb_io_in_valid_3 ;  
   reg s1_valid ;  
   reg s1_probe ;  
   reg [1:0] probe_bits_param ;  
   reg [3:0] probe_bits_size ;  
   reg probe_bits_source ;  
   reg [31:0] probe_bits_address ;  
   wire s1_valid_masked=s1_valid&~io_cpu_s1_kill ;  
   reg [33:0] s1_vaddr ;  
   reg [5:0] s1_req_tag ;  
   reg [4:0] s1_req_cmd ;  
   reg [1:0] s1_req_size ;  
   reg s1_req_signed ;  
   reg [1:0] s1_req_dprv ;  
   reg s1_req_dv ;  
   reg [1:0] s1_tlb_req_size ;  
   reg [4:0] s1_tlb_req_cmd ;  
   reg [1:0] s1_tlb_req_prv ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_1=s1_req_cmd==5'h0 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_2=s1_req_cmd==5'h10 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_3=s1_req_cmd==5'h6 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_29=s1_req_cmd==5'h7 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_31=s1_req_cmd==5'h4 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_32=s1_req_cmd==5'h9 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_33=s1_req_cmd==5'hA ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_34=s1_req_cmd==5'hB ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_38=s1_req_cmd==5'h8 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_39=s1_req_cmd==5'hC ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_40=s1_req_cmd==5'hD ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_41=s1_req_cmd==5'hE ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_42=s1_req_cmd==5'hF ;  
   wire s1_read=_io_cpu_perf_canAcceptLoadThenLoad_T_1|_io_cpu_perf_canAcceptLoadThenLoad_T_2|_io_cpu_perf_canAcceptLoadThenLoad_T_3|_io_cpu_perf_canAcceptLoadThenLoad_T_29|_io_cpu_perf_canAcceptLoadThenLoad_T_31|_io_cpu_perf_canAcceptLoadThenLoad_T_32|_io_cpu_perf_canAcceptLoadThenLoad_T_33|_io_cpu_perf_canAcceptLoadThenLoad_T_34|_io_cpu_perf_canAcceptLoadThenLoad_T_38|_io_cpu_perf_canAcceptLoadThenLoad_T_39|_io_cpu_perf_canAcceptLoadThenLoad_T_40|_io_cpu_perf_canAcceptLoadThenLoad_T_41|_io_cpu_perf_canAcceptLoadThenLoad_T_42 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_26=s1_req_cmd==5'h1 ;  
   wire _io_cpu_perf_canAcceptLoadThenLoad_T_51=s1_req_cmd==5'h11 ;  
   wire s1_write=_io_cpu_perf_canAcceptLoadThenLoad_T_26|_io_cpu_perf_canAcceptLoadThenLoad_T_51|_io_cpu_perf_canAcceptLoadThenLoad_T_29|_io_cpu_perf_canAcceptLoadThenLoad_T_31|_io_cpu_perf_canAcceptLoadThenLoad_T_32|_io_cpu_perf_canAcceptLoadThenLoad_T_33|_io_cpu_perf_canAcceptLoadThenLoad_T_34|_io_cpu_perf_canAcceptLoadThenLoad_T_38|_io_cpu_perf_canAcceptLoadThenLoad_T_39|_io_cpu_perf_canAcceptLoadThenLoad_T_40|_io_cpu_perf_canAcceptLoadThenLoad_T_41|_io_cpu_perf_canAcceptLoadThenLoad_T_42 ;  
   reg s1_flush_valid ;  
   reg cached_grant_wait ;  
   reg release_ack_wait ;  
   reg [31:0] release_ack_addr ;  
   reg [3:0] release_state ;  
   wire _canAcceptCachedGrant_T=release_state==4'h1 ;  
   wire _inWriteback_T_1=release_state==4'h2 ;  
   wire inWriteback=_canAcceptCachedGrant_T|_inWriteback_T_1 ;  
   wire _io_cpu_req_ready_T_4=release_state==4'h0&~cached_grant_wait&~s1_nack ;  
   reg uncachedInFlight_0 ;  
   reg [33:0] uncachedReqs_addr_0 ;  
   reg [5:0] uncachedReqs_tag_0 ;  
   reg [1:0] uncachedReqs_size_0 ;  
   reg uncachedReqs_signed_0 ;  
   wire _pstore_drain_opportunistic_T=io_cpu_req_bits_cmd==5'h0 ;  
   wire _pstore_drain_opportunistic_T_1=io_cpu_req_bits_cmd==5'h10 ;  
   wire _pstore_drain_opportunistic_T_2=io_cpu_req_bits_cmd==5'h6 ;  
   wire _pstore_drain_opportunistic_T_28=io_cpu_req_bits_cmd==5'h7 ;  
   wire _pstore_drain_opportunistic_T_30=io_cpu_req_bits_cmd==5'h4 ;  
   wire _pstore_drain_opportunistic_T_31=io_cpu_req_bits_cmd==5'h9 ;  
   wire _pstore_drain_opportunistic_T_32=io_cpu_req_bits_cmd==5'hA ;  
   wire _pstore_drain_opportunistic_T_33=io_cpu_req_bits_cmd==5'hB ;  
   wire _pstore_drain_opportunistic_T_37=io_cpu_req_bits_cmd==5'h8 ;  
   wire _pstore_drain_opportunistic_T_38=io_cpu_req_bits_cmd==5'hC ;  
   wire _pstore_drain_opportunistic_T_39=io_cpu_req_bits_cmd==5'hD ;  
   wire _pstore_drain_opportunistic_T_40=io_cpu_req_bits_cmd==5'hE ;  
   wire _pstore_drain_opportunistic_T_41=io_cpu_req_bits_cmd==5'hF ;  
   wire _pstore_drain_opportunistic_T_25=io_cpu_req_bits_cmd==5'h1 ;  
   wire _pstore_drain_opportunistic_res_T_1=io_cpu_req_bits_cmd==5'h3 ;  
   wire _dataArb_io_in_3_valid_res_T_2=_pstore_drain_opportunistic_T_25|_pstore_drain_opportunistic_res_T_1 ;  
   wire _pstore_drain_opportunistic_T_50=io_cpu_req_bits_cmd==5'h11 ;  
  assign dataArb_io_in_valid_3=io_cpu_req_valid&~_dataArb_io_in_3_valid_res_T_2; 
  assign dataArb_io_in_bits_addr_3=io_cpu_req_bits_addr[11:0]; 
   wire _GEN_0=dataArb__grant_T_1&(_pstore_drain_opportunistic_T|_pstore_drain_opportunistic_T_1|_pstore_drain_opportunistic_T_2|_pstore_drain_opportunistic_T_28|_pstore_drain_opportunistic_T_30|_pstore_drain_opportunistic_T_31|_pstore_drain_opportunistic_T_32|_pstore_drain_opportunistic_T_33|_pstore_drain_opportunistic_T_37|_pstore_drain_opportunistic_T_38|_pstore_drain_opportunistic_T_39|_pstore_drain_opportunistic_T_40|_pstore_drain_opportunistic_T_41) ;  
   reg s1_did_read ;  
  assign metaArb_io_in_bits_idx_7=io_cpu_req_bits_addr[11:6]; 
  assign writeEnable=metaArb_io_out_valid&metaArb_io_out_bits_write; 
  assign readEnable=metaArb_io_out_valid&~metaArb_io_out_bits_write; 
   wire [1:0] _s1_mask_xwr_T={s1_vaddr[0]|(|s1_req_size),~(s1_vaddr[0])} ;  
   wire [3:0] _s1_mask_xwr_T_1={(s1_vaddr[1] ? _s1_mask_xwr_T:2'h0)|{2{s1_req_size[1]}},s1_vaddr[1] ? 2'h0:_s1_mask_xwr_T} ;  
   wire [7:0] s1_mask_xwr={(s1_vaddr[2] ? _s1_mask_xwr_T_1:4'h0)|{4{&s1_req_size}},s1_vaddr[2] ? 4'h0:_s1_mask_xwr_T_1} ;  
   reg s2_valid ;  
   wire s2_valid_no_xcpt=s2_valid&{io_cpu_s2_xcpt_ma_ld_0,io_cpu_s2_xcpt_ma_st_0,io_cpu_s2_xcpt_pf_ld_0,io_cpu_s2_xcpt_pf_st_0,io_cpu_s2_xcpt_ae_ld_0,io_cpu_s2_xcpt_ae_st_0}==6'h0 ;  
   reg s2_probe ;  
   wire releaseInFlight=s1_probe|s2_probe|(|release_state) ;  
   reg s2_not_nacked_in_s1 ;  
   wire s2_valid_masked=s2_valid_no_xcpt&s2_not_nacked_in_s1 ;  
   reg [5:0] s2_req_tag ;  
   reg [4:0] s2_req_cmd ;  
   reg [1:0] s2_req_size ;  
   reg s2_req_signed ;  
   reg [1:0] s2_req_dprv ;  
   reg s2_req_dv ;  
   reg s2_tlb_xcpt_pf_ld ;  
   reg s2_tlb_xcpt_pf_st ;  
   reg s2_tlb_xcpt_ae_ld ;  
   reg s2_tlb_xcpt_ae_st ;  
   reg s2_tlb_xcpt_ma_ld ;  
   reg s2_tlb_xcpt_ma_st ;  
   reg s2_pma_cacheable ;  
   reg [33:0] s2_uncached_resp_addr ;  
   reg [33:0] s2_vaddr_r ;  
   wire s2_lr=s2_req_cmd==5'h6 ;  
   wire s2_sc=s2_req_cmd==5'h7 ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_28=s2_req_cmd==5'h4 ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_29=s2_req_cmd==5'h9 ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_30=s2_req_cmd==5'hA ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_31=s2_req_cmd==5'hB ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_35=s2_req_cmd==5'h8 ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_36=s2_req_cmd==5'hC ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_37=s2_req_cmd==5'hD ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_38=s2_req_cmd==5'hE ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_39=s2_req_cmd==5'hF ;  
   wire s2_read=s2_req_cmd==5'h0|s2_req_cmd==5'h10|s2_lr|s2_sc|_metaArb_io_in_3_bits_data_c_cat_T_28|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_39 ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_23=s2_req_cmd==5'h1 ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_24=s2_req_cmd==5'h11 ;  
   wire s2_write=_metaArb_io_in_3_bits_data_c_cat_T_23|_metaArb_io_in_3_bits_data_c_cat_T_24|s2_sc|_metaArb_io_in_3_bits_data_c_cat_T_28|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_39 ;  
   wire s2_readwrite=s2_read|s2_write ;  
   reg s2_flush_valid ;  
   reg [21:0] s2_meta_corrected_r ;  
   reg [63:0] s2_data ;  
   reg [1:0] s2_probe_state_state ;  
   reg [1:0] s2_hit_state_state ;  
   wire _metaArb_io_in_3_bits_data_c_cat_T_46=s2_req_cmd==5'h3 ;  
   wire [3:0] _GEN_1={_metaArb_io_in_3_bits_data_c_cat_T_23|_metaArb_io_in_3_bits_data_c_cat_T_24|s2_sc|_metaArb_io_in_3_bits_data_c_cat_T_28|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_39,_metaArb_io_in_3_bits_data_c_cat_T_23|_metaArb_io_in_3_bits_data_c_cat_T_24|s2_sc|_metaArb_io_in_3_bits_data_c_cat_T_28|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_39|_metaArb_io_in_3_bits_data_c_cat_T_46|s2_lr,s2_hit_state_state} ;  
   wire s2_hit=_GEN_1==4'h3|_GEN_1==4'h2|_GEN_1==4'h1|_GEN_1==4'h7|_GEN_1==4'h6|(&_GEN_1)|_GEN_1==4'hE ;  
   reg [1:0] casez_tmp ;  
   wire [1:0] _GEN_2={1'h0,_GEN_1==4'hC} ;  
  always @(*)
       begin 
         casez (_GEN_1)
          4 'b0000:
             casez_tmp =2'h0;
          4 'b0001:
             casez_tmp =2'h1;
          4 'b0010:
             casez_tmp =2'h2;
          4 'b0011:
             casez_tmp =2'h3;
          4 'b0100:
             casez_tmp =2'h1;
          4 'b0101:
             casez_tmp =2'h2;
          4 'b0110:
             casez_tmp =2'h2;
          4 'b0111:
             casez_tmp =2'h3;
          4 'b1000:
             casez_tmp =_GEN_2;
          4 'b1001:
             casez_tmp =_GEN_2;
          4 'b1010:
             casez_tmp =_GEN_2;
          4 'b1011:
             casez_tmp =_GEN_2;
          4 'b1100:
             casez_tmp =_GEN_2;
          4 'b1101:
             casez_tmp =2'h2;
          4 'b1110:
             casez_tmp =2'h3;
          default :
             casez_tmp =2'h3;
         endcase 
       end
  
   wire s2_valid_hit_maybe_flush_pre_data_ecc_and_waw=s2_valid_masked&s2_hit ;  
   wire s2_valid_hit_pre_data_ecc_and_waw=s2_valid_hit_maybe_flush_pre_data_ecc_and_waw&s2_readwrite ;  
   wire s2_valid_flush_line=s2_valid_hit_maybe_flush_pre_data_ecc_and_waw&s2_req_cmd==5'h5&s2_req_size[0] ;  
   wire s2_valid_miss=s2_valid_masked&s2_readwrite&~s2_hit ;  
   wire s2_valid_cached_miss=s2_valid_miss&s2_pma_cacheable&~uncachedInFlight_0 ;  
   wire s2_want_victimize=s2_valid_cached_miss|s2_valid_flush_line|s2_flush_valid ;  
   wire s2_valid_uncached_pending=s2_valid_miss&~s2_pma_cacheable&~uncachedInFlight_0 ;  
   wire [1:0] s2_victim_state_state=(|s2_hit_state_state) ? s2_hit_state_state:s2_meta_corrected_r[21:20] ;  
   wire [3:0] _GEN_3={probe_bits_param,s2_probe_state_state} ;  
   wire _GEN_4=_GEN_3==4'hB ;  
   wire _GEN_5=_GEN_3==4'h4 ;  
   wire _GEN_6=_GEN_3==4'h5 ;  
   wire _GEN_7=_GEN_3==4'h6 ;  
   wire _GEN_8=_GEN_3==4'h7 ;  
   wire _GEN_9=_GEN_3==4'h0 ;  
   wire _GEN_10=_GEN_3==4'h1 ;  
   wire _GEN_11=_GEN_3==4'h2 ;  
   wire _GEN_12=_GEN_3==4'h3 ;  
   wire s2_prb_ack_data=_GEN_12|~(_GEN_11|_GEN_10|_GEN_9)&(_GEN_8|~(_GEN_7|_GEN_6|_GEN_5)&_GEN_4) ;  
   wire _GEN_13=_GEN_12|_GEN_11 ;  
   wire s2_victim_dirty=&s2_victim_state_state ;  
   wire io_cpu_s2_nack_0=s2_valid_no_xcpt&~(s2_valid_uncached_pending&auto_out_a_ready)&~(s2_valid_masked&s2_req_cmd==5'h17)&~s2_valid_hit_pre_data_ecc_and_waw ;  
  assign metaArb_io_in_valid_2=s2_valid_hit_pre_data_ecc_and_waw&s2_hit_state_state!=casez_tmp; 
   wire _GEN_14=io_cpu_s2_nack_0|metaArb_io_in_valid_2 ;  
  assign metaArb_io_in_bits_idx_4=probe_bits_address[11:6]; 
  assign metaArb_io_in_bits_idx_3=s2_req_addr[11:6]; 
  assign metaArb_io_in_bits_data_2={casez_tmp,s2_req_addr[31:12]}; 
   reg [6:0] lrscCount ;  
   reg [27:0] lrscAddr ;  
   wire s2_sc_fail=s2_sc&~((|(lrscCount[6:2]))&lrscAddr==s2_req_addr[33:6]) ;  
   reg [4:0] pstore1_cmd ;  
   reg [33:0] pstore1_addr ;  
   reg [63:0] pstore1_data ;  
   reg [7:0] pstore1_mask ;  
   reg pstore1_rmw ;  
   wire _pstore1_held_T=s2_valid_hit_pre_data_ecc_and_waw&s2_write ;  
   reg pstore2_valid ;  
   wire _pstore_drain_opportunistic_res_T_2=_pstore_drain_opportunistic_T_25|_pstore_drain_opportunistic_res_T_1 ;  
   reg pstore_drain_on_miss_REG ;  
   reg pstore1_held ;  
   wire pstore1_valid_likely=s2_valid&s2_write|pstore1_held ;  
   wire pstore1_valid=_pstore1_held_T&~s2_sc_fail|pstore1_held ;  
   wire pstore_drain_structural=pstore1_valid_likely&pstore2_valid&(s1_valid&s1_write|pstore1_rmw) ;  
   wire _dataArb_io_in_0_valid_T_4=s2_valid_hit_pre_data_ecc_and_waw&s2_write ;  
   wire _dataArb_io_in_0_valid_T_9=~(io_cpu_req_valid&~_pstore_drain_opportunistic_res_T_2)|releaseInFlight|pstore_drain_on_miss_REG ;  
  assign pstore_drain=pstore_drain_structural|((_dataArb_io_in_0_valid_T_4|pstore1_held)&~pstore1_rmw|pstore2_valid)&_dataArb_io_in_0_valid_T_9; 
   reg [33:0] pstore2_addr ;  
   reg [7:0] pstore2_storegen_data_r ;  
   reg [7:0] pstore2_storegen_data_r_1 ;  
   reg [7:0] pstore2_storegen_data_r_2 ;  
   reg [7:0] pstore2_storegen_data_r_3 ;  
   reg [7:0] pstore2_storegen_data_r_4 ;  
   reg [7:0] pstore2_storegen_data_r_5 ;  
   reg [7:0] pstore2_storegen_data_r_6 ;  
   reg [7:0] pstore2_storegen_data_r_7 ;  
   reg [7:0] pstore2_storegen_mask ;  
  assign dataArb_io_in_valid_0=pstore_drain_structural|((_dataArb_io_in_0_valid_T_4|pstore1_held)&~pstore1_rmw|pstore2_valid)&_dataArb_io_in_0_valid_T_9; 
  assign _dataArb_io_in_0_bits_wordMask_wordMask_T=pstore2_valid ? pstore2_addr[11:0]:pstore1_addr[11:0]; 
  assign dataArb_io_in_bits_wdata_0=pstore2_valid ? {pstore2_storegen_data_r_7,pstore2_storegen_data_r_6,pstore2_storegen_data_r_5,pstore2_storegen_data_r_4,pstore2_storegen_data_r_3,pstore2_storegen_data_r_2,pstore2_storegen_data_r_1,pstore2_storegen_data_r}:pstore1_data; 
  assign dataArb_io_in_bits_eccMask_0=pstore2_valid ? pstore2_storegen_mask:pstore1_mask; 
   wire _GEN_15=s1_valid&s1_read&(pstore1_valid_likely&pstore1_addr[11:3]==s1_vaddr[11:3]&(s1_write ? (|(pstore1_mask&s1_mask_xwr)):(|(pstore1_mask&s1_mask_xwr)))|pstore2_valid&pstore2_addr[11:3]==s1_vaddr[11:3]&(s1_write ? (|(pstore2_storegen_mask&s1_mask_xwr)):(|(pstore2_storegen_mask&s1_mask_xwr)))) ;  
   wire get_a_mask_size=s2_req_size==2'h2 ;  
   wire get_a_mask_acc=(&s2_req_size)|get_a_mask_size&~(s2_req_addr[2]) ;  
   wire get_a_mask_acc_1=(&s2_req_size)|get_a_mask_size&s2_req_addr[2] ;  
   wire get_a_mask_size_1=s2_req_size==2'h1 ;  
   wire get_a_mask_eq_2=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire get_a_mask_acc_2=get_a_mask_acc|get_a_mask_size_1&get_a_mask_eq_2 ;  
   wire get_a_mask_eq_3=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire get_a_mask_acc_3=get_a_mask_acc|get_a_mask_size_1&get_a_mask_eq_3 ;  
   wire get_a_mask_eq_4=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire get_a_mask_acc_4=get_a_mask_acc_1|get_a_mask_size_1&get_a_mask_eq_4 ;  
   wire get_a_mask_eq_5=s2_req_addr[2]&s2_req_addr[1] ;  
   wire get_a_mask_acc_5=get_a_mask_acc_1|get_a_mask_size_1&get_a_mask_eq_5 ;  
   wire put_a_mask_size=s2_req_size==2'h2 ;  
   wire put_a_mask_acc=(&s2_req_size)|put_a_mask_size&~(s2_req_addr[2]) ;  
   wire put_a_mask_acc_1=(&s2_req_size)|put_a_mask_size&s2_req_addr[2] ;  
   wire put_a_mask_size_1=s2_req_size==2'h1 ;  
   wire put_a_mask_eq_2=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire put_a_mask_acc_2=put_a_mask_acc|put_a_mask_size_1&put_a_mask_eq_2 ;  
   wire put_a_mask_eq_3=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire put_a_mask_acc_3=put_a_mask_acc|put_a_mask_size_1&put_a_mask_eq_3 ;  
   wire put_a_mask_eq_4=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire put_a_mask_acc_4=put_a_mask_acc_1|put_a_mask_size_1&put_a_mask_eq_4 ;  
   wire put_a_mask_eq_5=s2_req_addr[2]&s2_req_addr[1] ;  
   wire put_a_mask_acc_5=put_a_mask_acc_1|put_a_mask_size_1&put_a_mask_eq_5 ;  
   wire atomics_a_mask_size=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc=(&s2_req_size)|atomics_a_mask_size&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_1=(&s2_req_size)|atomics_a_mask_size&s2_req_addr[2] ;  
   wire atomics_a_mask_size_1=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_2=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_2=atomics_a_mask_acc|atomics_a_mask_size_1&atomics_a_mask_eq_2 ;  
   wire atomics_a_mask_eq_3=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_3=atomics_a_mask_acc|atomics_a_mask_size_1&atomics_a_mask_eq_3 ;  
   wire atomics_a_mask_eq_4=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_4=atomics_a_mask_acc_1|atomics_a_mask_size_1&atomics_a_mask_eq_4 ;  
   wire atomics_a_mask_eq_5=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_5=atomics_a_mask_acc_1|atomics_a_mask_size_1&atomics_a_mask_eq_5 ;  
   wire atomics_a_mask_size_3=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_14=(&s2_req_size)|atomics_a_mask_size_3&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_15=(&s2_req_size)|atomics_a_mask_size_3&s2_req_addr[2] ;  
   wire atomics_a_mask_size_4=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_16=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_16=atomics_a_mask_acc_14|atomics_a_mask_size_4&atomics_a_mask_eq_16 ;  
   wire atomics_a_mask_eq_17=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_17=atomics_a_mask_acc_14|atomics_a_mask_size_4&atomics_a_mask_eq_17 ;  
   wire atomics_a_mask_eq_18=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_18=atomics_a_mask_acc_15|atomics_a_mask_size_4&atomics_a_mask_eq_18 ;  
   wire atomics_a_mask_eq_19=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_19=atomics_a_mask_acc_15|atomics_a_mask_size_4&atomics_a_mask_eq_19 ;  
   wire atomics_a_mask_size_6=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_28=(&s2_req_size)|atomics_a_mask_size_6&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_29=(&s2_req_size)|atomics_a_mask_size_6&s2_req_addr[2] ;  
   wire atomics_a_mask_size_7=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_30=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_30=atomics_a_mask_acc_28|atomics_a_mask_size_7&atomics_a_mask_eq_30 ;  
   wire atomics_a_mask_eq_31=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_31=atomics_a_mask_acc_28|atomics_a_mask_size_7&atomics_a_mask_eq_31 ;  
   wire atomics_a_mask_eq_32=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_32=atomics_a_mask_acc_29|atomics_a_mask_size_7&atomics_a_mask_eq_32 ;  
   wire atomics_a_mask_eq_33=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_33=atomics_a_mask_acc_29|atomics_a_mask_size_7&atomics_a_mask_eq_33 ;  
   wire atomics_a_mask_size_9=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_42=(&s2_req_size)|atomics_a_mask_size_9&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_43=(&s2_req_size)|atomics_a_mask_size_9&s2_req_addr[2] ;  
   wire atomics_a_mask_size_10=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_44=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_44=atomics_a_mask_acc_42|atomics_a_mask_size_10&atomics_a_mask_eq_44 ;  
   wire atomics_a_mask_eq_45=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_45=atomics_a_mask_acc_42|atomics_a_mask_size_10&atomics_a_mask_eq_45 ;  
   wire atomics_a_mask_eq_46=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_46=atomics_a_mask_acc_43|atomics_a_mask_size_10&atomics_a_mask_eq_46 ;  
   wire atomics_a_mask_eq_47=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_47=atomics_a_mask_acc_43|atomics_a_mask_size_10&atomics_a_mask_eq_47 ;  
   wire atomics_a_mask_size_12=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_56=(&s2_req_size)|atomics_a_mask_size_12&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_57=(&s2_req_size)|atomics_a_mask_size_12&s2_req_addr[2] ;  
   wire atomics_a_mask_size_13=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_58=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_58=atomics_a_mask_acc_56|atomics_a_mask_size_13&atomics_a_mask_eq_58 ;  
   wire atomics_a_mask_eq_59=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_59=atomics_a_mask_acc_56|atomics_a_mask_size_13&atomics_a_mask_eq_59 ;  
   wire atomics_a_mask_eq_60=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_60=atomics_a_mask_acc_57|atomics_a_mask_size_13&atomics_a_mask_eq_60 ;  
   wire atomics_a_mask_eq_61=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_61=atomics_a_mask_acc_57|atomics_a_mask_size_13&atomics_a_mask_eq_61 ;  
   wire atomics_a_mask_size_15=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_70=(&s2_req_size)|atomics_a_mask_size_15&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_71=(&s2_req_size)|atomics_a_mask_size_15&s2_req_addr[2] ;  
   wire atomics_a_mask_size_16=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_72=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_72=atomics_a_mask_acc_70|atomics_a_mask_size_16&atomics_a_mask_eq_72 ;  
   wire atomics_a_mask_eq_73=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_73=atomics_a_mask_acc_70|atomics_a_mask_size_16&atomics_a_mask_eq_73 ;  
   wire atomics_a_mask_eq_74=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_74=atomics_a_mask_acc_71|atomics_a_mask_size_16&atomics_a_mask_eq_74 ;  
   wire atomics_a_mask_eq_75=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_75=atomics_a_mask_acc_71|atomics_a_mask_size_16&atomics_a_mask_eq_75 ;  
   wire atomics_a_mask_size_18=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_84=(&s2_req_size)|atomics_a_mask_size_18&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_85=(&s2_req_size)|atomics_a_mask_size_18&s2_req_addr[2] ;  
   wire atomics_a_mask_size_19=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_86=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_86=atomics_a_mask_acc_84|atomics_a_mask_size_19&atomics_a_mask_eq_86 ;  
   wire atomics_a_mask_eq_87=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_87=atomics_a_mask_acc_84|atomics_a_mask_size_19&atomics_a_mask_eq_87 ;  
   wire atomics_a_mask_eq_88=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_88=atomics_a_mask_acc_85|atomics_a_mask_size_19&atomics_a_mask_eq_88 ;  
   wire atomics_a_mask_eq_89=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_89=atomics_a_mask_acc_85|atomics_a_mask_size_19&atomics_a_mask_eq_89 ;  
   wire atomics_a_mask_size_21=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_98=(&s2_req_size)|atomics_a_mask_size_21&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_99=(&s2_req_size)|atomics_a_mask_size_21&s2_req_addr[2] ;  
   wire atomics_a_mask_size_22=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_100=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_100=atomics_a_mask_acc_98|atomics_a_mask_size_22&atomics_a_mask_eq_100 ;  
   wire atomics_a_mask_eq_101=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_101=atomics_a_mask_acc_98|atomics_a_mask_size_22&atomics_a_mask_eq_101 ;  
   wire atomics_a_mask_eq_102=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_102=atomics_a_mask_acc_99|atomics_a_mask_size_22&atomics_a_mask_eq_102 ;  
   wire atomics_a_mask_eq_103=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_103=atomics_a_mask_acc_99|atomics_a_mask_size_22&atomics_a_mask_eq_103 ;  
   wire atomics_a_mask_size_24=s2_req_size==2'h2 ;  
   wire atomics_a_mask_acc_112=(&s2_req_size)|atomics_a_mask_size_24&~(s2_req_addr[2]) ;  
   wire atomics_a_mask_acc_113=(&s2_req_size)|atomics_a_mask_size_24&s2_req_addr[2] ;  
   wire atomics_a_mask_size_25=s2_req_size==2'h1 ;  
   wire atomics_a_mask_eq_114=~(s2_req_addr[2])&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_114=atomics_a_mask_acc_112|atomics_a_mask_size_25&atomics_a_mask_eq_114 ;  
   wire atomics_a_mask_eq_115=~(s2_req_addr[2])&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_115=atomics_a_mask_acc_112|atomics_a_mask_size_25&atomics_a_mask_eq_115 ;  
   wire atomics_a_mask_eq_116=s2_req_addr[2]&~(s2_req_addr[1]) ;  
   wire atomics_a_mask_acc_116=atomics_a_mask_acc_113|atomics_a_mask_size_25&atomics_a_mask_eq_116 ;  
   wire atomics_a_mask_eq_117=s2_req_addr[2]&s2_req_addr[1] ;  
   wire atomics_a_mask_acc_117=atomics_a_mask_acc_113|atomics_a_mask_size_25&atomics_a_mask_eq_117 ;  
   wire [7:0] atomics_mask=_metaArb_io_in_3_bits_data_c_cat_T_39 ? {atomics_a_mask_acc_117|atomics_a_mask_eq_117&s2_req_addr[0],atomics_a_mask_acc_117|atomics_a_mask_eq_117&~(s2_req_addr[0]),atomics_a_mask_acc_116|atomics_a_mask_eq_116&s2_req_addr[0],atomics_a_mask_acc_116|atomics_a_mask_eq_116&~(s2_req_addr[0]),atomics_a_mask_acc_115|atomics_a_mask_eq_115&s2_req_addr[0],atomics_a_mask_acc_115|atomics_a_mask_eq_115&~(s2_req_addr[0]),atomics_a_mask_acc_114|atomics_a_mask_eq_114&s2_req_addr[0],atomics_a_mask_acc_114|atomics_a_mask_eq_114&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_38 ? {atomics_a_mask_acc_103|atomics_a_mask_eq_103&s2_req_addr[0],atomics_a_mask_acc_103|atomics_a_mask_eq_103&~(s2_req_addr[0]),atomics_a_mask_acc_102|atomics_a_mask_eq_102&s2_req_addr[0],atomics_a_mask_acc_102|atomics_a_mask_eq_102&~(s2_req_addr[0]),atomics_a_mask_acc_101|atomics_a_mask_eq_101&s2_req_addr[0],atomics_a_mask_acc_101|atomics_a_mask_eq_101&~(s2_req_addr[0]),atomics_a_mask_acc_100|atomics_a_mask_eq_100&s2_req_addr[0],atomics_a_mask_acc_100|atomics_a_mask_eq_100&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_37 ? {atomics_a_mask_acc_89|atomics_a_mask_eq_89&s2_req_addr[0],atomics_a_mask_acc_89|atomics_a_mask_eq_89&~(s2_req_addr[0]),atomics_a_mask_acc_88|atomics_a_mask_eq_88&s2_req_addr[0],atomics_a_mask_acc_88|atomics_a_mask_eq_88&~(s2_req_addr[0]),atomics_a_mask_acc_87|atomics_a_mask_eq_87&s2_req_addr[0],atomics_a_mask_acc_87|atomics_a_mask_eq_87&~(s2_req_addr[0]),atomics_a_mask_acc_86|atomics_a_mask_eq_86&s2_req_addr[0],atomics_a_mask_acc_86|atomics_a_mask_eq_86&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_36 ? {atomics_a_mask_acc_75|atomics_a_mask_eq_75&s2_req_addr[0],atomics_a_mask_acc_75|atomics_a_mask_eq_75&~(s2_req_addr[0]),atomics_a_mask_acc_74|atomics_a_mask_eq_74&s2_req_addr[0],atomics_a_mask_acc_74|atomics_a_mask_eq_74&~(s2_req_addr[0]),atomics_a_mask_acc_73|atomics_a_mask_eq_73&s2_req_addr[0],atomics_a_mask_acc_73|atomics_a_mask_eq_73&~(s2_req_addr[0]),atomics_a_mask_acc_72|atomics_a_mask_eq_72&s2_req_addr[0],atomics_a_mask_acc_72|atomics_a_mask_eq_72&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_35 ? {atomics_a_mask_acc_61|atomics_a_mask_eq_61&s2_req_addr[0],atomics_a_mask_acc_61|atomics_a_mask_eq_61&~(s2_req_addr[0]),atomics_a_mask_acc_60|atomics_a_mask_eq_60&s2_req_addr[0],atomics_a_mask_acc_60|atomics_a_mask_eq_60&~(s2_req_addr[0]),atomics_a_mask_acc_59|atomics_a_mask_eq_59&s2_req_addr[0],atomics_a_mask_acc_59|atomics_a_mask_eq_59&~(s2_req_addr[0]),atomics_a_mask_acc_58|atomics_a_mask_eq_58&s2_req_addr[0],atomics_a_mask_acc_58|atomics_a_mask_eq_58&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_31 ? {atomics_a_mask_acc_47|atomics_a_mask_eq_47&s2_req_addr[0],atomics_a_mask_acc_47|atomics_a_mask_eq_47&~(s2_req_addr[0]),atomics_a_mask_acc_46|atomics_a_mask_eq_46&s2_req_addr[0],atomics_a_mask_acc_46|atomics_a_mask_eq_46&~(s2_req_addr[0]),atomics_a_mask_acc_45|atomics_a_mask_eq_45&s2_req_addr[0],atomics_a_mask_acc_45|atomics_a_mask_eq_45&~(s2_req_addr[0]),atomics_a_mask_acc_44|atomics_a_mask_eq_44&s2_req_addr[0],atomics_a_mask_acc_44|atomics_a_mask_eq_44&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_30 ? {atomics_a_mask_acc_33|atomics_a_mask_eq_33&s2_req_addr[0],atomics_a_mask_acc_33|atomics_a_mask_eq_33&~(s2_req_addr[0]),atomics_a_mask_acc_32|atomics_a_mask_eq_32&s2_req_addr[0],atomics_a_mask_acc_32|atomics_a_mask_eq_32&~(s2_req_addr[0]),atomics_a_mask_acc_31|atomics_a_mask_eq_31&s2_req_addr[0],atomics_a_mask_acc_31|atomics_a_mask_eq_31&~(s2_req_addr[0]),atomics_a_mask_acc_30|atomics_a_mask_eq_30&s2_req_addr[0],atomics_a_mask_acc_30|atomics_a_mask_eq_30&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_29 ? {atomics_a_mask_acc_19|atomics_a_mask_eq_19&s2_req_addr[0],atomics_a_mask_acc_19|atomics_a_mask_eq_19&~(s2_req_addr[0]),atomics_a_mask_acc_18|atomics_a_mask_eq_18&s2_req_addr[0],atomics_a_mask_acc_18|atomics_a_mask_eq_18&~(s2_req_addr[0]),atomics_a_mask_acc_17|atomics_a_mask_eq_17&s2_req_addr[0],atomics_a_mask_acc_17|atomics_a_mask_eq_17&~(s2_req_addr[0]),atomics_a_mask_acc_16|atomics_a_mask_eq_16&s2_req_addr[0],atomics_a_mask_acc_16|atomics_a_mask_eq_16&~(s2_req_addr[0])}:_metaArb_io_in_3_bits_data_c_cat_T_28 ? {atomics_a_mask_acc_5|atomics_a_mask_eq_5&s2_req_addr[0],atomics_a_mask_acc_5|atomics_a_mask_eq_5&~(s2_req_addr[0]),atomics_a_mask_acc_4|atomics_a_mask_eq_4&s2_req_addr[0],atomics_a_mask_acc_4|atomics_a_mask_eq_4&~(s2_req_addr[0]),atomics_a_mask_acc_3|atomics_a_mask_eq_3&s2_req_addr[0],atomics_a_mask_acc_3|atomics_a_mask_eq_3&~(s2_req_addr[0]),atomics_a_mask_acc_2|atomics_a_mask_eq_2&s2_req_addr[0],atomics_a_mask_acc_2|atomics_a_mask_eq_2&~(s2_req_addr[0])}:8'h0 ;  
   wire tl_out_a_valid=s2_valid_uncached_pending|s2_valid_cached_miss&~(release_ack_wait&(s2_req_addr[20:6]^release_ack_addr[20:6])==15'h0)&~s2_victim_dirty ;  
   wire _GEN_16=~s2_write|_metaArb_io_in_3_bits_data_c_cat_T_24|~s2_read|_metaArb_io_in_3_bits_data_c_cat_T_39|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_28 ;  
   wire _io_errors_bus_valid_T=nodeOut_d_ready&auto_out_d_valid ;  
   wire [26:0] _beats1_decode_T_1=27'hFFF<<auto_out_d_bits_size ;  
   wire [8:0] beats1=auto_out_d_bits_opcode[0] ? ~(_beats1_decode_T_1[11:3]):9'h0 ;  
   reg [8:0] counter ;  
   wire [8:0] _counter1_T=counter-9'h1 ;  
   wire d_last=counter==9'h1|beats1==9'h0 ;  
   wire [8:0] count=beats1&~_counter1_T ;  
   wire grantIsUncachedData=auto_out_d_bits_opcode==3'h1 ;  
   wire grantIsUncached=grantIsUncachedData|auto_out_d_bits_opcode==3'h0|auto_out_d_bits_opcode==3'h2 ;  
   wire grantIsRefill=auto_out_d_bits_opcode==3'h5 ;  
   wire grantIsCached=auto_out_d_bits_opcode==3'h4|grantIsRefill ;  
   wire grantIsVoluntary=auto_out_d_bits_opcode==3'h6 ;  
   reg grantInProgress ;  
   reg [2:0] blockProbeAfterGrantCount ;  
   wire _metaArb_io_in_4_valid_T=release_state==4'h6 ;  
   wire _nodeOut_c_valid_T_1=release_state==4'h9 ;  
   wire _canAcceptCachedGrant_T_4=_canAcceptCachedGrant_T|_metaArb_io_in_4_valid_T|_nodeOut_c_valid_T_1 ;  
   wire _GEN_17=_io_errors_bus_valid_T&grantIsCached ;  
   wire _GEN_18=auto_out_d_bits_source&d_last ;  
   wire _GEN_19=~_io_errors_bus_valid_T|grantIsCached|~(grantIsUncached&grantIsUncachedData) ;  
   wire _GEN_20=grantIsRefill&dataArb_io_in_valid_0 ;  
   wire nodeOut_e_valid=~_GEN_20&auto_out_d_valid&~(|counter)&grantIsCached&~_canAcceptCachedGrant_T_4 ;  
  assign dataArb_io_in_bits_addr_1={s2_req_addr[11:6]|count[8:3],count[2:0],3'h0}; 
  assign metaArb_io_in_valid_3=grantIsCached&d_last&_io_errors_bus_valid_T&~auto_out_d_bits_denied; 
   wire [3:0] _metaArb_io_in_3_bits_data_T_1={_metaArb_io_in_3_bits_data_c_cat_T_23|_metaArb_io_in_3_bits_data_c_cat_T_24|s2_sc|_metaArb_io_in_3_bits_data_c_cat_T_28|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_39,_metaArb_io_in_3_bits_data_c_cat_T_23|_metaArb_io_in_3_bits_data_c_cat_T_24|s2_sc|_metaArb_io_in_3_bits_data_c_cat_T_28|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_39|_metaArb_io_in_3_bits_data_c_cat_T_46|s2_lr,auto_out_d_bits_param} ;  
  assign metaArb_io_in_bits_data_3={_metaArb_io_in_3_bits_data_T_1==4'hC ? 2'h3:_metaArb_io_in_3_bits_data_T_1==4'h4|_metaArb_io_in_3_bits_data_T_1==4'h0 ? 2'h2:{1'h0,_metaArb_io_in_3_bits_data_T_1==4'h1},s2_req_addr[31:12]}; 
   reg blockUncachedGrant ;  
   wire _GEN_21=grantIsUncachedData&(blockUncachedGrant|s1_valid) ;  
  assign nodeOut_d_ready=~(_GEN_21|_GEN_20)&(~grantIsCached|((|counter)|auto_out_e_ready)&~_canAcceptCachedGrant_T_4); 
   wire io_cpu_req_ready_0=_GEN_21 ? ~(auto_out_d_valid|metaArb__grant_T_5|_GEN_0)&_io_cpu_req_ready_T_4:~(metaArb__grant_T_5|_GEN_0)&_io_cpu_req_ready_T_4 ;  
   wire _GEN_22=_GEN_21&auto_out_d_valid ;  
  assign dataArb_io_in_valid_1=_GEN_22|auto_out_d_valid&grantIsRefill&~_canAcceptCachedGrant_T_4; 
  assign dataArb_io_in_bits_write_1=~_GEN_21|~auto_out_d_valid; 
   wire block_probe_for_core_progress=(|blockProbeAfterGrantCount)|(|(lrscCount[6:2])) ;  
   wire nodeOut_b_ready=~metaArb__grant_T_3&~(block_probe_for_core_progress|releaseInFlight|release_ack_wait&(auto_out_b_bits_address[20:6]^release_ack_addr[20:6])==15'h0|grantInProgress|s1_valid|s2_valid) ;  
   wire _io_cpu_perf_release_T=auto_out_c_ready&nodeOut_c_valid ;  
   wire [26:0] _GEN_23={23'h0,nodeOut_c_bits_size} ;  
   wire [26:0] _beats1_decode_T_5=27'hFFF<<_GEN_23 ;  
   wire [8:0] beats1_1=nodeOut_c_bits_opcode[0] ? ~(_beats1_decode_T_5[11:3]):9'h0 ;  
   reg [8:0] counter_1 ;  
   wire [8:0] _counter1_T_1=counter_1-9'h1 ;  
   wire c_first=counter_1==9'h0 ;  
   wire releaseDone=(counter_1==9'h1|beats1_1==9'h0)&_io_cpu_perf_release_T ;  
   reg s1_release_data_valid ;  
   reg s2_release_data_valid ;  
   wire releaseRejected=s2_release_data_valid&~_io_cpu_perf_release_T ;  
   wire [9:0] _releaseDataBeat_T_5={1'h0,beats1_1&~_counter1_T_1}+{8'h0,releaseRejected ? 2'h0:{1'h0,s1_release_data_valid}+{1'h0,s2_release_data_valid}} ;  
  assign s1_nack=s2_probe ? s2_prb_ack_data|(|s2_probe_state_state)|~releaseDone|_GEN_15|_GEN_14:_GEN_15|_GEN_14; 
   wire _GEN_24=release_state==4'h4 ;  
  assign metaArb_io_in_valid_6=_GEN_24|auto_out_b_valid&(~block_probe_for_core_progress|(|lrscCount)&~(|(lrscCount[6:2]))); 
  assign metaArb_io_in_bits_idx_6=_GEN_24 ? metaArb_io_in_bits_idx_4:auto_out_b_bits_address[11:6]; 
   wire _GEN_25=release_state==4'h5 ;  
   wire _GEN_26=release_state==4'h3 ;  
  assign nodeOut_c_valid=_GEN_26|_GEN_25|s2_probe&~s2_prb_ack_data|s2_release_data_valid&~(c_first&release_ack_wait); 
   wire _GEN_27=_canAcceptCachedGrant_T|_metaArb_io_in_4_valid_T|_nodeOut_c_valid_T_1 ;  
  assign nodeOut_c_bits_opcode=_GEN_27 ? {2'h3,~_nodeOut_c_valid_T_1}:{2'h2,_inWriteback_T_1}; 
  assign nodeOut_c_bits_size=_GEN_27 ? 4'h6:probe_bits_size; 
  assign dataArb_io_in_valid_2=inWriteback&_releaseDataBeat_T_5<10'h8; 
  assign dataArb_io_in_bits_addr_2={metaArb_io_in_bits_idx_4,_releaseDataBeat_T_5[2:0],3'h0}; 
  assign metaArb_io_in_valid_4=_metaArb_io_in_4_valid_T|release_state==4'h7; 
  assign metaArb_io_in_bits_data_7={_GEN_27 ? 2'h0:_GEN_13 ? 2'h2:_GEN_10 ? 2'h1:_GEN_9 ? 2'h0:{1'h0,_GEN_8|_GEN_7|_GEN_6},probe_bits_address[31:12]}; 
   reg io_cpu_s2_xcpt_REG ;  
  assign io_cpu_s2_xcpt_pf_ld_0=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_pf_ld; 
  assign io_cpu_s2_xcpt_pf_st_0=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_pf_st; 
  assign io_cpu_s2_xcpt_ae_ld_0=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ae_ld; 
  assign io_cpu_s2_xcpt_ae_st_0=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ae_st; 
  assign io_cpu_s2_xcpt_ma_ld_0=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ma_ld; 
  assign io_cpu_s2_xcpt_ma_st_0=io_cpu_s2_xcpt_REG&s2_tlb_xcpt_ma_st; 
   reg doUncachedResp ;  
   wire io_cpu_replay_next_0=_io_errors_bus_valid_T&grantIsUncachedData ;  
   wire _GEN_28=_io_errors_bus_valid_T&~grantIsCached ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~(_pstore_drain_opportunistic_T|_pstore_drain_opportunistic_T_1|_pstore_drain_opportunistic_T_2|_pstore_drain_opportunistic_T_28|_pstore_drain_opportunistic_T_30|_pstore_drain_opportunistic_T_31|_pstore_drain_opportunistic_T_32|_pstore_drain_opportunistic_T_33|_pstore_drain_opportunistic_T_37|_pstore_drain_opportunistic_T_38|_pstore_drain_opportunistic_T_39|_pstore_drain_opportunistic_T_40|_pstore_drain_opportunistic_T_41|(_pstore_drain_opportunistic_T_25|_pstore_drain_opportunistic_T_50|_pstore_drain_opportunistic_T_28|_pstore_drain_opportunistic_T_30|_pstore_drain_opportunistic_T_31|_pstore_drain_opportunistic_T_32|_pstore_drain_opportunistic_T_33|_pstore_drain_opportunistic_T_37|_pstore_drain_opportunistic_T_38|_pstore_drain_opportunistic_T_39|_pstore_drain_opportunistic_T_40|_pstore_drain_opportunistic_T_41)&_pstore_drain_opportunistic_T_50)|~_dataArb_io_in_3_valid_res_T_2))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
              if (1)$display("");
            end 
         if (~reset&~(~(s1_valid_masked&_io_cpu_perf_canAcceptLoadThenLoad_T_51)|(&(s1_mask_xwr|~io_cpu_s1_data_mask))))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:306 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n");
              if (1)$display("");
            end 
         if (~reset&~(~(_pstore_drain_opportunistic_T|_pstore_drain_opportunistic_T_1|_pstore_drain_opportunistic_T_2|_pstore_drain_opportunistic_T_28|_pstore_drain_opportunistic_T_30|_pstore_drain_opportunistic_T_31|_pstore_drain_opportunistic_T_32|_pstore_drain_opportunistic_T_33|_pstore_drain_opportunistic_T_37|_pstore_drain_opportunistic_T_38|_pstore_drain_opportunistic_T_39|_pstore_drain_opportunistic_T_40|_pstore_drain_opportunistic_T_41|(_pstore_drain_opportunistic_T_25|_pstore_drain_opportunistic_T_50|_pstore_drain_opportunistic_T_28|_pstore_drain_opportunistic_T_30|_pstore_drain_opportunistic_T_31|_pstore_drain_opportunistic_T_32|_pstore_drain_opportunistic_T_33|_pstore_drain_opportunistic_T_37|_pstore_drain_opportunistic_T_38|_pstore_drain_opportunistic_T_39|_pstore_drain_opportunistic_T_40|_pstore_drain_opportunistic_T_41)&_pstore_drain_opportunistic_T_50)|~_pstore_drain_opportunistic_res_T_2))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
              if (1)$display("");
            end 
         if (~reset&~(pstore1_rmw|(_dataArb_io_in_0_valid_T_4|pstore1_held)==pstore1_valid))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:487 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~reset&~cached_grant_wait)
            begin 
              if (1)$display("Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:654 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n");
              if (1)$display("");
            end 
         if (_GEN_28&grantIsUncached&_GEN_18&~reset&~uncachedInFlight_0)
            begin 
              if (1)$display("Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:664 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n");
              if (1)$display("");
            end 
         if (_GEN_28&~grantIsUncached&grantIsVoluntary&~reset&~release_ack_wait)
            begin 
              if (1)$display("Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:685 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n");
              if (1)$display("");
            end 
         if (~reset&(auto_out_e_ready&nodeOut_e_valid)!=(_io_errors_bus_valid_T&~(|counter)&grantIsCached))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:693 assert(tl_out.e.fire === (tl_out.d.fire && d_first && grantIsCached))\n");
              if (1)$display("");
            end 
         if (s2_want_victimize&~reset&~(s2_valid_flush_line|s2_flush_valid|io_cpu_s2_nack_0))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:794 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n");
              if (1)$display("");
            end 
         if (doUncachedResp&~reset&s2_valid_hit_pre_data_ecc_and_waw)
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:928 assert(!s2_valid_hit)\n");
              if (1)$display("");
            end 
       end
  
   wire [31:0] io_cpu_resp_bits_data_zeroed=s2_req_addr[2] ? s2_data[63:32]:s2_data[31:0] ;  
   wire _io_cpu_resp_bits_data_word_bypass_T_1=s2_req_size==2'h2 ;  
   wire [15:0] io_cpu_resp_bits_data_zeroed_1=s2_req_addr[1] ? io_cpu_resp_bits_data_zeroed[31:16]:io_cpu_resp_bits_data_zeroed[15:0] ;  
   wire [7:0] io_cpu_resp_bits_data_zeroed_2=s2_sc ? 8'h0:s2_req_addr[0] ? io_cpu_resp_bits_data_zeroed_1[15:8]:io_cpu_resp_bits_data_zeroed_1[7:0] ;  
   wire [31:0] io_cpu_resp_bits_data_word_bypass_zeroed=s2_req_addr[2] ? s2_data[63:32]:s2_data[31:0] ;  
   reg REG ;  
   wire [26:0] _io_cpu_perf_release_beats1_decode_T_1=27'hFFF<<_GEN_23 ;  
   wire [8:0] io_cpu_perf_release_beats1=nodeOut_c_bits_opcode[0] ? ~(_io_cpu_perf_release_beats1_decode_T_1[11:3]):9'h0 ;  
   reg [8:0] io_cpu_perf_release_counter ;  
   wire [3:0] _release_state_T_14=s2_victim_dirty&~(s2_valid_flush_line&s2_req_size[1]) ? 4'h1:4'h6 ;  
   wire [3:0] _release_state_T_15={1'h0,releaseDone,2'h3} ;  
   wire [3:0] _GEN_29=s2_prb_ack_data ? 4'h2:(|s2_probe_state_state) ? 4'h3:4'h5 ;  
   wire [3:0] _GEN_30=s2_want_victimize ? _release_state_T_14:release_state ;  
   wire [3:0] _GEN_31=s2_probe ? _GEN_29:_GEN_30 ;  
   wire _GEN_32=_io_errors_bus_valid_T&grantIsCached&d_last ;  
   wire _GEN_33=_GEN_24&~metaArb__grant_T_3 ;  
   wire [6:0] flushCounterNext={1'h0,flushCounter}+7'h1 ;  
   wire _GEN_34=_GEN_25&releaseDone|_GEN_33 ;  
   wire [33:0] s0_req_addr={resetting ? {io_cpu_req_bits_addr[33:12],flushCounter}:_GEN ? {io_cpu_req_bits_addr[33:12],s2_req_addr[11:6]}:metaArb_io_in_valid_4 ? {io_cpu_req_bits_addr[33:12],probe_bits_address[11:6]}:metaArb_io_in_valid_6 ? {io_cpu_req_bits_addr[33:32],_GEN_24 ? probe_bits_address[31:6]:auto_out_b_bits_address[31:6]}:io_cpu_req_bits_addr[33:6],io_cpu_req_bits_addr[5:0]} ;  
   wire [9:0] _GEN_35=s1_tlb_req_vaddr[25:16]^10'h200 ;  
   wire [3:0] _GEN_36=s1_tlb_req_vaddr[31:28]^4'h8 ;  
   wire tlb_legal_address={s1_tlb_req_vaddr[33:14],~(s1_tlb_req_vaddr[13:12])}==22'h0|{s1_tlb_req_vaddr[33:28],~(s1_tlb_req_vaddr[27:26])}==8'h0|{s1_tlb_req_vaddr[33:26],_GEN_35}==18'h0|~(|(s1_tlb_req_vaddr[33:12]))|{s1_tlb_req_vaddr[33:17],~(s1_tlb_req_vaddr[16])}==18'h0|{s1_tlb_req_vaddr[33:32],_GEN_36}==6'h0|{s1_tlb_req_vaddr[33:31],~(s1_tlb_req_vaddr[30:29])}==5'h0 ;  
   wire tlb_cacheable=tlb_legal_address&~(_GEN_36[3]) ;  
   wire tlb_deny_access_to_debug=~io_ptw_status_debug&~(|(s1_tlb_req_vaddr[33:12])) ;  
   wire [3:0] _GEN_37={s1_tlb_req_vaddr[31:30],s1_tlb_req_vaddr[27],s1_tlb_req_vaddr[16]} ;  
   wire [2:0] _GEN_38={s1_tlb_req_vaddr[31:30],~(s1_tlb_req_vaddr[27])} ;  
   wire [1:0] _GEN_39={s1_tlb_req_vaddr[31],~(s1_tlb_req_vaddr[30])} ;  
   wire [3:0] _GEN_40=s1_tlb_req_vaddr[3:0]&(4'h1<<s1_tlb_req_size)-4'h1 ;  
   wire tlb__cmd_lrsc_T=s1_tlb_req_cmd==5'h6 ;  
   wire tlb__cmd_lrsc_T_1=s1_tlb_req_cmd==5'h7 ;  
   wire tlb__cmd_read_T_7=s1_tlb_req_cmd==5'h4 ;  
   wire tlb__cmd_read_T_8=s1_tlb_req_cmd==5'h9 ;  
   wire tlb__cmd_read_T_9=s1_tlb_req_cmd==5'hA ;  
   wire tlb__cmd_read_T_10=s1_tlb_req_cmd==5'hB ;  
   wire tlb__cmd_read_T_14=s1_tlb_req_cmd==5'h8 ;  
   wire tlb__cmd_read_T_15=s1_tlb_req_cmd==5'hC ;  
   wire tlb__cmd_read_T_16=s1_tlb_req_cmd==5'hD ;  
   wire tlb__cmd_read_T_17=s1_tlb_req_cmd==5'hE ;  
   wire tlb__cmd_read_T_18=s1_tlb_req_cmd==5'hF ;  
   wire tlb_cmd_put_partial=s1_tlb_req_cmd==5'h11 ;  
   wire tlb_cmd_read=s1_tlb_req_cmd==5'h0|s1_tlb_req_cmd==5'h10|tlb__cmd_lrsc_T|tlb__cmd_lrsc_T_1|tlb__cmd_read_T_7|tlb__cmd_read_T_8|tlb__cmd_read_T_9|tlb__cmd_read_T_10|tlb__cmd_read_T_14|tlb__cmd_read_T_15|tlb__cmd_read_T_16|tlb__cmd_read_T_17|tlb__cmd_read_T_18 ;  
   wire tlb_cmd_write=s1_tlb_req_cmd==5'h1|tlb_cmd_put_partial|tlb__cmd_lrsc_T_1|tlb__cmd_read_T_7|tlb__cmd_read_T_8|tlb__cmd_read_T_9|tlb__cmd_read_T_10|tlb__cmd_read_T_14|tlb__cmd_read_T_15|tlb__cmd_read_T_16|tlb__cmd_read_T_17|tlb__cmd_read_T_18 ;  
   wire tlb_ae_array=(|_GEN_40)&tlb_legal_address&({s1_tlb_req_vaddr[31:30],s1_tlb_req_vaddr[27],s1_tlb_req_vaddr[25],s1_tlb_req_vaddr[16],s1_tlb_req_vaddr[13]}==6'h0|{s1_tlb_req_vaddr[31:30],s1_tlb_req_vaddr[27],_GEN_35[9],s1_tlb_req_vaddr[16]}==5'h0|~(|_GEN_38)|~(|_GEN_39))|(tlb__cmd_lrsc_T|tlb__cmd_lrsc_T_1)&~tlb_cacheable ;  
   wire [1:0] _s2_data_T_1=io_cpu_replay_next_0|inWriteback|s1_did_read ? (_GEN_19 ? 2'h1:2'h2):2'h0 ;  
   wire _probe_bits_T=nodeOut_b_ready&auto_out_b_valid ;  
   wire s1_valid_not_nacked=s1_valid&~s1_nack ;  
   wire _s1_meta_hit_state_T_2=_tag_array_0_ext_RW0_rdata[19:0]==s1_tlb_req_vaddr[31:12]&~s1_flush_valid ;  
   wire _s2_victim_way_T=s1_valid_not_nacked|s1_flush_valid ;  
   wire _GEN_41=s2_valid_hit_pre_data_ecc_and_waw&s2_lr&~cached_grant_wait|s2_valid_cached_miss ;  
   wire advance_pstore1=pstore1_valid&pstore2_valid==pstore_drain ;  
   wire _io_cpu_perf_acquire_T=auto_out_a_ready&tl_out_a_valid ;  
   wire _GEN_42=_io_cpu_perf_acquire_T&~s2_pma_cacheable ;  
   wire _GEN_43=_GEN_27&_io_cpu_perf_release_T&c_first ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              s1_valid <=1'h0;
              s1_probe <=1'h0;
              cached_grant_wait <=1'h0;
              resetting <=1'h0;
              flushCounter <=6'h0;
              release_ack_wait <=1'h0;
              release_state <=4'h0;
              uncachedInFlight_0 <=1'h0;
              s2_valid <=1'h0;
              s2_probe <=1'h0;
              lrscCount <=7'h0;
              pstore2_valid <=1'h0;
              pstore1_held <=1'h0;
              counter <=9'h0;
              grantInProgress <=1'h0;
              blockProbeAfterGrantCount <=3'h0;
              counter_1 <=9'h0;
              io_cpu_perf_release_counter <=9'h0;
            end 
          else 
            begin 
              s1_valid <=io_cpu_req_ready_0&io_cpu_req_valid;
              s1_probe <=_GEN_33|_probe_bits_T;
              cached_grant_wait <=~_GEN_32&(_io_cpu_perf_acquire_T&s2_pma_cacheable|cached_grant_wait);
              resetting <=~(resetting&flushCounterNext[6])&(REG|resetting);
              if (resetting)
                 flushCounter <=flushCounterNext[5:0];
              release_ack_wait <=_GEN_43|(~_io_errors_bus_valid_T|grantIsCached|grantIsUncached|~grantIsVoluntary)&release_ack_wait;
              if (~metaArb__grant_T_2&metaArb_io_in_valid_4)
                 release_state <=4'h0;
               else 
                 if (_GEN_27)
                    begin 
                      if (releaseDone)
                         release_state <=4'h6;
                       else 
                         if (_GEN_26)
                            release_state <=_inWriteback_T_1 ? (_GEN_34 ? 4'h0:_GEN_31):_GEN_25 ? (releaseDone|_GEN_33 ? 4'h0:_GEN_31):_GEN_33 ? 4'h0:s2_probe ? (s2_prb_ack_data ? 4'h2:(|s2_probe_state_state) ? 4'h3:releaseDone ? 4'h0:4'h5):_GEN_30;
                          else 
                            if (_GEN_34)
                               release_state <=4'h0;
                             else 
                               if (s2_probe)
                                  begin 
                                    if (s2_prb_ack_data)
                                       release_state <=4'h2;
                                     else 
                                       if (|s2_probe_state_state)
                                          release_state <=_release_state_T_15;
                                        else 
                                          if (releaseDone)
                                             release_state <=4'h0;
                                           else 
                                             release_state <=4'h5;
                                  end 
                                else 
                                  if (s2_want_victimize)
                                     release_state <=_release_state_T_14;
                    end 
                  else 
                    if (_inWriteback_T_1)
                       begin 
                         if (releaseDone)
                            release_state <=4'h7;
                          else 
                            if (_GEN_34)
                               release_state <=4'h0;
                             else 
                               if (s2_probe)
                                  release_state <=_GEN_29;
                                else 
                                  if (s2_want_victimize)
                                     release_state <=_release_state_T_14;
                       end 
                     else 
                       if (_GEN_26)
                          begin 
                            if (releaseDone)
                               release_state <=4'h7;
                             else 
                               if (_GEN_34)
                                  release_state <=4'h0;
                                else 
                                  if (s2_probe)
                                     release_state <=_GEN_29;
                                   else 
                                     if (s2_want_victimize)
                                        release_state <=_release_state_T_14;
                          end 
                        else 
                          if (_GEN_34)
                             release_state <=4'h0;
                           else 
                             if (s2_probe)
                                begin 
                                  if (s2_prb_ack_data)
                                     release_state <=4'h2;
                                   else 
                                     if (|s2_probe_state_state)
                                        release_state <=_release_state_T_15;
                                      else 
                                        if (releaseDone)
                                           release_state <=4'h0;
                                         else 
                                           release_state <=4'h5;
                                end 
                              else 
                                if (s2_want_victimize)
                                   release_state <=_release_state_T_14;
              uncachedInFlight_0 <=(~_io_errors_bus_valid_T|grantIsCached|~(grantIsUncached&_GEN_18))&(_GEN_42|uncachedInFlight_0);
              s2_valid <=s1_valid_masked&~(s1_req_cmd==5'h14|s1_req_cmd==5'h15|s1_req_cmd==5'h16);
              s2_probe <=s1_probe;
              if (s1_probe)
                 lrscCount <=7'h0;
               else 
                 if (s2_valid_masked&(|(lrscCount[6:2])))
                    lrscCount <=7'h3;
                  else 
                    if (|lrscCount)
                       lrscCount <=lrscCount-7'h1;
                     else 
                       if (_GEN_41)
                          lrscCount <=s2_hit ? 7'h4F:7'h0;
              pstore2_valid <=pstore2_valid&~pstore_drain|advance_pstore1;
              pstore1_held <=(_pstore1_held_T&~s2_sc_fail|pstore1_held)&pstore2_valid&~pstore_drain;
              if (_io_errors_bus_valid_T)
                 begin 
                   if (|counter)
                      counter <=_counter1_T;
                    else 
                      counter <=beats1;
                 end 
              if (_GEN_17)
                 grantInProgress <=~d_last;
              if (_GEN_32)
                 blockProbeAfterGrantCount <=3'h7;
               else 
                 if (|blockProbeAfterGrantCount)
                    blockProbeAfterGrantCount <=blockProbeAfterGrantCount-3'h1;
              if (_io_cpu_perf_release_T)
                 begin 
                   if (c_first)
                      counter_1 <=beats1_1;
                    else 
                      counter_1 <=_counter1_T_1;
                   if (io_cpu_perf_release_counter==9'h0)
                      io_cpu_perf_release_counter <=io_cpu_perf_release_beats1;
                    else 
                      io_cpu_perf_release_counter <=io_cpu_perf_release_counter-9'h1;
                 end 
            end 
         if (s2_want_victimize)
            begin 
              probe_bits_param <=2'h0;
              probe_bits_size <=4'h0;
              probe_bits_address <={s2_valid_flush_line ? s2_req_addr[31:12]:s2_meta_corrected_r[19:0],s2_req_addr[11:6],6'h0};
            end 
          else 
            if (_probe_bits_T)
               begin 
                 probe_bits_param <=auto_out_b_bits_param;
                 probe_bits_size <=auto_out_b_bits_size;
                 probe_bits_address <=auto_out_b_bits_address;
               end 
         probe_bits_source <=~s2_want_victimize&(_probe_bits_T ? auto_out_b_bits_source:probe_bits_source);
         if (metaArb_io_out_valid&~metaArb_io_out_bits_write)
            begin 
              s1_vaddr <=s0_req_addr;
              s1_req_tag <=io_cpu_req_bits_tag;
              s1_req_cmd <=io_cpu_req_bits_cmd;
              s1_req_size <=io_cpu_req_bits_size;
              s1_req_signed <=io_cpu_req_bits_signed;
              s1_req_dprv <=2'h3;
              s1_req_dv <=io_cpu_req_bits_dv;
              s1_tlb_req_vaddr <=s0_req_addr;
              s1_tlb_req_size <=io_cpu_req_bits_size;
              s1_tlb_req_cmd <=io_cpu_req_bits_cmd;
              s1_tlb_req_prv <=2'h3;
              s1_did_read <=~dataArb__grant_T_1&io_cpu_req_valid&(_pstore_drain_opportunistic_T|_pstore_drain_opportunistic_T_1|_pstore_drain_opportunistic_T_2|_pstore_drain_opportunistic_T_28|_pstore_drain_opportunistic_T_30|_pstore_drain_opportunistic_T_31|_pstore_drain_opportunistic_T_32|_pstore_drain_opportunistic_T_33|_pstore_drain_opportunistic_T_37|_pstore_drain_opportunistic_T_38|_pstore_drain_opportunistic_T_39|_pstore_drain_opportunistic_T_40|_pstore_drain_opportunistic_T_41|(_pstore_drain_opportunistic_T_25|_pstore_drain_opportunistic_T_50|_pstore_drain_opportunistic_T_28|_pstore_drain_opportunistic_T_30|_pstore_drain_opportunistic_T_31|_pstore_drain_opportunistic_T_32|_pstore_drain_opportunistic_T_33|_pstore_drain_opportunistic_T_37|_pstore_drain_opportunistic_T_38|_pstore_drain_opportunistic_T_39|_pstore_drain_opportunistic_T_40|_pstore_drain_opportunistic_T_41)&_pstore_drain_opportunistic_T_50);
            end 
         s1_flush_valid <=1'h0;
         if (_GEN_43)
            release_ack_addr <=probe_bits_address;
         if (_GEN_42)
            begin 
              uncachedReqs_addr_0 <=s2_req_addr;
              uncachedReqs_tag_0 <=s2_req_tag;
              uncachedReqs_size_0 <=s2_req_size;
              uncachedReqs_signed_0 <=s2_req_signed;
            end 
         s2_not_nacked_in_s1 <=~s1_nack;
         if (_GEN_19)
            begin 
              if (_s2_victim_way_T)
                 begin 
                   s2_req_addr <={2'h0,s1_tlb_req_vaddr[31:12],s1_vaddr[11:0]};
                   s2_req_tag <=s1_req_tag;
                   s2_req_cmd <=s1_req_cmd;
                   s2_req_size <=s1_req_size;
                   s2_req_signed <=s1_req_signed;
                 end 
            end 
          else 
            begin 
              s2_req_addr <={2'h0,s1_tlb_req_vaddr[31:12],s1_vaddr[11:3],uncachedReqs_addr_0[2:0]};
              s2_req_tag <=uncachedReqs_tag_0;
              s2_req_cmd <=5'h0;
              s2_req_size <=uncachedReqs_size_0;
              s2_req_signed <=uncachedReqs_signed_0;
            end 
         if (_s2_victim_way_T)
            begin 
              s2_req_dprv <=s1_req_dprv;
              s2_req_dv <=s1_req_dv;
              s2_tlb_xcpt_ae_ld <=tlb_cmd_read&(tlb_ae_array|~(tlb_legal_address&~tlb_deny_access_to_debug&_tlb_pmp_io_r));
              s2_tlb_xcpt_ae_st <=(tlb_cmd_write|s1_tlb_req_cmd==5'h5|s1_tlb_req_cmd==5'h17)&(tlb_ae_array|~(tlb_legal_address&(~(|_GEN_37)|~(|_GEN_38)|~(|_GEN_39)|~(|(_GEN_36[3:2])))&~tlb_deny_access_to_debug&_tlb_pmp_io_w))|tlb_cmd_put_partial&~(tlb_legal_address&(~(|_GEN_37)|~(|_GEN_38)|~(|_GEN_39)|~(|(_GEN_36[3:2])))|tlb_cacheable)|(tlb__cmd_read_T_7|tlb__cmd_read_T_8|tlb__cmd_read_T_9|tlb__cmd_read_T_10)&~(tlb_legal_address&(~(|_GEN_37)|~(|_GEN_38))|tlb_cacheable)|(tlb__cmd_read_T_14|tlb__cmd_read_T_15|tlb__cmd_read_T_16|tlb__cmd_read_T_17|tlb__cmd_read_T_18)&~(tlb_legal_address&(~(|_GEN_37)|~(|_GEN_38))|tlb_cacheable);
              s2_tlb_xcpt_ma_ld <=(|_GEN_40)&tlb_cmd_read;
              s2_tlb_xcpt_ma_st <=(|_GEN_40)&tlb_cmd_write;
              s2_pma_cacheable <=tlb_cacheable;
              s2_vaddr_r <=s1_vaddr;
              if (_s1_meta_hit_state_T_2)
                 s2_hit_state_state <=_tag_array_0_ext_RW0_rdata[21:20];
               else 
                 s2_hit_state_state <=2'h0;
            end 
         s2_tlb_xcpt_pf_ld <=~_s2_victim_way_T&s2_tlb_xcpt_pf_ld;
         s2_tlb_xcpt_pf_st <=~_s2_victim_way_T&s2_tlb_xcpt_pf_st;
         if (_GEN_19)
            begin 
            end 
          else 
            s2_uncached_resp_addr <=uncachedReqs_addr_0;
         s2_flush_valid <=s1_flush_valid;
         if (_s2_victim_way_T|s1_probe)
            s2_meta_corrected_r <=_tag_array_0_ext_RW0_rdata;
         if (s1_valid|inWriteback|io_cpu_replay_next_0)
            s2_data <=(_s2_data_T_1[0] ? _data_io_resp_0:64'h0)|(_s2_data_T_1[1] ? auto_out_d_bits_data:64'h0);
         if (s1_probe)
            begin 
              if (_s1_meta_hit_state_T_2)
                 s2_probe_state_state <=_tag_array_0_ext_RW0_rdata[21:20];
               else 
                 s2_probe_state_state <=2'h0;
            end 
         if (_GEN_41)
            lrscAddr <=s2_req_addr[33:6];
         if (s1_valid_not_nacked&s1_write)
            begin 
              pstore1_cmd <=s1_req_cmd;
              pstore1_addr <=s1_vaddr;
              pstore1_data <=io_cpu_s1_data_data;
              pstore1_mask <=_io_cpu_perf_canAcceptLoadThenLoad_T_51 ? io_cpu_s1_data_mask:s1_mask_xwr;
              pstore1_rmw <=_io_cpu_perf_canAcceptLoadThenLoad_T_1|_io_cpu_perf_canAcceptLoadThenLoad_T_2|_io_cpu_perf_canAcceptLoadThenLoad_T_3|_io_cpu_perf_canAcceptLoadThenLoad_T_29|_io_cpu_perf_canAcceptLoadThenLoad_T_31|_io_cpu_perf_canAcceptLoadThenLoad_T_32|_io_cpu_perf_canAcceptLoadThenLoad_T_33|_io_cpu_perf_canAcceptLoadThenLoad_T_34|_io_cpu_perf_canAcceptLoadThenLoad_T_38|_io_cpu_perf_canAcceptLoadThenLoad_T_39|_io_cpu_perf_canAcceptLoadThenLoad_T_40|_io_cpu_perf_canAcceptLoadThenLoad_T_41|_io_cpu_perf_canAcceptLoadThenLoad_T_42|(_io_cpu_perf_canAcceptLoadThenLoad_T_26|_io_cpu_perf_canAcceptLoadThenLoad_T_51|_io_cpu_perf_canAcceptLoadThenLoad_T_29|_io_cpu_perf_canAcceptLoadThenLoad_T_31|_io_cpu_perf_canAcceptLoadThenLoad_T_32|_io_cpu_perf_canAcceptLoadThenLoad_T_33|_io_cpu_perf_canAcceptLoadThenLoad_T_34|_io_cpu_perf_canAcceptLoadThenLoad_T_38|_io_cpu_perf_canAcceptLoadThenLoad_T_39|_io_cpu_perf_canAcceptLoadThenLoad_T_40|_io_cpu_perf_canAcceptLoadThenLoad_T_41|_io_cpu_perf_canAcceptLoadThenLoad_T_42)&_io_cpu_perf_canAcceptLoadThenLoad_T_51;
            end 
         pstore_drain_on_miss_REG <=io_cpu_s2_nack_0;
         if (advance_pstore1)
            begin 
              pstore2_addr <=pstore1_addr;
              pstore2_storegen_data_r <=_amoalus_0_io_out[7:0];
              pstore2_storegen_data_r_1 <=_amoalus_0_io_out[15:8];
              pstore2_storegen_data_r_2 <=_amoalus_0_io_out[23:16];
              pstore2_storegen_data_r_3 <=_amoalus_0_io_out[31:24];
              pstore2_storegen_data_r_4 <=_amoalus_0_io_out[39:32];
              pstore2_storegen_data_r_5 <=_amoalus_0_io_out[47:40];
              pstore2_storegen_data_r_6 <=_amoalus_0_io_out[55:48];
              pstore2_storegen_data_r_7 <=_amoalus_0_io_out[63:56];
              pstore2_storegen_mask <=pstore1_mask;
            end 
         if (_GEN_22)
            blockUncachedGrant <=dataArb_io_in_valid_0;
          else 
            blockUncachedGrant <=dataArb_io_out_valid;
         s1_release_data_valid <=~dataArb__grant_T&dataArb_io_in_valid_2;
         s2_release_data_valid <=s1_release_data_valid&~releaseRejected;
         io_cpu_s2_xcpt_REG <=s1_valid&~io_cpu_s1_kill&(s1_read|s1_write|s1_req_cmd==5'h5&s1_req_size[0]|s1_req_cmd==5'h17)&~s1_nack;
         doUncachedResp <=io_cpu_replay_next_0;
         REG <=reset;
       end
  
  PMPChecker tlb_pmp(.io_prv(s1_tlb_req_prv),.io_pmp_cfg_l_0(io_ptw_pmp_cfg_l_0),.io_pmp_cfg_l_1(io_ptw_pmp_cfg_l_1),.io_pmp_cfg_l_2(io_ptw_pmp_cfg_l_2),.io_pmp_cfg_l_3(io_ptw_pmp_cfg_l_3),.io_pmp_cfg_l_4(io_ptw_pmp_cfg_l_4),.io_pmp_cfg_l_5(io_ptw_pmp_cfg_l_5),.io_pmp_cfg_l_6(io_ptw_pmp_cfg_l_6),.io_pmp_cfg_l_7(io_ptw_pmp_cfg_l_7),.io_pmp_cfg_a_0(io_ptw_pmp_cfg_a_0),.io_pmp_cfg_a_1(io_ptw_pmp_cfg_a_1),.io_pmp_cfg_a_2(io_ptw_pmp_cfg_a_2),.io_pmp_cfg_a_3(io_ptw_pmp_cfg_a_3),.io_pmp_cfg_a_4(io_ptw_pmp_cfg_a_4),.io_pmp_cfg_a_5(io_ptw_pmp_cfg_a_5),.io_pmp_cfg_a_6(io_ptw_pmp_cfg_a_6),.io_pmp_cfg_a_7(io_ptw_pmp_cfg_a_7),.io_pmp_cfg_w_0(io_ptw_pmp_cfg_w_0),.io_pmp_cfg_w_1(io_ptw_pmp_cfg_w_1),.io_pmp_cfg_w_2(io_ptw_pmp_cfg_w_2),.io_pmp_cfg_w_3(io_ptw_pmp_cfg_w_3),.io_pmp_cfg_w_4(io_ptw_pmp_cfg_w_4),.io_pmp_cfg_w_5(io_ptw_pmp_cfg_w_5),.io_pmp_cfg_w_6(io_ptw_pmp_cfg_w_6),.io_pmp_cfg_w_7(io_ptw_pmp_cfg_w_7),.io_pmp_cfg_r_0(io_ptw_pmp_cfg_r_0),.io_pmp_cfg_r_1(io_ptw_pmp_cfg_r_1),.io_pmp_cfg_r_2(io_ptw_pmp_cfg_r_2),.io_pmp_cfg_r_3(io_ptw_pmp_cfg_r_3),.io_pmp_cfg_r_4(io_ptw_pmp_cfg_r_4),.io_pmp_cfg_r_5(io_ptw_pmp_cfg_r_5),.io_pmp_cfg_r_6(io_ptw_pmp_cfg_r_6),.io_pmp_cfg_r_7(io_ptw_pmp_cfg_r_7),.io_pmp_addr_0(io_ptw_pmp_addr_0),.io_pmp_addr_1(io_ptw_pmp_addr_1),.io_pmp_addr_2(io_ptw_pmp_addr_2),.io_pmp_addr_3(io_ptw_pmp_addr_3),.io_pmp_addr_4(io_ptw_pmp_addr_4),.io_pmp_addr_5(io_ptw_pmp_addr_5),.io_pmp_addr_6(io_ptw_pmp_addr_6),.io_pmp_addr_7(io_ptw_pmp_addr_7),.io_pmp_mask_0(io_ptw_pmp_mask_0),.io_pmp_mask_1(io_ptw_pmp_mask_1),.io_pmp_mask_2(io_ptw_pmp_mask_2),.io_pmp_mask_3(io_ptw_pmp_mask_3),.io_pmp_mask_4(io_ptw_pmp_mask_4),.io_pmp_mask_5(io_ptw_pmp_mask_5),.io_pmp_mask_6(io_ptw_pmp_mask_6),.io_pmp_mask_7(io_ptw_pmp_mask_7),.io_addr(s1_tlb_req_vaddr[31:0]),.io_size(s1_tlb_req_size),.io_r(_tlb_pmp_io_r),.io_w(_tlb_pmp_io_w)); 
  OptimizationBarrier tlb_entries_barrier(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier tlb_entries_barrier_1(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier tlb_entries_barrier_2(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier tlb_entries_barrier_3(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier tlb_entries_barrier_4(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier tlb_entries_barrier_5(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier pma_checker_entries_barrier(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier pma_checker_entries_barrier_1(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier pma_checker_entries_barrier_2(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier pma_checker_entries_barrier_3(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier pma_checker_entries_barrier_4(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  tag_array_0_64x22 tag_array_0_ext(.RW0_addr(resetting ? flushCounter:_GEN ? metaArb_io_in_bits_idx_3:metaArb_io_in_valid_4 ? metaArb_io_in_bits_idx_4:metaArb_io_in_valid_6 ? metaArb_io_in_bits_idx_6:metaArb_io_in_bits_idx_7),.RW0_en(readEnable|writeEnable),.RW0_clk(clock),.RW0_wmode(metaArb_io_out_bits_write),.RW0_wdata(resetting ? 22'h0:metaArb_io_in_valid_2 ? metaArb_io_in_bits_data_2:metaArb_io_in_valid_3 ? metaArb_io_in_bits_data_3:metaArb_io_in_bits_data_7),.RW0_rdata(_tag_array_0_ext_RW0_rdata)); 
  DCacheDataArray data(.clock(clock),.io_req_valid(dataArb_io_out_valid),.io_req_bits_addr(dataArb_io_in_valid_0 ? _dataArb_io_in_0_bits_wordMask_wordMask_T:dataArb_io_in_valid_1 ? dataArb_io_in_bits_addr_1:dataArb_io_in_valid_2 ? dataArb_io_in_bits_addr_2:dataArb_io_in_bits_addr_3),.io_req_bits_write(dataArb_io_in_valid_0 ? pstore_drain:dataArb_io_in_valid_1&dataArb_io_in_bits_write_1),.io_req_bits_wdata(dataArb_io_in_valid_0 ? dataArb_io_in_bits_wdata_0:auto_out_d_bits_data),.io_req_bits_eccMask(dataArb_io_in_valid_0 ? dataArb_io_in_bits_eccMask_0:8'hFF),.io_resp_0(_data_io_resp_0)); 
  AMOALU amoalus_0(.io_mask(pstore1_mask),.io_cmd(pstore1_cmd),.io_lhs(s2_data),.io_rhs(pstore1_data),.io_out(_amoalus_0_io_out)); 
  assign auto_out_a_valid=tl_out_a_valid; 
  assign auto_out_a_bits_opcode=s2_pma_cacheable ? 3'h6:s2_write ? (_metaArb_io_in_3_bits_data_c_cat_T_24 ? 3'h1:s2_read ? (_metaArb_io_in_3_bits_data_c_cat_T_39|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_35 ? 3'h2:_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_28 ? 3'h3:3'h0):3'h0):3'h4; 
  assign auto_out_a_bits_param=s2_pma_cacheable ? {1'h0,casez_tmp}:~s2_write|_metaArb_io_in_3_bits_data_c_cat_T_24|~s2_read ? 3'h0:_metaArb_io_in_3_bits_data_c_cat_T_39 ? 3'h3:_metaArb_io_in_3_bits_data_c_cat_T_38 ? 3'h2:_metaArb_io_in_3_bits_data_c_cat_T_37 ? 3'h1:_metaArb_io_in_3_bits_data_c_cat_T_36 ? 3'h0:_metaArb_io_in_3_bits_data_c_cat_T_35 ? 3'h4:_metaArb_io_in_3_bits_data_c_cat_T_31 ? 3'h2:_metaArb_io_in_3_bits_data_c_cat_T_30 ? 3'h1:_metaArb_io_in_3_bits_data_c_cat_T_29|~_metaArb_io_in_3_bits_data_c_cat_T_28 ? 3'h0:3'h3; 
  assign auto_out_a_bits_size=s2_pma_cacheable ? 4'h6:_GEN_16 ? {2'h0,s2_req_size}:4'h0; 
  assign auto_out_a_bits_source=~s2_pma_cacheable&(~s2_write|_metaArb_io_in_3_bits_data_c_cat_T_24|~s2_read|_metaArb_io_in_3_bits_data_c_cat_T_39|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_28); 
  assign auto_out_a_bits_address=s2_pma_cacheable ? {s2_req_addr[31:6],6'h0}:_GEN_16 ? s2_req_addr[31:0]:32'h0; 
  assign auto_out_a_bits_mask=s2_pma_cacheable ? 8'hFF:s2_write ? (_metaArb_io_in_3_bits_data_c_cat_T_24 ? pstore1_mask:s2_read ? atomics_mask:{put_a_mask_acc_5|put_a_mask_eq_5&s2_req_addr[0],put_a_mask_acc_5|put_a_mask_eq_5&~(s2_req_addr[0]),put_a_mask_acc_4|put_a_mask_eq_4&s2_req_addr[0],put_a_mask_acc_4|put_a_mask_eq_4&~(s2_req_addr[0]),put_a_mask_acc_3|put_a_mask_eq_3&s2_req_addr[0],put_a_mask_acc_3|put_a_mask_eq_3&~(s2_req_addr[0]),put_a_mask_acc_2|put_a_mask_eq_2&s2_req_addr[0],put_a_mask_acc_2|put_a_mask_eq_2&~(s2_req_addr[0])}):{get_a_mask_acc_5|get_a_mask_eq_5&s2_req_addr[0],get_a_mask_acc_5|get_a_mask_eq_5&~(s2_req_addr[0]),get_a_mask_acc_4|get_a_mask_eq_4&s2_req_addr[0],get_a_mask_acc_4|get_a_mask_eq_4&~(s2_req_addr[0]),get_a_mask_acc_3|get_a_mask_eq_3&s2_req_addr[0],get_a_mask_acc_3|get_a_mask_eq_3&~(s2_req_addr[0]),get_a_mask_acc_2|get_a_mask_eq_2&s2_req_addr[0],get_a_mask_acc_2|get_a_mask_eq_2&~(s2_req_addr[0])}; 
  assign auto_out_a_bits_data=s2_pma_cacheable|~s2_write|~(_metaArb_io_in_3_bits_data_c_cat_T_24|~s2_read|_metaArb_io_in_3_bits_data_c_cat_T_39|_metaArb_io_in_3_bits_data_c_cat_T_38|_metaArb_io_in_3_bits_data_c_cat_T_37|_metaArb_io_in_3_bits_data_c_cat_T_36|_metaArb_io_in_3_bits_data_c_cat_T_35|_metaArb_io_in_3_bits_data_c_cat_T_31|_metaArb_io_in_3_bits_data_c_cat_T_30|_metaArb_io_in_3_bits_data_c_cat_T_29|_metaArb_io_in_3_bits_data_c_cat_T_28) ? 64'h0:pstore1_data; 
  assign auto_out_b_ready=nodeOut_b_ready; 
  assign auto_out_c_valid=nodeOut_c_valid; 
  assign auto_out_c_bits_opcode=nodeOut_c_bits_opcode; 
  assign auto_out_c_bits_param=_GEN_27 ? ((&s2_victim_state_state)|s2_victim_state_state==2'h2 ? 3'h1:s2_victim_state_state==2'h1 ? 3'h2:s2_victim_state_state==2'h0 ? 3'h5:3'h0):_inWriteback_T_1|_GEN_26|~(~s2_probe|s2_prb_ack_data|~(|s2_probe_state_state)) ? (_GEN_13 ? 3'h3:_GEN_10 ? 3'h4:_GEN_9 ? 3'h5:_GEN_8|_GEN_7 ? 3'h0:_GEN_6 ? 3'h4:_GEN_5 ? 3'h5:_GEN_4|_GEN_3==4'hA ? 3'h1:_GEN_3==4'h9 ? 3'h2:_GEN_3==4'h8 ? 3'h5:3'h0):3'h5; 
  assign auto_out_c_bits_size=nodeOut_c_bits_size; 
  assign auto_out_c_bits_source=probe_bits_source; 
  assign auto_out_c_bits_address=probe_bits_address; 
  assign auto_out_c_bits_data=s2_data; 
  assign auto_out_d_ready=nodeOut_d_ready; 
  assign auto_out_e_valid=nodeOut_e_valid; 
  assign auto_out_e_bits_sink=auto_out_d_bits_sink; 
  assign io_cpu_req_ready=io_cpu_req_ready_0; 
  assign io_cpu_s2_nack=io_cpu_s2_nack_0; 
  assign io_cpu_resp_valid=s2_valid_hit_pre_data_ecc_and_waw|doUncachedResp; 
  assign io_cpu_resp_bits_addr=doUncachedResp ? s2_uncached_resp_addr:s2_req_addr; 
  assign io_cpu_resp_bits_tag=s2_req_tag; 
  assign io_cpu_resp_bits_cmd=s2_req_cmd; 
  assign io_cpu_resp_bits_size=s2_req_size; 
  assign io_cpu_resp_bits_signed=s2_req_signed; 
  assign io_cpu_resp_bits_dprv=s2_req_dprv; 
  assign io_cpu_resp_bits_dv=s2_req_dv; 
  assign io_cpu_resp_bits_data={s2_req_size==2'h0|s2_sc ? {56{s2_req_signed&io_cpu_resp_bits_data_zeroed_2[7]}}:{s2_req_size==2'h1 ? {48{s2_req_signed&io_cpu_resp_bits_data_zeroed_1[15]}}:{_io_cpu_resp_bits_data_word_bypass_T_1 ? {32{s2_req_signed&io_cpu_resp_bits_data_zeroed[31]}}:s2_data[63:32],io_cpu_resp_bits_data_zeroed[31:16]},io_cpu_resp_bits_data_zeroed_1[15:8]},io_cpu_resp_bits_data_zeroed_2[7:1],io_cpu_resp_bits_data_zeroed_2[0]|s2_sc_fail}; 
  assign io_cpu_resp_bits_mask=8'h0; 
  assign io_cpu_resp_bits_replay=doUncachedResp; 
  assign io_cpu_resp_bits_has_data=s2_read; 
  assign io_cpu_resp_bits_data_word_bypass={_io_cpu_resp_bits_data_word_bypass_T_1 ? {32{s2_req_signed&io_cpu_resp_bits_data_word_bypass_zeroed[31]}}:s2_data[63:32],io_cpu_resp_bits_data_word_bypass_zeroed}; 
  assign io_cpu_resp_bits_data_raw=s2_data; 
  assign io_cpu_resp_bits_store_data=pstore1_data; 
  assign io_cpu_replay_next=io_cpu_replay_next_0; 
  assign io_cpu_s2_xcpt_ma_ld=io_cpu_s2_xcpt_ma_ld_0; 
  assign io_cpu_s2_xcpt_ma_st=io_cpu_s2_xcpt_ma_st_0; 
  assign io_cpu_s2_xcpt_pf_ld=io_cpu_s2_xcpt_pf_ld_0; 
  assign io_cpu_s2_xcpt_pf_st=io_cpu_s2_xcpt_pf_st_0; 
  assign io_cpu_s2_xcpt_ae_ld=io_cpu_s2_xcpt_ae_ld_0; 
  assign io_cpu_s2_xcpt_ae_st=io_cpu_s2_xcpt_ae_st_0; 
  assign io_cpu_ordered=~(s1_valid|s2_valid|cached_grant_wait|uncachedInFlight_0); 
  assign io_cpu_perf_release=(io_cpu_perf_release_counter==9'h1|io_cpu_perf_release_beats1==9'h0)&_io_cpu_perf_release_T; 
  assign io_cpu_perf_grant=auto_out_d_valid&d_last; 
  assign io_ptw_req_bits_bits_need_gpa=1'h0; 
  assign io_ptw_req_bits_bits_stage2=1'h0; 
endmodule
 
module tag_array_0_64x21 (
  input [5:0] RW0_addr,
  input RW0_en,
  input RW0_clk,
  input RW0_wmode,
  input [20:0] RW0_wdata,
  output [20:0] RW0_rdata) ; 
   reg [20:0] Memory[0:63] ;  
   reg [5:0] _RW0_raddr_d0 ;  
   reg _RW0_ren_d0 ;  
   reg _RW0_rmode_d0 ;  
  always @( posedge RW0_clk)
       begin 
         _RW0_raddr_d0 <=RW0_addr;
         _RW0_ren_d0 <=RW0_en;
         _RW0_rmode_d0 <=RW0_wmode;
         if (RW0_en&RW0_wmode&1'h1)
            Memory [RW0_addr]<=RW0_wdata;
       end
  
  assign RW0_rdata=_RW0_ren_d0&~_RW0_rmode_d0 ? Memory[_RW0_raddr_d0]:21'bx; 
endmodule
 
module data_arrays_512x32 (
  input [8:0] RW0_addr,
  input RW0_en,
  input RW0_clk,
  input RW0_wmode,
  input [31:0] RW0_wdata,
  output [31:0] RW0_rdata) ; 
   reg [31:0] Memory[0:511] ;  
   reg [8:0] _RW0_raddr_d0 ;  
   reg _RW0_ren_d0 ;  
   reg _RW0_rmode_d0 ;  
  always @( posedge RW0_clk)
       begin 
         _RW0_raddr_d0 <=RW0_addr;
         _RW0_ren_d0 <=RW0_en;
         _RW0_rmode_d0 <=RW0_wmode;
         if (RW0_en&RW0_wmode&1'h1)
            Memory [RW0_addr]<=RW0_wdata;
       end
  
  assign RW0_rdata=_RW0_ren_d0&~_RW0_rmode_d0 ? Memory[_RW0_raddr_d0]:32'bx; 
endmodule
 
module ICache (
  input clock,
  input reset,
  input auto_master_out_a_ready,
  output auto_master_out_a_valid,
  output [31:0] auto_master_out_a_bits_address,
  input auto_master_out_d_valid,
  input [2:0] auto_master_out_d_bits_opcode,
  input [3:0] auto_master_out_d_bits_size,
  input [63:0] auto_master_out_d_bits_data,
  input auto_master_out_d_bits_corrupt,
  input io_req_valid,
  input [32:0] io_req_bits_addr,
  input [31:0] io_s1_paddr,
  input io_s1_kill,
  input io_s2_kill,
  output io_resp_valid,
  output [31:0] io_resp_bits_data,
  output io_resp_bits_ae,
  input io_invalidate) ; 
   wire readEnable ;  
   wire writeEnable ;  
   wire readEnable_0 ;  
   wire wen ;  
   wire readEnable_1 ;  
   wire [5:0] _tag_rdata_T ;  
   wire io_req_ready ;  
   wire [31:0] _data_arrays_1_0_ext_RW0_rdata ;  
   wire [31:0] _data_arrays_0_0_ext_RW0_rdata ;  
   wire [20:0] _tag_array_0_ext_RW0_rdata ;  
   wire s0_valid=io_req_ready&io_req_valid ;  
   reg s1_valid ;  
   reg s2_valid ;  
   reg s2_hit ;  
   reg invalidated ;  
   reg refill_valid ;  
   wire s2_miss=s2_valid&~s2_hit&~io_s2_kill ;  
   reg s2_request_refill_REG ;  
   wire s2_request_refill=s2_miss&s2_request_refill_REG ;  
   reg [31:0] refill_paddr ;  
   wire refill_one_beat=auto_master_out_d_valid&auto_master_out_d_bits_opcode[0] ;  
  assign io_req_ready=~refill_one_beat; 
   wire [26:0] _beats1_decode_T_1=27'hFFF<<auto_master_out_d_bits_size ;  
   wire [8:0] beats1=auto_master_out_d_bits_opcode[0] ? ~(_beats1_decode_T_1[11:3]):9'h0 ;  
   reg [8:0] counter ;  
   wire [8:0] _counter1_T=counter-9'h1 ;  
   wire [8:0] refill_cnt=beats1&~_counter1_T ;  
   wire writeEnable_0=refill_one_beat&(counter==9'h1|beats1==9'h0)&auto_master_out_d_valid ;  
  assign _tag_rdata_T=io_req_bits_addr[11:6]; 
  assign readEnable_1=~writeEnable_0&s0_valid; 
   reg accruedRefillError ;  
   wire refillError=auto_master_out_d_bits_corrupt|(|refill_cnt)&accruedRefillError ;  
   reg [63:0] vb_array ;  
   wire [63:0] _s1_vb_T_1=vb_array>>io_s1_paddr[11:6] ;  
   wire s1_hit=_s1_vb_T_1[0]&_tag_array_0_ext_RW0_rdata[19:0]==io_s1_paddr[31:12] ;  
  assign wen=refill_one_beat&~invalidated; 
   wire [8:0] _mem_idx_T_6={refill_paddr[11:6],3'h0} ;  
  assign readEnable_0=~wen&s0_valid&~(io_req_bits_addr[2]); 
  assign writeEnable=refill_one_beat&~invalidated; 
  assign readEnable=~writeEnable&s0_valid&io_req_bits_addr[2]; 
   reg [31:0] s2_dout_0 ;  
   reg s2_tl_error ;  
   wire [127:0] _vb_array_T_3=128'h1<<refill_paddr[11:6] ;  
   wire _s1_can_request_refill_T=s2_miss|refill_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              s1_valid <=1'h0;
              s2_valid <=1'h0;
              refill_valid <=1'h0;
              counter <=9'h0;
              vb_array <=64'h0;
            end 
          else 
            begin 
              s1_valid <=s0_valid;
              s2_valid <=s1_valid&~io_s1_kill;
              refill_valid <=~writeEnable_0&(auto_master_out_a_ready&s2_request_refill|refill_valid);
              if (auto_master_out_d_valid)
                 begin 
                   if (counter==9'h0)
                      counter <=beats1;
                    else 
                      counter <=_counter1_T;
                 end 
              if (io_invalidate)
                 vb_array <=64'h0;
               else 
                 if (refill_one_beat)
                    vb_array <=writeEnable_0&~invalidated ? vb_array|_vb_array_T_3[63:0]:~(~vb_array|_vb_array_T_3[63:0]);
            end 
         s2_hit <=s1_hit;
         invalidated <=refill_valid&(io_invalidate|invalidated);
         s2_request_refill_REG <=~_s1_can_request_refill_T;
         if (s1_valid&~_s1_can_request_refill_T)
            refill_paddr <=io_s1_paddr;
         if (refill_one_beat)
            accruedRefillError <=refillError;
         if (s1_valid)
            begin 
              s2_dout_0 <=io_s1_paddr[2] ? _data_arrays_1_0_ext_RW0_rdata:_data_arrays_0_0_ext_RW0_rdata;
              s2_tl_error <=s1_hit&_tag_array_0_ext_RW0_rdata[20];
            end 
       end
  
  tag_array_0_64x21 tag_array_0_ext(.RW0_addr(writeEnable_0 ? refill_paddr[11:6]:_tag_rdata_T),.RW0_en(readEnable_1|writeEnable_0),.RW0_clk(clock),.RW0_wmode(refill_one_beat),.RW0_wdata({refillError,refill_paddr[31:12]}),.RW0_rdata(_tag_array_0_ext_RW0_rdata)); 
  data_arrays_512x32 data_arrays_0_0_ext(.RW0_addr(refill_one_beat ? _mem_idx_T_6|refill_cnt:io_req_bits_addr[11:3]),.RW0_en(readEnable_0|wen),.RW0_clk(clock),.RW0_wmode(refill_one_beat),.RW0_wdata(auto_master_out_d_bits_data[31:0]),.RW0_rdata(_data_arrays_0_0_ext_RW0_rdata)); 
  data_arrays_512x32 data_arrays_1_0_ext(.RW0_addr(refill_one_beat ? _mem_idx_T_6|refill_cnt:io_req_bits_addr[11:3]),.RW0_en(readEnable|writeEnable),.RW0_clk(clock),.RW0_wmode(refill_one_beat),.RW0_wdata(auto_master_out_d_bits_data[63:32]),.RW0_rdata(_data_arrays_1_0_ext_RW0_rdata)); 
  assign auto_master_out_a_valid=s2_request_refill; 
  assign auto_master_out_a_bits_address={refill_paddr[31:6],6'h0}; 
  assign io_resp_valid=s2_valid&s2_hit; 
  assign io_resp_bits_data=s2_dout_0; 
  assign io_resp_bits_ae=s2_tl_error; 
endmodule
 
module ShiftQueue (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [33:0] io_enq_bits_pc,
  input [31:0] io_enq_bits_data,
  input io_enq_bits_xcpt_pf_inst,
  input io_enq_bits_xcpt_ae_inst,
  input io_enq_bits_replay,
  input io_deq_ready,
  output io_deq_valid,
  output [33:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_data,
  output io_deq_bits_xcpt_pf_inst,
  output io_deq_bits_xcpt_gf_inst,
  output io_deq_bits_xcpt_ae_inst,
  output io_deq_bits_replay,
  output [4:0] io_mask) ; 
   reg valid_0 ;  
   reg valid_1 ;  
   reg valid_2 ;  
   reg valid_3 ;  
   reg valid_4 ;  
   reg [33:0] elts_pc_0 ;  
   reg [33:0] elts_pc_1 ;  
   reg [33:0] elts_pc_2 ;  
   reg [33:0] elts_pc_3 ;  
   reg [33:0] elts_pc_4 ;  
   reg [31:0] elts_data_0 ;  
   reg [31:0] elts_data_1 ;  
   reg [31:0] elts_data_2 ;  
   reg [31:0] elts_data_3 ;  
   reg [31:0] elts_data_4 ;  
   reg elts_xcpt_pf_inst_0 ;  
   reg elts_xcpt_pf_inst_1 ;  
   reg elts_xcpt_pf_inst_2 ;  
   reg elts_xcpt_pf_inst_3 ;  
   reg elts_xcpt_pf_inst_4 ;  
   reg elts_xcpt_gf_inst_0 ;  
   reg elts_xcpt_gf_inst_1 ;  
   reg elts_xcpt_gf_inst_2 ;  
   reg elts_xcpt_gf_inst_3 ;  
   reg elts_xcpt_gf_inst_4 ;  
   reg elts_xcpt_ae_inst_0 ;  
   reg elts_xcpt_ae_inst_1 ;  
   reg elts_xcpt_ae_inst_2 ;  
   reg elts_xcpt_ae_inst_3 ;  
   reg elts_xcpt_ae_inst_4 ;  
   reg elts_replay_0 ;  
   reg elts_replay_1 ;  
   reg elts_replay_2 ;  
   reg elts_replay_3 ;  
   reg elts_replay_4 ;  
   wire _valid_4_T_4=~valid_4&io_enq_valid ;  
   wire wen_4=io_deq_ready ? _valid_4_T_4&valid_4:_valid_4_T_4&valid_3&~valid_4 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              valid_0 <=1'h0;
              valid_1 <=1'h0;
              valid_2 <=1'h0;
              valid_3 <=1'h0;
              valid_4 <=1'h0;
            end 
          else 
            if (io_deq_ready)
               begin 
                 valid_0 <=valid_1|_valid_4_T_4&valid_0;
                 valid_1 <=valid_2|_valid_4_T_4&valid_1;
                 valid_2 <=valid_3|_valid_4_T_4&valid_2;
                 valid_3 <=valid_4|_valid_4_T_4&valid_3;
                 valid_4 <=_valid_4_T_4&valid_4;
               end 
             else 
               begin 
                 valid_0 <=_valid_4_T_4|valid_0;
                 valid_1 <=_valid_4_T_4&valid_0|valid_1;
                 valid_2 <=_valid_4_T_4&valid_1|valid_2;
                 valid_3 <=_valid_4_T_4&valid_2|valid_3;
                 valid_4 <=_valid_4_T_4&valid_3|valid_4;
               end 
         if (io_deq_ready ? valid_1|_valid_4_T_4&valid_0:_valid_4_T_4&~valid_0)
            begin 
              elts_pc_0 <=valid_1 ? elts_pc_1:io_enq_bits_pc;
              elts_data_0 <=valid_1 ? elts_data_1:io_enq_bits_data;
              elts_xcpt_pf_inst_0 <=valid_1 ? elts_xcpt_pf_inst_1:io_enq_bits_xcpt_pf_inst;
              elts_xcpt_gf_inst_0 <=valid_1&elts_xcpt_gf_inst_1;
              elts_xcpt_ae_inst_0 <=valid_1 ? elts_xcpt_ae_inst_1:io_enq_bits_xcpt_ae_inst;
              elts_replay_0 <=valid_1 ? elts_replay_1:io_enq_bits_replay;
            end 
         if (io_deq_ready ? valid_2|_valid_4_T_4&valid_1:_valid_4_T_4&valid_0&~valid_1)
            begin 
              elts_pc_1 <=valid_2 ? elts_pc_2:io_enq_bits_pc;
              elts_data_1 <=valid_2 ? elts_data_2:io_enq_bits_data;
              elts_xcpt_pf_inst_1 <=valid_2 ? elts_xcpt_pf_inst_2:io_enq_bits_xcpt_pf_inst;
              elts_xcpt_gf_inst_1 <=valid_2&elts_xcpt_gf_inst_2;
              elts_xcpt_ae_inst_1 <=valid_2 ? elts_xcpt_ae_inst_2:io_enq_bits_xcpt_ae_inst;
              elts_replay_1 <=valid_2 ? elts_replay_2:io_enq_bits_replay;
            end 
         if (io_deq_ready ? valid_3|_valid_4_T_4&valid_2:_valid_4_T_4&valid_1&~valid_2)
            begin 
              elts_pc_2 <=valid_3 ? elts_pc_3:io_enq_bits_pc;
              elts_data_2 <=valid_3 ? elts_data_3:io_enq_bits_data;
              elts_xcpt_pf_inst_2 <=valid_3 ? elts_xcpt_pf_inst_3:io_enq_bits_xcpt_pf_inst;
              elts_xcpt_gf_inst_2 <=valid_3&elts_xcpt_gf_inst_3;
              elts_xcpt_ae_inst_2 <=valid_3 ? elts_xcpt_ae_inst_3:io_enq_bits_xcpt_ae_inst;
              elts_replay_2 <=valid_3 ? elts_replay_3:io_enq_bits_replay;
            end 
         if (io_deq_ready ? valid_4|_valid_4_T_4&valid_3:_valid_4_T_4&valid_2&~valid_3)
            begin 
              elts_pc_3 <=valid_4 ? elts_pc_4:io_enq_bits_pc;
              elts_data_3 <=valid_4 ? elts_data_4:io_enq_bits_data;
              elts_xcpt_pf_inst_3 <=valid_4 ? elts_xcpt_pf_inst_4:io_enq_bits_xcpt_pf_inst;
              elts_xcpt_gf_inst_3 <=valid_4&elts_xcpt_gf_inst_4;
              elts_xcpt_ae_inst_3 <=valid_4 ? elts_xcpt_ae_inst_4:io_enq_bits_xcpt_ae_inst;
              elts_replay_3 <=valid_4 ? elts_replay_4:io_enq_bits_replay;
            end 
         if (wen_4)
            begin 
              elts_pc_4 <=io_enq_bits_pc;
              elts_data_4 <=io_enq_bits_data;
              elts_xcpt_pf_inst_4 <=io_enq_bits_xcpt_pf_inst;
              elts_xcpt_ae_inst_4 <=io_enq_bits_xcpt_ae_inst;
              elts_replay_4 <=io_enq_bits_replay;
            end 
         elts_xcpt_gf_inst_4 <=~wen_4&elts_xcpt_gf_inst_4;
       end
  
  assign io_enq_ready=~valid_4; 
  assign io_deq_valid=io_enq_valid|valid_0; 
  assign io_deq_bits_pc=valid_0 ? elts_pc_0:io_enq_bits_pc; 
  assign io_deq_bits_data=valid_0 ? elts_data_0:io_enq_bits_data; 
  assign io_deq_bits_xcpt_pf_inst=valid_0 ? elts_xcpt_pf_inst_0:io_enq_bits_xcpt_pf_inst; 
  assign io_deq_bits_xcpt_gf_inst=valid_0&elts_xcpt_gf_inst_0; 
  assign io_deq_bits_xcpt_ae_inst=valid_0 ? elts_xcpt_ae_inst_0:io_enq_bits_xcpt_ae_inst; 
  assign io_deq_bits_replay=valid_0 ? elts_replay_0:io_enq_bits_replay; 
  assign io_mask={valid_4,valid_3,valid_2,valid_1,valid_0}; 
endmodule
 
module PMPChecker_2 (
  input [1:0] io_prv,
  input io_pmp_cfg_l_0,
  input io_pmp_cfg_l_1,
  input io_pmp_cfg_l_2,
  input io_pmp_cfg_l_3,
  input io_pmp_cfg_l_4,
  input io_pmp_cfg_l_5,
  input io_pmp_cfg_l_6,
  input io_pmp_cfg_l_7,
  input [1:0] io_pmp_cfg_a_0,
  input [1:0] io_pmp_cfg_a_1,
  input [1:0] io_pmp_cfg_a_2,
  input [1:0] io_pmp_cfg_a_3,
  input [1:0] io_pmp_cfg_a_4,
  input [1:0] io_pmp_cfg_a_5,
  input [1:0] io_pmp_cfg_a_6,
  input [1:0] io_pmp_cfg_a_7,
  input io_pmp_cfg_x_0,
  input io_pmp_cfg_x_1,
  input io_pmp_cfg_x_2,
  input io_pmp_cfg_x_3,
  input io_pmp_cfg_x_4,
  input io_pmp_cfg_x_5,
  input io_pmp_cfg_x_6,
  input io_pmp_cfg_x_7,
  input [29:0] io_pmp_addr_0,
  input [29:0] io_pmp_addr_1,
  input [29:0] io_pmp_addr_2,
  input [29:0] io_pmp_addr_3,
  input [29:0] io_pmp_addr_4,
  input [29:0] io_pmp_addr_5,
  input [29:0] io_pmp_addr_6,
  input [29:0] io_pmp_addr_7,
  input [31:0] io_pmp_mask_0,
  input [31:0] io_pmp_mask_1,
  input [31:0] io_pmp_mask_2,
  input [31:0] io_pmp_mask_3,
  input [31:0] io_pmp_mask_4,
  input [31:0] io_pmp_mask_5,
  input [31:0] io_pmp_mask_6,
  input [31:0] io_pmp_mask_7,
  input [31:0] io_addr,
  output io_x) ; 
  assign io_x=(io_pmp_cfg_a_0[1] ? ((io_addr^{io_pmp_addr_0,2'h0})&~io_pmp_mask_0)==32'h0:io_pmp_cfg_a_0[0]&io_addr<{io_pmp_addr_0,2'h0}) ? io_pmp_cfg_x_0|io_prv[1]&~io_pmp_cfg_l_0:(io_pmp_cfg_a_1[1] ? ((io_addr^{io_pmp_addr_1,2'h0})&~io_pmp_mask_1)==32'h0:io_pmp_cfg_a_1[0]&io_addr>={io_pmp_addr_0,2'h0}&io_addr<{io_pmp_addr_1,2'h0}) ? io_pmp_cfg_x_1|io_prv[1]&~io_pmp_cfg_l_1:(io_pmp_cfg_a_2[1] ? ((io_addr^{io_pmp_addr_2,2'h0})&~io_pmp_mask_2)==32'h0:io_pmp_cfg_a_2[0]&io_addr>={io_pmp_addr_1,2'h0}&io_addr<{io_pmp_addr_2,2'h0}) ? io_pmp_cfg_x_2|io_prv[1]&~io_pmp_cfg_l_2:(io_pmp_cfg_a_3[1] ? ((io_addr^{io_pmp_addr_3,2'h0})&~io_pmp_mask_3)==32'h0:io_pmp_cfg_a_3[0]&io_addr>={io_pmp_addr_2,2'h0}&io_addr<{io_pmp_addr_3,2'h0}) ? io_pmp_cfg_x_3|io_prv[1]&~io_pmp_cfg_l_3:(io_pmp_cfg_a_4[1] ? ((io_addr^{io_pmp_addr_4,2'h0})&~io_pmp_mask_4)==32'h0:io_pmp_cfg_a_4[0]&io_addr>={io_pmp_addr_3,2'h0}&io_addr<{io_pmp_addr_4,2'h0}) ? io_pmp_cfg_x_4|io_prv[1]&~io_pmp_cfg_l_4:(io_pmp_cfg_a_5[1] ? ((io_addr^{io_pmp_addr_5,2'h0})&~io_pmp_mask_5)==32'h0:io_pmp_cfg_a_5[0]&io_addr>={io_pmp_addr_4,2'h0}&io_addr<{io_pmp_addr_5,2'h0}) ? io_pmp_cfg_x_5|io_prv[1]&~io_pmp_cfg_l_5:(io_pmp_cfg_a_6[1] ? ((io_addr^{io_pmp_addr_6,2'h0})&~io_pmp_mask_6)==32'h0:io_pmp_cfg_a_6[0]&io_addr>={io_pmp_addr_5,2'h0}&io_addr<{io_pmp_addr_6,2'h0}) ? io_pmp_cfg_x_6|io_prv[1]&~io_pmp_cfg_l_6:(io_pmp_cfg_a_7[1] ? ((io_addr^{io_pmp_addr_7,2'h0})&~io_pmp_mask_7)==32'h0:io_pmp_cfg_a_7[0]&io_addr>={io_pmp_addr_6,2'h0}&io_addr<{io_pmp_addr_7,2'h0}) ? io_pmp_cfg_x_7|io_prv[1]&~io_pmp_cfg_l_7:io_prv[1]; 
endmodule
 
module TLB_1 (
  input [33:0] io_req_bits_vaddr,
  output [31:0] io_resp_paddr,
  output io_resp_pf_inst,
  output io_resp_ae_inst,
  output io_resp_cacheable,
  output io_ptw_req_bits_bits_need_gpa,
  output io_ptw_req_bits_bits_stage2,
  input io_ptw_status_debug,
  input io_ptw_pmp_cfg_l_0,
  input io_ptw_pmp_cfg_l_1,
  input io_ptw_pmp_cfg_l_2,
  input io_ptw_pmp_cfg_l_3,
  input io_ptw_pmp_cfg_l_4,
  input io_ptw_pmp_cfg_l_5,
  input io_ptw_pmp_cfg_l_6,
  input io_ptw_pmp_cfg_l_7,
  input [1:0] io_ptw_pmp_cfg_a_0,
  input [1:0] io_ptw_pmp_cfg_a_1,
  input [1:0] io_ptw_pmp_cfg_a_2,
  input [1:0] io_ptw_pmp_cfg_a_3,
  input [1:0] io_ptw_pmp_cfg_a_4,
  input [1:0] io_ptw_pmp_cfg_a_5,
  input [1:0] io_ptw_pmp_cfg_a_6,
  input [1:0] io_ptw_pmp_cfg_a_7,
  input io_ptw_pmp_cfg_x_0,
  input io_ptw_pmp_cfg_x_1,
  input io_ptw_pmp_cfg_x_2,
  input io_ptw_pmp_cfg_x_3,
  input io_ptw_pmp_cfg_x_4,
  input io_ptw_pmp_cfg_x_5,
  input io_ptw_pmp_cfg_x_6,
  input io_ptw_pmp_cfg_x_7,
  input [29:0] io_ptw_pmp_addr_0,
  input [29:0] io_ptw_pmp_addr_1,
  input [29:0] io_ptw_pmp_addr_2,
  input [29:0] io_ptw_pmp_addr_3,
  input [29:0] io_ptw_pmp_addr_4,
  input [29:0] io_ptw_pmp_addr_5,
  input [29:0] io_ptw_pmp_addr_6,
  input [29:0] io_ptw_pmp_addr_7,
  input [31:0] io_ptw_pmp_mask_0,
  input [31:0] io_ptw_pmp_mask_1,
  input [31:0] io_ptw_pmp_mask_2,
  input [31:0] io_ptw_pmp_mask_3,
  input [31:0] io_ptw_pmp_mask_4,
  input [31:0] io_ptw_pmp_mask_5,
  input [31:0] io_ptw_pmp_mask_6,
  input [31:0] io_ptw_pmp_mask_7) ; 
   wire _pmp_io_x ;  
   wire [3:0] _GEN=io_req_bits_vaddr[31:28]^4'h8 ;  
   wire legal_address={io_req_bits_vaddr[33:14],~(io_req_bits_vaddr[13:12])}==22'h0|{io_req_bits_vaddr[33:28],~(io_req_bits_vaddr[27:26])}==8'h0|{io_req_bits_vaddr[33:26],io_req_bits_vaddr[25:16]^10'h200}==18'h0|~(|(io_req_bits_vaddr[33:12]))|{io_req_bits_vaddr[33:17],~(io_req_bits_vaddr[16])}==18'h0|{io_req_bits_vaddr[33:32],_GEN}==6'h0|{io_req_bits_vaddr[33:31],~(io_req_bits_vaddr[30:29])}==5'h0 ;  
  PMPChecker_2 pmp(.io_prv(2'h3),.io_pmp_cfg_l_0(io_ptw_pmp_cfg_l_0),.io_pmp_cfg_l_1(io_ptw_pmp_cfg_l_1),.io_pmp_cfg_l_2(io_ptw_pmp_cfg_l_2),.io_pmp_cfg_l_3(io_ptw_pmp_cfg_l_3),.io_pmp_cfg_l_4(io_ptw_pmp_cfg_l_4),.io_pmp_cfg_l_5(io_ptw_pmp_cfg_l_5),.io_pmp_cfg_l_6(io_ptw_pmp_cfg_l_6),.io_pmp_cfg_l_7(io_ptw_pmp_cfg_l_7),.io_pmp_cfg_a_0(io_ptw_pmp_cfg_a_0),.io_pmp_cfg_a_1(io_ptw_pmp_cfg_a_1),.io_pmp_cfg_a_2(io_ptw_pmp_cfg_a_2),.io_pmp_cfg_a_3(io_ptw_pmp_cfg_a_3),.io_pmp_cfg_a_4(io_ptw_pmp_cfg_a_4),.io_pmp_cfg_a_5(io_ptw_pmp_cfg_a_5),.io_pmp_cfg_a_6(io_ptw_pmp_cfg_a_6),.io_pmp_cfg_a_7(io_ptw_pmp_cfg_a_7),.io_pmp_cfg_x_0(io_ptw_pmp_cfg_x_0),.io_pmp_cfg_x_1(io_ptw_pmp_cfg_x_1),.io_pmp_cfg_x_2(io_ptw_pmp_cfg_x_2),.io_pmp_cfg_x_3(io_ptw_pmp_cfg_x_3),.io_pmp_cfg_x_4(io_ptw_pmp_cfg_x_4),.io_pmp_cfg_x_5(io_ptw_pmp_cfg_x_5),.io_pmp_cfg_x_6(io_ptw_pmp_cfg_x_6),.io_pmp_cfg_x_7(io_ptw_pmp_cfg_x_7),.io_pmp_addr_0(io_ptw_pmp_addr_0),.io_pmp_addr_1(io_ptw_pmp_addr_1),.io_pmp_addr_2(io_ptw_pmp_addr_2),.io_pmp_addr_3(io_ptw_pmp_addr_3),.io_pmp_addr_4(io_ptw_pmp_addr_4),.io_pmp_addr_5(io_ptw_pmp_addr_5),.io_pmp_addr_6(io_ptw_pmp_addr_6),.io_pmp_addr_7(io_ptw_pmp_addr_7),.io_pmp_mask_0(io_ptw_pmp_mask_0),.io_pmp_mask_1(io_ptw_pmp_mask_1),.io_pmp_mask_2(io_ptw_pmp_mask_2),.io_pmp_mask_3(io_ptw_pmp_mask_3),.io_pmp_mask_4(io_ptw_pmp_mask_4),.io_pmp_mask_5(io_ptw_pmp_mask_5),.io_pmp_mask_6(io_ptw_pmp_mask_6),.io_pmp_mask_7(io_ptw_pmp_mask_7),.io_addr(io_req_bits_vaddr[31:0]),.io_x(_pmp_io_x)); 
  OptimizationBarrier entries_barrier(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier entries_barrier_1(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier entries_barrier_2(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier entries_barrier_3(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier entries_barrier_4(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  OptimizationBarrier entries_barrier_5(.io_x_u(1'h0),.io_x_ae_ptw(1'h0),.io_x_ae_final(1'h0),.io_x_pf(1'h0),.io_x_gf(1'h0),.io_x_sw(1'h0),.io_x_sx(1'h0),.io_x_sr(1'h0),.io_x_pw(1'h0),.io_x_px(1'h0),.io_x_pr(1'h0),.io_x_ppp(1'h0),.io_x_pal(1'h0),.io_x_paa(1'h0),.io_x_eff(1'h0),.io_x_c(1'h0),.io_y_u(),.io_y_ae_ptw(),.io_y_ae_final(),.io_y_pf(),.io_y_gf(),.io_y_sw(),.io_y_sx(),.io_y_sr(),.io_y_pw(),.io_y_px(),.io_y_pr(),.io_y_ppp(),.io_y_pal(),.io_y_paa(),.io_y_eff(),.io_y_c()); 
  assign io_resp_paddr=io_req_bits_vaddr[31:0]; 
  assign io_resp_pf_inst=1'h0; 
  assign io_resp_ae_inst=~(legal_address&({io_req_bits_vaddr[31:30],io_req_bits_vaddr[27],io_req_bits_vaddr[25]}==4'h0|{io_req_bits_vaddr[31],~(io_req_bits_vaddr[30])}==2'h0|_GEN[3:2]==2'h0)&~(~io_ptw_status_debug&~(|(io_req_bits_vaddr[33:12])))&_pmp_io_x); 
  assign io_resp_cacheable=legal_address&~(_GEN[3]); 
  assign io_ptw_req_bits_bits_need_gpa=1'h0; 
  assign io_ptw_req_bits_bits_stage2=1'h0; 
endmodule
 
module Frontend (
  input clock,
  input reset,
  input auto_icache_master_out_a_ready,
  output auto_icache_master_out_a_valid,
  output [31:0] auto_icache_master_out_a_bits_address,
  input auto_icache_master_out_d_valid,
  input [2:0] auto_icache_master_out_d_bits_opcode,
  input [3:0] auto_icache_master_out_d_bits_size,
  input [63:0] auto_icache_master_out_d_bits_data,
  input auto_icache_master_out_d_bits_corrupt,
  input io_cpu_might_request,
  input io_cpu_req_valid,
  input [33:0] io_cpu_req_bits_pc,
  input io_cpu_req_bits_speculative,
  input io_cpu_resp_ready,
  output io_cpu_resp_valid,
  output [33:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output io_cpu_resp_bits_xcpt_pf_inst,
  output io_cpu_resp_bits_xcpt_gf_inst,
  output io_cpu_resp_bits_xcpt_ae_inst,
  output io_cpu_resp_bits_replay,
  input io_cpu_btb_update_valid,
  input io_cpu_bht_update_valid,
  input io_cpu_flush_icache,
  output io_ptw_req_bits_bits_need_gpa,
  output io_ptw_req_bits_bits_stage2,
  input io_ptw_status_debug,
  input io_ptw_pmp_cfg_l_0,
  input io_ptw_pmp_cfg_l_1,
  input io_ptw_pmp_cfg_l_2,
  input io_ptw_pmp_cfg_l_3,
  input io_ptw_pmp_cfg_l_4,
  input io_ptw_pmp_cfg_l_5,
  input io_ptw_pmp_cfg_l_6,
  input io_ptw_pmp_cfg_l_7,
  input [1:0] io_ptw_pmp_cfg_a_0,
  input [1:0] io_ptw_pmp_cfg_a_1,
  input [1:0] io_ptw_pmp_cfg_a_2,
  input [1:0] io_ptw_pmp_cfg_a_3,
  input [1:0] io_ptw_pmp_cfg_a_4,
  input [1:0] io_ptw_pmp_cfg_a_5,
  input [1:0] io_ptw_pmp_cfg_a_6,
  input [1:0] io_ptw_pmp_cfg_a_7,
  input io_ptw_pmp_cfg_x_0,
  input io_ptw_pmp_cfg_x_1,
  input io_ptw_pmp_cfg_x_2,
  input io_ptw_pmp_cfg_x_3,
  input io_ptw_pmp_cfg_x_4,
  input io_ptw_pmp_cfg_x_5,
  input io_ptw_pmp_cfg_x_6,
  input io_ptw_pmp_cfg_x_7,
  input [29:0] io_ptw_pmp_addr_0,
  input [29:0] io_ptw_pmp_addr_1,
  input [29:0] io_ptw_pmp_addr_2,
  input [29:0] io_ptw_pmp_addr_3,
  input [29:0] io_ptw_pmp_addr_4,
  input [29:0] io_ptw_pmp_addr_5,
  input [29:0] io_ptw_pmp_addr_6,
  input [29:0] io_ptw_pmp_addr_7,
  input [31:0] io_ptw_pmp_mask_0,
  input [31:0] io_ptw_pmp_mask_1,
  input [31:0] io_ptw_pmp_mask_2,
  input [31:0] io_ptw_pmp_mask_3,
  input [31:0] io_ptw_pmp_mask_4,
  input [31:0] io_ptw_pmp_mask_5,
  input [31:0] io_ptw_pmp_mask_6,
  input [31:0] io_ptw_pmp_mask_7,
  input [63:0] io_ptw_customCSRs_csrs_0_value) ; 
   wire [32:0] _io_cpu_npc_T ;  
   wire fq_io_enq_valid ;  
   wire [31:0] _tlb_io_resp_paddr ;  
   wire _tlb_io_resp_pf_inst ;  
   wire _tlb_io_resp_ae_inst ;  
   wire _tlb_io_resp_cacheable ;  
   wire _fq_io_enq_ready ;  
   wire [4:0] _fq_io_mask ;  
   wire _icache_io_resp_valid ;  
   wire [31:0] _icache_io_resp_bits_data ;  
   wire _icache_io_resp_bits_ae ;  
   reg s1_valid ;  
   reg s2_valid ;  
   wire s0_valid=io_cpu_req_valid|~(_fq_io_mask[2])|~(_fq_io_mask[3])&(~s1_valid|~s2_valid)|~(_fq_io_mask[4])&~s1_valid&~s2_valid ;  
   reg [33:0] s1_pc ;  
   reg s1_speculative ;  
   reg [33:0] s2_pc ;  
   reg s2_tlb_resp_pf_inst ;  
   reg s2_tlb_resp_ae_inst ;  
   reg s2_tlb_resp_cacheable ;  
   wire _s2_xcpt_T=s2_tlb_resp_ae_inst|s2_tlb_resp_pf_inst ;  
   reg s2_speculative ;  
   wire [33:0] predicted_npc={s1_pc[33:2],2'h0}+34'h4 ;  
   reg s2_replay_REG ;  
   wire s2_replay=s2_valid&~(_fq_io_enq_ready&fq_io_enq_valid)|s2_replay_REG ;  
   wire icache_io_s2_kill=s2_speculative&~(s2_tlb_resp_cacheable&~(io_ptw_customCSRs_csrs_0_value[3]))|_s2_xcpt_T ;  
   reg fq_io_enq_valid_REG ;  
  assign fq_io_enq_valid=fq_io_enq_valid_REG&s2_valid&(_icache_io_resp_valid|icache_io_s2_kill); 
  assign _io_cpu_npc_T=io_cpu_req_valid ? io_cpu_req_bits_pc[33:1]:s2_replay ? s2_pc[33:1]:predicted_npc[33:1]; 
  always @( posedge clock)
       begin 
         if (~reset&~(~(io_cpu_req_valid|io_cpu_flush_icache|io_cpu_bht_update_valid|io_cpu_btb_update_valid)|io_cpu_might_request))
            begin 
              if (1)$display("Assertion failed\n    at Frontend.scala:92 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n");
              if (1)$display("");
            end 
         if (~reset&s2_speculative&io_ptw_customCSRs_csrs_0_value[3]&~icache_io_s2_kill)
            begin 
              if (1)$display("Assertion failed\n    at Frontend.scala:190 assert(!(s2_speculative && io.ptw.customCSRs.asInstanceOf[RocketCustomCSRs].disableSpeculativeICacheRefill && !icache.io.s2_kill))\n");
              if (1)$display("");
            end 
       end
  
  always @( posedge clock)
       begin 
         s1_valid <=s0_valid;
         s1_pc <={_io_cpu_npc_T,1'h0};
         if (io_cpu_req_valid)
            s1_speculative <=io_cpu_req_bits_speculative;
          else 
            if (s2_replay)
               s1_speculative <=s2_speculative;
             else 
               s1_speculative <=s1_speculative|s2_valid&~s2_speculative;
         if (~s2_replay)
            begin 
              s2_tlb_resp_pf_inst <=_tlb_io_resp_pf_inst;
              s2_tlb_resp_ae_inst <=_tlb_io_resp_ae_inst;
              s2_tlb_resp_cacheable <=_tlb_io_resp_cacheable;
            end 
         fq_io_enq_valid_REG <=s1_valid;
         if (reset)
            begin 
              s2_valid <=1'h0;
              s2_pc <=34'h10040;
              s2_speculative <=1'h0;
              s2_replay_REG <=1'h1;
            end 
          else 
            begin 
              s2_valid <=~s2_replay&~io_cpu_req_valid;
              if (~s2_replay)
                 begin 
                   s2_pc <=s1_pc;
                   s2_speculative <=s1_speculative;
                 end 
              s2_replay_REG <=s2_replay&~s0_valid;
            end 
       end
  
  ICache icache(.clock(clock),.reset(reset),.auto_master_out_a_ready(auto_icache_master_out_a_ready),.auto_master_out_a_valid(auto_icache_master_out_a_valid),.auto_master_out_a_bits_address(auto_icache_master_out_a_bits_address),.auto_master_out_d_valid(auto_icache_master_out_d_valid),.auto_master_out_d_bits_opcode(auto_icache_master_out_d_bits_opcode),.auto_master_out_d_bits_size(auto_icache_master_out_d_bits_size),.auto_master_out_d_bits_data(auto_icache_master_out_d_bits_data),.auto_master_out_d_bits_corrupt(auto_icache_master_out_d_bits_corrupt),.io_req_valid(s0_valid),.io_req_bits_addr({_io_cpu_npc_T[31:0],1'h0}),.io_s1_paddr(_tlb_io_resp_paddr),.io_s1_kill(io_cpu_req_valid|s2_replay),.io_s2_kill(icache_io_s2_kill),.io_resp_valid(_icache_io_resp_valid),.io_resp_bits_data(_icache_io_resp_bits_data),.io_resp_bits_ae(_icache_io_resp_bits_ae),.io_invalidate(io_cpu_flush_icache)); 
  ShiftQueue fq(.clock(clock),.reset(reset|io_cpu_req_valid),.io_enq_ready(_fq_io_enq_ready),.io_enq_valid(fq_io_enq_valid),.io_enq_bits_pc(s2_pc),.io_enq_bits_data(_icache_io_resp_bits_data),.io_enq_bits_xcpt_pf_inst(s2_tlb_resp_pf_inst),.io_enq_bits_xcpt_ae_inst(_icache_io_resp_valid&_icache_io_resp_bits_ae|s2_tlb_resp_ae_inst),.io_enq_bits_replay(icache_io_s2_kill&~_icache_io_resp_valid&~_s2_xcpt_T),.io_deq_ready(io_cpu_resp_ready),.io_deq_valid(io_cpu_resp_valid),.io_deq_bits_pc(io_cpu_resp_bits_pc),.io_deq_bits_data(io_cpu_resp_bits_data),.io_deq_bits_xcpt_pf_inst(io_cpu_resp_bits_xcpt_pf_inst),.io_deq_bits_xcpt_gf_inst(io_cpu_resp_bits_xcpt_gf_inst),.io_deq_bits_xcpt_ae_inst(io_cpu_resp_bits_xcpt_ae_inst),.io_deq_bits_replay(io_cpu_resp_bits_replay),.io_mask(_fq_io_mask)); 
  TLB_1 tlb(.io_req_bits_vaddr(s1_pc),.io_resp_paddr(_tlb_io_resp_paddr),.io_resp_pf_inst(_tlb_io_resp_pf_inst),.io_resp_ae_inst(_tlb_io_resp_ae_inst),.io_resp_cacheable(_tlb_io_resp_cacheable),.io_ptw_req_bits_bits_need_gpa(io_ptw_req_bits_bits_need_gpa),.io_ptw_req_bits_bits_stage2(io_ptw_req_bits_bits_stage2),.io_ptw_status_debug(io_ptw_status_debug),.io_ptw_pmp_cfg_l_0(io_ptw_pmp_cfg_l_0),.io_ptw_pmp_cfg_l_1(io_ptw_pmp_cfg_l_1),.io_ptw_pmp_cfg_l_2(io_ptw_pmp_cfg_l_2),.io_ptw_pmp_cfg_l_3(io_ptw_pmp_cfg_l_3),.io_ptw_pmp_cfg_l_4(io_ptw_pmp_cfg_l_4),.io_ptw_pmp_cfg_l_5(io_ptw_pmp_cfg_l_5),.io_ptw_pmp_cfg_l_6(io_ptw_pmp_cfg_l_6),.io_ptw_pmp_cfg_l_7(io_ptw_pmp_cfg_l_7),.io_ptw_pmp_cfg_a_0(io_ptw_pmp_cfg_a_0),.io_ptw_pmp_cfg_a_1(io_ptw_pmp_cfg_a_1),.io_ptw_pmp_cfg_a_2(io_ptw_pmp_cfg_a_2),.io_ptw_pmp_cfg_a_3(io_ptw_pmp_cfg_a_3),.io_ptw_pmp_cfg_a_4(io_ptw_pmp_cfg_a_4),.io_ptw_pmp_cfg_a_5(io_ptw_pmp_cfg_a_5),.io_ptw_pmp_cfg_a_6(io_ptw_pmp_cfg_a_6),.io_ptw_pmp_cfg_a_7(io_ptw_pmp_cfg_a_7),.io_ptw_pmp_cfg_x_0(io_ptw_pmp_cfg_x_0),.io_ptw_pmp_cfg_x_1(io_ptw_pmp_cfg_x_1),.io_ptw_pmp_cfg_x_2(io_ptw_pmp_cfg_x_2),.io_ptw_pmp_cfg_x_3(io_ptw_pmp_cfg_x_3),.io_ptw_pmp_cfg_x_4(io_ptw_pmp_cfg_x_4),.io_ptw_pmp_cfg_x_5(io_ptw_pmp_cfg_x_5),.io_ptw_pmp_cfg_x_6(io_ptw_pmp_cfg_x_6),.io_ptw_pmp_cfg_x_7(io_ptw_pmp_cfg_x_7),.io_ptw_pmp_addr_0(io_ptw_pmp_addr_0),.io_ptw_pmp_addr_1(io_ptw_pmp_addr_1),.io_ptw_pmp_addr_2(io_ptw_pmp_addr_2),.io_ptw_pmp_addr_3(io_ptw_pmp_addr_3),.io_ptw_pmp_addr_4(io_ptw_pmp_addr_4),.io_ptw_pmp_addr_5(io_ptw_pmp_addr_5),.io_ptw_pmp_addr_6(io_ptw_pmp_addr_6),.io_ptw_pmp_addr_7(io_ptw_pmp_addr_7),.io_ptw_pmp_mask_0(io_ptw_pmp_mask_0),.io_ptw_pmp_mask_1(io_ptw_pmp_mask_1),.io_ptw_pmp_mask_2(io_ptw_pmp_mask_2),.io_ptw_pmp_mask_3(io_ptw_pmp_mask_3),.io_ptw_pmp_mask_4(io_ptw_pmp_mask_4),.io_ptw_pmp_mask_5(io_ptw_pmp_mask_5),.io_ptw_pmp_mask_6(io_ptw_pmp_mask_6),.io_ptw_pmp_mask_7(io_ptw_pmp_mask_7)); 
endmodule
 
module HellaCacheArbiter (
  output io_requestor_0_req_ready,
  input io_requestor_0_req_valid,
  input [33:0] io_requestor_0_req_bits_addr,
  input [5:0] io_requestor_0_req_bits_tag,
  input [4:0] io_requestor_0_req_bits_cmd,
  input [1:0] io_requestor_0_req_bits_size,
  input io_requestor_0_req_bits_signed,
  input io_requestor_0_req_bits_dv,
  input io_requestor_0_s1_kill,
  input [63:0] io_requestor_0_s1_data_data,
  output io_requestor_0_s2_nack,
  output io_requestor_0_resp_valid,
  output [5:0] io_requestor_0_resp_bits_tag,
  output [63:0] io_requestor_0_resp_bits_data,
  output io_requestor_0_resp_bits_replay,
  output io_requestor_0_resp_bits_has_data,
  output [63:0] io_requestor_0_resp_bits_data_word_bypass,
  output io_requestor_0_replay_next,
  output io_requestor_0_s2_xcpt_ma_ld,
  output io_requestor_0_s2_xcpt_ma_st,
  output io_requestor_0_s2_xcpt_pf_ld,
  output io_requestor_0_s2_xcpt_pf_st,
  output io_requestor_0_s2_xcpt_ae_ld,
  output io_requestor_0_s2_xcpt_ae_st,
  output io_requestor_0_ordered,
  output io_requestor_0_perf_release,
  output io_requestor_0_perf_grant,
  input io_mem_req_ready,
  output io_mem_req_valid,
  output [33:0] io_mem_req_bits_addr,
  output [5:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [1:0] io_mem_req_bits_size,
  output io_mem_req_bits_signed,
  output io_mem_req_bits_dv,
  output io_mem_s1_kill,
  output [63:0] io_mem_s1_data_data,
  input io_mem_s2_nack,
  input io_mem_resp_valid,
  input [5:0] io_mem_resp_bits_tag,
  input [63:0] io_mem_resp_bits_data,
  input io_mem_resp_bits_replay,
  input io_mem_resp_bits_has_data,
  input [63:0] io_mem_resp_bits_data_word_bypass,
  input io_mem_replay_next,
  input io_mem_s2_xcpt_ma_ld,
  input io_mem_s2_xcpt_ma_st,
  input io_mem_s2_xcpt_pf_ld,
  input io_mem_s2_xcpt_pf_st,
  input io_mem_s2_xcpt_ae_ld,
  input io_mem_s2_xcpt_ae_st,
  input io_mem_ordered,
  input io_mem_perf_release,
  input io_mem_perf_grant) ; 
  assign io_requestor_0_req_ready=io_mem_req_ready; 
  assign io_requestor_0_s2_nack=io_mem_s2_nack; 
  assign io_requestor_0_resp_valid=io_mem_resp_valid; 
  assign io_requestor_0_resp_bits_tag=io_mem_resp_bits_tag; 
  assign io_requestor_0_resp_bits_data=io_mem_resp_bits_data; 
  assign io_requestor_0_resp_bits_replay=io_mem_resp_bits_replay; 
  assign io_requestor_0_resp_bits_has_data=io_mem_resp_bits_has_data; 
  assign io_requestor_0_resp_bits_data_word_bypass=io_mem_resp_bits_data_word_bypass; 
  assign io_requestor_0_replay_next=io_mem_replay_next; 
  assign io_requestor_0_s2_xcpt_ma_ld=io_mem_s2_xcpt_ma_ld; 
  assign io_requestor_0_s2_xcpt_ma_st=io_mem_s2_xcpt_ma_st; 
  assign io_requestor_0_s2_xcpt_pf_ld=io_mem_s2_xcpt_pf_ld; 
  assign io_requestor_0_s2_xcpt_pf_st=io_mem_s2_xcpt_pf_st; 
  assign io_requestor_0_s2_xcpt_ae_ld=io_mem_s2_xcpt_ae_ld; 
  assign io_requestor_0_s2_xcpt_ae_st=io_mem_s2_xcpt_ae_st; 
  assign io_requestor_0_ordered=io_mem_ordered; 
  assign io_requestor_0_perf_release=io_mem_perf_release; 
  assign io_requestor_0_perf_grant=io_mem_perf_grant; 
  assign io_mem_req_valid=io_requestor_0_req_valid; 
  assign io_mem_req_bits_addr=io_requestor_0_req_bits_addr; 
  assign io_mem_req_bits_tag=io_requestor_0_req_bits_tag; 
  assign io_mem_req_bits_cmd=io_requestor_0_req_bits_cmd; 
  assign io_mem_req_bits_size=io_requestor_0_req_bits_size; 
  assign io_mem_req_bits_signed=io_requestor_0_req_bits_signed; 
  assign io_mem_req_bits_dv=io_requestor_0_req_bits_dv; 
  assign io_mem_s1_kill=io_requestor_0_s1_kill; 
  assign io_mem_s1_data_data=io_requestor_0_s1_data_data; 
endmodule
 
module Arbiter (
  input io_in_0_bits_bits_need_gpa,
  input io_in_0_bits_bits_stage2,
  input io_in_1_bits_bits_need_gpa,
  input io_in_1_bits_bits_stage2,
  output io_out_bits_bits_need_gpa,
  output io_out_bits_bits_stage2) ; 
  assign io_out_bits_bits_need_gpa=io_in_1_bits_bits_need_gpa; 
  assign io_out_bits_bits_stage2=io_in_1_bits_bits_stage2; 
endmodule
 
module PTW (
  input clock,
  input io_requestor_0_req_bits_bits_need_gpa,
  input io_requestor_0_req_bits_bits_stage2,
  output io_requestor_0_status_debug,
  output io_requestor_0_pmp_cfg_l_0,
  output io_requestor_0_pmp_cfg_l_1,
  output io_requestor_0_pmp_cfg_l_2,
  output io_requestor_0_pmp_cfg_l_3,
  output io_requestor_0_pmp_cfg_l_4,
  output io_requestor_0_pmp_cfg_l_5,
  output io_requestor_0_pmp_cfg_l_6,
  output io_requestor_0_pmp_cfg_l_7,
  output [1:0] io_requestor_0_pmp_cfg_a_0,
  output [1:0] io_requestor_0_pmp_cfg_a_1,
  output [1:0] io_requestor_0_pmp_cfg_a_2,
  output [1:0] io_requestor_0_pmp_cfg_a_3,
  output [1:0] io_requestor_0_pmp_cfg_a_4,
  output [1:0] io_requestor_0_pmp_cfg_a_5,
  output [1:0] io_requestor_0_pmp_cfg_a_6,
  output [1:0] io_requestor_0_pmp_cfg_a_7,
  output io_requestor_0_pmp_cfg_w_0,
  output io_requestor_0_pmp_cfg_w_1,
  output io_requestor_0_pmp_cfg_w_2,
  output io_requestor_0_pmp_cfg_w_3,
  output io_requestor_0_pmp_cfg_w_4,
  output io_requestor_0_pmp_cfg_w_5,
  output io_requestor_0_pmp_cfg_w_6,
  output io_requestor_0_pmp_cfg_w_7,
  output io_requestor_0_pmp_cfg_r_0,
  output io_requestor_0_pmp_cfg_r_1,
  output io_requestor_0_pmp_cfg_r_2,
  output io_requestor_0_pmp_cfg_r_3,
  output io_requestor_0_pmp_cfg_r_4,
  output io_requestor_0_pmp_cfg_r_5,
  output io_requestor_0_pmp_cfg_r_6,
  output io_requestor_0_pmp_cfg_r_7,
  output [29:0] io_requestor_0_pmp_addr_0,
  output [29:0] io_requestor_0_pmp_addr_1,
  output [29:0] io_requestor_0_pmp_addr_2,
  output [29:0] io_requestor_0_pmp_addr_3,
  output [29:0] io_requestor_0_pmp_addr_4,
  output [29:0] io_requestor_0_pmp_addr_5,
  output [29:0] io_requestor_0_pmp_addr_6,
  output [29:0] io_requestor_0_pmp_addr_7,
  output [31:0] io_requestor_0_pmp_mask_0,
  output [31:0] io_requestor_0_pmp_mask_1,
  output [31:0] io_requestor_0_pmp_mask_2,
  output [31:0] io_requestor_0_pmp_mask_3,
  output [31:0] io_requestor_0_pmp_mask_4,
  output [31:0] io_requestor_0_pmp_mask_5,
  output [31:0] io_requestor_0_pmp_mask_6,
  output [31:0] io_requestor_0_pmp_mask_7,
  input io_requestor_1_req_bits_bits_need_gpa,
  input io_requestor_1_req_bits_bits_stage2,
  output io_requestor_1_status_debug,
  output io_requestor_1_pmp_cfg_l_0,
  output io_requestor_1_pmp_cfg_l_1,
  output io_requestor_1_pmp_cfg_l_2,
  output io_requestor_1_pmp_cfg_l_3,
  output io_requestor_1_pmp_cfg_l_4,
  output io_requestor_1_pmp_cfg_l_5,
  output io_requestor_1_pmp_cfg_l_6,
  output io_requestor_1_pmp_cfg_l_7,
  output [1:0] io_requestor_1_pmp_cfg_a_0,
  output [1:0] io_requestor_1_pmp_cfg_a_1,
  output [1:0] io_requestor_1_pmp_cfg_a_2,
  output [1:0] io_requestor_1_pmp_cfg_a_3,
  output [1:0] io_requestor_1_pmp_cfg_a_4,
  output [1:0] io_requestor_1_pmp_cfg_a_5,
  output [1:0] io_requestor_1_pmp_cfg_a_6,
  output [1:0] io_requestor_1_pmp_cfg_a_7,
  output io_requestor_1_pmp_cfg_x_0,
  output io_requestor_1_pmp_cfg_x_1,
  output io_requestor_1_pmp_cfg_x_2,
  output io_requestor_1_pmp_cfg_x_3,
  output io_requestor_1_pmp_cfg_x_4,
  output io_requestor_1_pmp_cfg_x_5,
  output io_requestor_1_pmp_cfg_x_6,
  output io_requestor_1_pmp_cfg_x_7,
  output [29:0] io_requestor_1_pmp_addr_0,
  output [29:0] io_requestor_1_pmp_addr_1,
  output [29:0] io_requestor_1_pmp_addr_2,
  output [29:0] io_requestor_1_pmp_addr_3,
  output [29:0] io_requestor_1_pmp_addr_4,
  output [29:0] io_requestor_1_pmp_addr_5,
  output [29:0] io_requestor_1_pmp_addr_6,
  output [29:0] io_requestor_1_pmp_addr_7,
  output [31:0] io_requestor_1_pmp_mask_0,
  output [31:0] io_requestor_1_pmp_mask_1,
  output [31:0] io_requestor_1_pmp_mask_2,
  output [31:0] io_requestor_1_pmp_mask_3,
  output [31:0] io_requestor_1_pmp_mask_4,
  output [31:0] io_requestor_1_pmp_mask_5,
  output [31:0] io_requestor_1_pmp_mask_6,
  output [31:0] io_requestor_1_pmp_mask_7,
  output [63:0] io_requestor_1_customCSRs_csrs_0_value,
  input io_dpath_status_debug,
  input io_dpath_pmp_cfg_l_0,
  input io_dpath_pmp_cfg_l_1,
  input io_dpath_pmp_cfg_l_2,
  input io_dpath_pmp_cfg_l_3,
  input io_dpath_pmp_cfg_l_4,
  input io_dpath_pmp_cfg_l_5,
  input io_dpath_pmp_cfg_l_6,
  input io_dpath_pmp_cfg_l_7,
  input [1:0] io_dpath_pmp_cfg_a_0,
  input [1:0] io_dpath_pmp_cfg_a_1,
  input [1:0] io_dpath_pmp_cfg_a_2,
  input [1:0] io_dpath_pmp_cfg_a_3,
  input [1:0] io_dpath_pmp_cfg_a_4,
  input [1:0] io_dpath_pmp_cfg_a_5,
  input [1:0] io_dpath_pmp_cfg_a_6,
  input [1:0] io_dpath_pmp_cfg_a_7,
  input io_dpath_pmp_cfg_x_0,
  input io_dpath_pmp_cfg_x_1,
  input io_dpath_pmp_cfg_x_2,
  input io_dpath_pmp_cfg_x_3,
  input io_dpath_pmp_cfg_x_4,
  input io_dpath_pmp_cfg_x_5,
  input io_dpath_pmp_cfg_x_6,
  input io_dpath_pmp_cfg_x_7,
  input io_dpath_pmp_cfg_w_0,
  input io_dpath_pmp_cfg_w_1,
  input io_dpath_pmp_cfg_w_2,
  input io_dpath_pmp_cfg_w_3,
  input io_dpath_pmp_cfg_w_4,
  input io_dpath_pmp_cfg_w_5,
  input io_dpath_pmp_cfg_w_6,
  input io_dpath_pmp_cfg_w_7,
  input io_dpath_pmp_cfg_r_0,
  input io_dpath_pmp_cfg_r_1,
  input io_dpath_pmp_cfg_r_2,
  input io_dpath_pmp_cfg_r_3,
  input io_dpath_pmp_cfg_r_4,
  input io_dpath_pmp_cfg_r_5,
  input io_dpath_pmp_cfg_r_6,
  input io_dpath_pmp_cfg_r_7,
  input [29:0] io_dpath_pmp_addr_0,
  input [29:0] io_dpath_pmp_addr_1,
  input [29:0] io_dpath_pmp_addr_2,
  input [29:0] io_dpath_pmp_addr_3,
  input [29:0] io_dpath_pmp_addr_4,
  input [29:0] io_dpath_pmp_addr_5,
  input [29:0] io_dpath_pmp_addr_6,
  input [29:0] io_dpath_pmp_addr_7,
  input [31:0] io_dpath_pmp_mask_0,
  input [31:0] io_dpath_pmp_mask_1,
  input [31:0] io_dpath_pmp_mask_2,
  input [31:0] io_dpath_pmp_mask_3,
  input [31:0] io_dpath_pmp_mask_4,
  input [31:0] io_dpath_pmp_mask_5,
  input [31:0] io_dpath_pmp_mask_6,
  input [31:0] io_dpath_pmp_mask_7,
  input [63:0] io_dpath_customCSRs_csrs_0_value) ; 
  Arbiter arb(.io_in_0_bits_bits_need_gpa(io_requestor_0_req_bits_bits_need_gpa),.io_in_0_bits_bits_stage2(io_requestor_0_req_bits_bits_stage2),.io_in_1_bits_bits_need_gpa(io_requestor_1_req_bits_bits_need_gpa),.io_in_1_bits_bits_stage2(io_requestor_1_req_bits_bits_stage2),.io_out_bits_bits_need_gpa(),.io_out_bits_bits_stage2()); 
  assign io_requestor_0_status_debug=io_dpath_status_debug; 
  assign io_requestor_0_pmp_cfg_l_0=io_dpath_pmp_cfg_l_0; 
  assign io_requestor_0_pmp_cfg_l_1=io_dpath_pmp_cfg_l_1; 
  assign io_requestor_0_pmp_cfg_l_2=io_dpath_pmp_cfg_l_2; 
  assign io_requestor_0_pmp_cfg_l_3=io_dpath_pmp_cfg_l_3; 
  assign io_requestor_0_pmp_cfg_l_4=io_dpath_pmp_cfg_l_4; 
  assign io_requestor_0_pmp_cfg_l_5=io_dpath_pmp_cfg_l_5; 
  assign io_requestor_0_pmp_cfg_l_6=io_dpath_pmp_cfg_l_6; 
  assign io_requestor_0_pmp_cfg_l_7=io_dpath_pmp_cfg_l_7; 
  assign io_requestor_0_pmp_cfg_a_0=io_dpath_pmp_cfg_a_0; 
  assign io_requestor_0_pmp_cfg_a_1=io_dpath_pmp_cfg_a_1; 
  assign io_requestor_0_pmp_cfg_a_2=io_dpath_pmp_cfg_a_2; 
  assign io_requestor_0_pmp_cfg_a_3=io_dpath_pmp_cfg_a_3; 
  assign io_requestor_0_pmp_cfg_a_4=io_dpath_pmp_cfg_a_4; 
  assign io_requestor_0_pmp_cfg_a_5=io_dpath_pmp_cfg_a_5; 
  assign io_requestor_0_pmp_cfg_a_6=io_dpath_pmp_cfg_a_6; 
  assign io_requestor_0_pmp_cfg_a_7=io_dpath_pmp_cfg_a_7; 
  assign io_requestor_0_pmp_cfg_w_0=io_dpath_pmp_cfg_w_0; 
  assign io_requestor_0_pmp_cfg_w_1=io_dpath_pmp_cfg_w_1; 
  assign io_requestor_0_pmp_cfg_w_2=io_dpath_pmp_cfg_w_2; 
  assign io_requestor_0_pmp_cfg_w_3=io_dpath_pmp_cfg_w_3; 
  assign io_requestor_0_pmp_cfg_w_4=io_dpath_pmp_cfg_w_4; 
  assign io_requestor_0_pmp_cfg_w_5=io_dpath_pmp_cfg_w_5; 
  assign io_requestor_0_pmp_cfg_w_6=io_dpath_pmp_cfg_w_6; 
  assign io_requestor_0_pmp_cfg_w_7=io_dpath_pmp_cfg_w_7; 
  assign io_requestor_0_pmp_cfg_r_0=io_dpath_pmp_cfg_r_0; 
  assign io_requestor_0_pmp_cfg_r_1=io_dpath_pmp_cfg_r_1; 
  assign io_requestor_0_pmp_cfg_r_2=io_dpath_pmp_cfg_r_2; 
  assign io_requestor_0_pmp_cfg_r_3=io_dpath_pmp_cfg_r_3; 
  assign io_requestor_0_pmp_cfg_r_4=io_dpath_pmp_cfg_r_4; 
  assign io_requestor_0_pmp_cfg_r_5=io_dpath_pmp_cfg_r_5; 
  assign io_requestor_0_pmp_cfg_r_6=io_dpath_pmp_cfg_r_6; 
  assign io_requestor_0_pmp_cfg_r_7=io_dpath_pmp_cfg_r_7; 
  assign io_requestor_0_pmp_addr_0=io_dpath_pmp_addr_0; 
  assign io_requestor_0_pmp_addr_1=io_dpath_pmp_addr_1; 
  assign io_requestor_0_pmp_addr_2=io_dpath_pmp_addr_2; 
  assign io_requestor_0_pmp_addr_3=io_dpath_pmp_addr_3; 
  assign io_requestor_0_pmp_addr_4=io_dpath_pmp_addr_4; 
  assign io_requestor_0_pmp_addr_5=io_dpath_pmp_addr_5; 
  assign io_requestor_0_pmp_addr_6=io_dpath_pmp_addr_6; 
  assign io_requestor_0_pmp_addr_7=io_dpath_pmp_addr_7; 
  assign io_requestor_0_pmp_mask_0=io_dpath_pmp_mask_0; 
  assign io_requestor_0_pmp_mask_1=io_dpath_pmp_mask_1; 
  assign io_requestor_0_pmp_mask_2=io_dpath_pmp_mask_2; 
  assign io_requestor_0_pmp_mask_3=io_dpath_pmp_mask_3; 
  assign io_requestor_0_pmp_mask_4=io_dpath_pmp_mask_4; 
  assign io_requestor_0_pmp_mask_5=io_dpath_pmp_mask_5; 
  assign io_requestor_0_pmp_mask_6=io_dpath_pmp_mask_6; 
  assign io_requestor_0_pmp_mask_7=io_dpath_pmp_mask_7; 
  assign io_requestor_1_status_debug=io_dpath_status_debug; 
  assign io_requestor_1_pmp_cfg_l_0=io_dpath_pmp_cfg_l_0; 
  assign io_requestor_1_pmp_cfg_l_1=io_dpath_pmp_cfg_l_1; 
  assign io_requestor_1_pmp_cfg_l_2=io_dpath_pmp_cfg_l_2; 
  assign io_requestor_1_pmp_cfg_l_3=io_dpath_pmp_cfg_l_3; 
  assign io_requestor_1_pmp_cfg_l_4=io_dpath_pmp_cfg_l_4; 
  assign io_requestor_1_pmp_cfg_l_5=io_dpath_pmp_cfg_l_5; 
  assign io_requestor_1_pmp_cfg_l_6=io_dpath_pmp_cfg_l_6; 
  assign io_requestor_1_pmp_cfg_l_7=io_dpath_pmp_cfg_l_7; 
  assign io_requestor_1_pmp_cfg_a_0=io_dpath_pmp_cfg_a_0; 
  assign io_requestor_1_pmp_cfg_a_1=io_dpath_pmp_cfg_a_1; 
  assign io_requestor_1_pmp_cfg_a_2=io_dpath_pmp_cfg_a_2; 
  assign io_requestor_1_pmp_cfg_a_3=io_dpath_pmp_cfg_a_3; 
  assign io_requestor_1_pmp_cfg_a_4=io_dpath_pmp_cfg_a_4; 
  assign io_requestor_1_pmp_cfg_a_5=io_dpath_pmp_cfg_a_5; 
  assign io_requestor_1_pmp_cfg_a_6=io_dpath_pmp_cfg_a_6; 
  assign io_requestor_1_pmp_cfg_a_7=io_dpath_pmp_cfg_a_7; 
  assign io_requestor_1_pmp_cfg_x_0=io_dpath_pmp_cfg_x_0; 
  assign io_requestor_1_pmp_cfg_x_1=io_dpath_pmp_cfg_x_1; 
  assign io_requestor_1_pmp_cfg_x_2=io_dpath_pmp_cfg_x_2; 
  assign io_requestor_1_pmp_cfg_x_3=io_dpath_pmp_cfg_x_3; 
  assign io_requestor_1_pmp_cfg_x_4=io_dpath_pmp_cfg_x_4; 
  assign io_requestor_1_pmp_cfg_x_5=io_dpath_pmp_cfg_x_5; 
  assign io_requestor_1_pmp_cfg_x_6=io_dpath_pmp_cfg_x_6; 
  assign io_requestor_1_pmp_cfg_x_7=io_dpath_pmp_cfg_x_7; 
  assign io_requestor_1_pmp_addr_0=io_dpath_pmp_addr_0; 
  assign io_requestor_1_pmp_addr_1=io_dpath_pmp_addr_1; 
  assign io_requestor_1_pmp_addr_2=io_dpath_pmp_addr_2; 
  assign io_requestor_1_pmp_addr_3=io_dpath_pmp_addr_3; 
  assign io_requestor_1_pmp_addr_4=io_dpath_pmp_addr_4; 
  assign io_requestor_1_pmp_addr_5=io_dpath_pmp_addr_5; 
  assign io_requestor_1_pmp_addr_6=io_dpath_pmp_addr_6; 
  assign io_requestor_1_pmp_addr_7=io_dpath_pmp_addr_7; 
  assign io_requestor_1_pmp_mask_0=io_dpath_pmp_mask_0; 
  assign io_requestor_1_pmp_mask_1=io_dpath_pmp_mask_1; 
  assign io_requestor_1_pmp_mask_2=io_dpath_pmp_mask_2; 
  assign io_requestor_1_pmp_mask_3=io_dpath_pmp_mask_3; 
  assign io_requestor_1_pmp_mask_4=io_dpath_pmp_mask_4; 
  assign io_requestor_1_pmp_mask_5=io_dpath_pmp_mask_5; 
  assign io_requestor_1_pmp_mask_6=io_dpath_pmp_mask_6; 
  assign io_requestor_1_pmp_mask_7=io_dpath_pmp_mask_7; 
  assign io_requestor_1_customCSRs_csrs_0_value=io_dpath_customCSRs_csrs_0_value; 
endmodule
 
module RVCExpander (
  input [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0] io_out_rd,
  output [4:0] io_out_rs1,
  output [4:0] io_out_rs2,
  output io_rvc) ; 
   reg [2:0] casez_tmp ;  
   wire [2:0] _io_out_s_funct_T_2={io_in[12],io_in[6:5]} ;  
   wire [2:0] _io_out_s_funct_T_4={_io_out_s_funct_T_2==3'h1,2'h0} ;  
  always @(*)
       begin 
         casez (_io_out_s_funct_T_2)
          3 'b000:
             casez_tmp =_io_out_s_funct_T_4;
          3 'b001:
             casez_tmp =_io_out_s_funct_T_4;
          3 'b010:
             casez_tmp =3'h6;
          3 'b011:
             casez_tmp =3'h7;
          3 'b100:
             casez_tmp =3'h0;
          3 'b101:
             casez_tmp =3'h0;
          3 'b110:
             casez_tmp =3'h2;
          default :
             casez_tmp =3'h3;
         endcase 
       end
  
   wire [3:0] _GEN={4{io_in[12]}} ;  
   wire [6:0] io_out_s_load_opc=(|(io_in[11:7])) ? 7'h3:7'h1F ;  
   wire [4:0] _io_out_T_2={io_in[1:0],io_in[15:13]} ;  
   wire _io_out_T_29=_io_out_T_2==5'hE ;  
   wire _io_out_T_31=_io_out_T_2==5'hF ;  
   wire _io_out_T_33=_io_out_T_2==5'h10 ;  
   wire _io_out_T_35=_io_out_T_2==5'h11 ;  
   wire _io_out_T_37=_io_out_T_2==5'h12 ;  
   wire _io_out_T_39=_io_out_T_2==5'h13 ;  
   wire _io_out_T_41=_io_out_T_2==5'h14 ;  
   wire [31:0] _io_out_T_42_bits=_io_out_T_41 ? {7'h0,io_in[12] ? ((|(io_in[6:2])) ? {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}:(|(io_in[11:7])) ? {io_in[6:2],io_in[11:7],15'hE7}:{io_in[6:3],1'h1,io_in[11:7],15'h73}):{io_in[6:2],(|(io_in[6:2])) ? {8'h0,io_in[11:7],7'h33}:{io_in[11:7],(|(io_in[11:7])) ? 15'h67:15'h1F}}}:_io_out_T_39 ? {3'h0,io_in[4:2],io_in[12],io_in[6:5],11'h13,io_in[11:7],io_out_s_load_opc}:_io_out_T_37 ? {4'h0,io_in[3:2],io_in[12],io_in[6:4],10'h12,io_in[11:7],io_out_s_load_opc}:_io_out_T_35 ? {3'h0,io_in[4:2],io_in[12],io_in[6:5],11'h13,io_in[11:7],7'h7}:_io_out_T_33 ? {6'h0,io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}:_io_out_T_31 ? {_GEN,io_in[6:5],io_in[2],7'h1,io_in[9:7],3'h1,io_in[11:10],io_in[4:3],io_in[12],7'h63}:_io_out_T_29 ? {_GEN,io_in[6:5],io_in[2],7'h1,io_in[9:7],3'h0,io_in[11:10],io_in[4:3],io_in[12],7'h63}:_io_out_T_2==5'hD ? {io_in[12],io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],{9{io_in[12]}},12'h6F}:_io_out_T_2==5'hC ? ((&(io_in[11:10])) ? {1'h0,io_in[6:5]==2'h0,7'h1,io_in[4:2],2'h1,io_in[9:7],casez_tmp,2'h1,io_in[9:7],3'h3,io_in[12],3'h3}:{io_in[11:10]==2'h2 ? {{7{io_in[12]}},io_in[6:2],2'h1,io_in[9:7],5'h1D}:{1'h0,io_in[11:10]==2'h1,4'h0,io_in[12],io_in[6:2],2'h1,io_in[9:7],5'h15},io_in[9:7],7'h13}):_io_out_T_2==5'hB ? {{3{io_in[12]}},io_in[11:7]==5'h0|io_in[11:7]==5'h2 ? {io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:7],(|{{7{io_in[12]}},io_in[6:2]}) ? 7'h13:7'h1F}:{{12{io_in[12]}},io_in[6:2],io_in[11:7],3'h3,{{7{io_in[12]}},io_in[6:2]}==12'h0,3'h7}}:_io_out_T_2==5'hA ? {{7{io_in[12]}},io_in[6:2],8'h0,io_in[11:7],7'h13}:_io_out_T_2==5'h9 ? {{7{io_in[12]}},io_in[6:2],io_in[11:7],3'h0,io_in[11:7],4'h3,io_in[11:7]==5'h0,2'h3}:_io_out_T_2==5'h8 ? {{7{io_in[12]}},io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}:_io_out_T_2==5'h7 ? {4'h0,io_in[6:5],io_in[12],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,io_in[11:10],10'h23}:_io_out_T_2==5'h6 ? {5'h0,io_in[5],io_in[12],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,io_in[11:10],io_in[6],9'h23}:_io_out_T_2==5'h5 ? {4'h0,io_in[6:5],io_in[12],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,io_in[11:10],10'h27}:_io_out_T_2==5'h4 ? {5'h0,io_in[5],io_in[12],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,io_in[11:10],io_in[6],9'h3F}:_io_out_T_2==5'h3 ? {4'h0,io_in[6:5],io_in[12:10],5'h1,io_in[9:7],5'hD,io_in[4:2],7'h3}:_io_out_T_2==5'h2 ? {5'h0,io_in[5],io_in[12:10],io_in[6],4'h1,io_in[9:7],5'h9,io_in[4:2],7'h3}:_io_out_T_2==5'h1 ? {4'h0,io_in[6:5],io_in[12:10],5'h1,io_in[9:7],5'hD,io_in[4:2],7'h7}:{2'h0,io_in[10:7],io_in[12:11],io_in[5],io_in[6],12'h41,io_in[4:2],(|(io_in[12:5])) ? 7'h13:7'h1F} ;  
   wire _io_out_T_43=_io_out_T_2==5'h15 ;  
   wire _io_out_T_45=_io_out_T_2==5'h16 ;  
   wire _io_out_T_47=_io_out_T_2==5'h17 ;  
   wire _io_out_T_49=_io_out_T_2==5'h18 ;  
   wire _io_out_T_51=_io_out_T_2==5'h19 ;  
   wire _io_out_T_53=_io_out_T_2==5'h1A ;  
   wire _io_out_T_55=_io_out_T_2==5'h1B ;  
   wire _io_out_T_57=_io_out_T_2==5'h1C ;  
   wire _io_out_T_59=_io_out_T_2==5'h1D ;  
   wire _io_out_T_61=_io_out_T_2==5'h1E ;  
   reg [4:0] casez_tmp_0 ;  
   wire [4:0] io_out_s_7_rd={2'h1,io_in[4:2]} ;  
  always @(*)
       begin 
         casez (_io_out_T_2)
          5 'b00000:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b00001:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b00010:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b00011:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b00100:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b00101:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b00110:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b00111:
             casez_tmp_0 =io_out_s_7_rd;
          5 'b01000:
             casez_tmp_0 =io_in[11:7];
          5 'b01001:
             casez_tmp_0 =io_in[11:7];
          5 'b01010:
             casez_tmp_0 =io_in[11:7];
          5 'b01011:
             casez_tmp_0 =io_in[11:7];
          5 'b01100:
             casez_tmp_0 ={2'h1,io_in[9:7]};
          5 'b01101:
             casez_tmp_0 =5'h0;
          5 'b01110:
             casez_tmp_0 ={2'h1,io_in[9:7]};
          5 'b01111:
             casez_tmp_0 =5'h0;
          5 'b10000:
             casez_tmp_0 =io_in[11:7];
          5 'b10001:
             casez_tmp_0 =io_in[11:7];
          5 'b10010:
             casez_tmp_0 =io_in[11:7];
          5 'b10011:
             casez_tmp_0 =io_in[11:7];
          5 'b10100:
             casez_tmp_0 =io_in[12] ? ((|(io_in[6:2])) ? io_in[11:7]:5'h1):(|(io_in[6:2])) ? io_in[11:7]:5'h0;
          5 'b10101:
             casez_tmp_0 =io_in[11:7];
          5 'b10110:
             casez_tmp_0 =io_in[11:7];
          5 'b10111:
             casez_tmp_0 =io_in[11:7];
          5 'b11000:
             casez_tmp_0 =io_in[11:7];
          5 'b11001:
             casez_tmp_0 =io_in[11:7];
          5 'b11010:
             casez_tmp_0 =io_in[11:7];
          5 'b11011:
             casez_tmp_0 =io_in[11:7];
          5 'b11100:
             casez_tmp_0 =io_in[11:7];
          5 'b11101:
             casez_tmp_0 =io_in[11:7];
          5 'b11110:
             casez_tmp_0 =io_in[11:7];
          default :
             casez_tmp_0 =io_in[11:7];
         endcase 
       end
  
   reg [4:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_io_out_T_2)
          5 'b00000:
             casez_tmp_1 =5'h2;
          5 'b00001:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b00010:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b00011:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b00100:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b00101:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b00110:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b00111:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b01000:
             casez_tmp_1 =io_in[11:7];
          5 'b01001:
             casez_tmp_1 =io_in[11:7];
          5 'b01010:
             casez_tmp_1 =5'h0;
          5 'b01011:
             casez_tmp_1 =io_in[11:7];
          5 'b01100:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b01101:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b01110:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b01111:
             casez_tmp_1 ={2'h1,io_in[9:7]};
          5 'b10000:
             casez_tmp_1 =io_in[11:7];
          5 'b10001:
             casez_tmp_1 =5'h2;
          5 'b10010:
             casez_tmp_1 =5'h2;
          5 'b10011:
             casez_tmp_1 =5'h2;
          5 'b10100:
             casez_tmp_1 =io_in[12]|~(|(io_in[6:2])) ? io_in[11:7]:5'h0;
          5 'b10101:
             casez_tmp_1 =5'h2;
          5 'b10110:
             casez_tmp_1 =5'h2;
          5 'b10111:
             casez_tmp_1 =5'h2;
          5 'b11000:
             casez_tmp_1 =io_in[19:15];
          5 'b11001:
             casez_tmp_1 =io_in[19:15];
          5 'b11010:
             casez_tmp_1 =io_in[19:15];
          5 'b11011:
             casez_tmp_1 =io_in[19:15];
          5 'b11100:
             casez_tmp_1 =io_in[19:15];
          5 'b11101:
             casez_tmp_1 =io_in[19:15];
          5 'b11110:
             casez_tmp_1 =io_in[19:15];
          default :
             casez_tmp_1 =io_in[19:15];
         endcase 
       end
  
  assign io_out_bits=(&_io_out_T_2)|_io_out_T_61|_io_out_T_59|_io_out_T_57|_io_out_T_55|_io_out_T_53|_io_out_T_51|_io_out_T_49 ? io_in:_io_out_T_47 ? {3'h0,io_in[9:7],io_in[12],io_in[6:2],8'h13,io_in[11:10],10'h23}:_io_out_T_45 ? {4'h0,io_in[8:7],io_in[12],io_in[6:2],8'h12,io_in[11:9],9'h23}:_io_out_T_43 ? {3'h0,io_in[9:7],io_in[12],io_in[6:2],8'h13,io_in[11:10],10'h27}:_io_out_T_42_bits; 
  assign io_out_rd=casez_tmp_0; 
  assign io_out_rs1=casez_tmp_1; 
  assign io_out_rs2=(&_io_out_T_2)|_io_out_T_61|_io_out_T_59|_io_out_T_57|_io_out_T_55|_io_out_T_53|_io_out_T_51|_io_out_T_49 ? io_in[24:20]:_io_out_T_47|_io_out_T_45|_io_out_T_43|_io_out_T_41|_io_out_T_39|_io_out_T_37|_io_out_T_35|_io_out_T_33 ? io_in[6:2]:_io_out_T_31|_io_out_T_29 ? 5'h0:{2'h1,io_in[4:2]}; 
  assign io_rvc=io_in[1:0]!=2'h3; 
endmodule
 
module IBuf (
  input clock,
  input reset,
  output io_imem_ready,
  input io_imem_valid,
  input [33:0] io_imem_bits_pc,
  input [31:0] io_imem_bits_data,
  input io_imem_bits_xcpt_pf_inst,
  input io_imem_bits_xcpt_gf_inst,
  input io_imem_bits_xcpt_ae_inst,
  input io_imem_bits_replay,
  input io_kill,
  output [33:0] io_pc,
  input io_inst_0_ready,
  output io_inst_0_valid,
  output io_inst_0_bits_xcpt0_pf_inst,
  output io_inst_0_bits_xcpt0_gf_inst,
  output io_inst_0_bits_xcpt0_ae_inst,
  output io_inst_0_bits_xcpt1_pf_inst,
  output io_inst_0_bits_xcpt1_gf_inst,
  output io_inst_0_bits_xcpt1_ae_inst,
  output io_inst_0_bits_replay,
  output io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0] io_inst_0_bits_inst_rd,
  output [4:0] io_inst_0_bits_inst_rs1,
  output [4:0] io_inst_0_bits_inst_rs2,
  output [31:0] io_inst_0_bits_raw) ; 
   wire [1:0] nReady ;  
   wire _exp_io_rvc ;  
   reg nBufValid ;  
   reg [33:0] buf_pc ;  
   reg [31:0] buf_data ;  
   reg buf_xcpt_pf_inst ;  
   reg buf_xcpt_gf_inst ;  
   reg buf_xcpt_ae_inst ;  
   reg buf_replay ;  
   wire [1:0] _GEN={1'h0,io_imem_bits_pc[1]} ;  
   wire [1:0] _nIC_T_2=2'h2-_GEN ;  
   wire [1:0] _GEN_0={1'h0,nBufValid} ;  
   wire [1:0] _nICReady_T=nReady-_GEN_0 ;  
   wire _nBufValid_T=nReady>=_GEN_0 ;  
   wire [1:0] _nBufValid_T_6=_nIC_T_2-_nICReady_T ;  
   wire [190:0] _icData_T_4={63'h0,{2{{2{io_imem_bits_data[31:16]}}}},io_imem_bits_data,{2{io_imem_bits_data[15:0]}}}<<{185'h0,_GEN_0-2'h2-_GEN,4'h0} ;  
   wire [62:0] _icMask_T_2=63'hFFFFFFFF<<{58'h0,nBufValid,4'h0} ;  
   wire [31:0] inst=_icData_T_4[95:64]&_icMask_T_2[31:0]|buf_data&~(_icMask_T_2[31:0]) ;  
   wire [3:0] _valid_T=4'h1<<(io_imem_valid ? _nIC_T_2:2'h0)+_GEN_0 ;  
   wire [1:0] _valid_T_1=_valid_T[1:0]-2'h1 ;  
   wire [1:0] _bufMask_T_1=(2'h1<<_GEN_0)-2'h1 ;  
   wire [1:0] buf_replay_0=buf_replay ? _bufMask_T_1:2'h0 ;  
   wire [1:0] ic_replay=buf_replay_0|(io_imem_bits_replay ? _valid_T_1&~_bufMask_T_1:2'h0) ;  
   wire full_insn=_exp_io_rvc|_valid_T_1[1]|buf_replay_0[0] ;  
   wire [2:0] _io_inst_0_bits_xcpt1_T_5=_exp_io_rvc ? 3'h0:{_bufMask_T_1[1] ? buf_xcpt_pf_inst:io_imem_bits_xcpt_pf_inst,_bufMask_T_1[1] ? buf_xcpt_gf_inst:io_imem_bits_xcpt_gf_inst,_bufMask_T_1[1] ? buf_xcpt_ae_inst:io_imem_bits_xcpt_ae_inst} ;  
  assign nReady=full_insn ? (_exp_io_rvc ? 2'h1:2'h2):2'h0; 
   wire [63:0] _buf_data_T_1={{2{io_imem_bits_data[31:16]}},io_imem_bits_data}>>{58'h0,_GEN+_nICReady_T,4'h0} ;  
   wire _GEN_1=io_imem_valid&_nBufValid_T&_nICReady_T<_nIC_T_2&~(_nBufValid_T_6[1]) ;  
  always @( posedge clock)
       begin 
         if (reset)
            nBufValid <=1'h0;
          else 
            nBufValid <=~io_kill&(io_inst_0_ready ? (_GEN_1 ? _nBufValid_T_6[0]:~(_nBufValid_T|~nBufValid)&nBufValid-nReady[0]):nBufValid);
         if (io_inst_0_ready&_GEN_1)
            begin 
              buf_pc <=io_imem_bits_pc&34'h3FFFFFFFC|io_imem_bits_pc+{31'h0,_nICReady_T,1'h0}&34'h3;
              buf_data <={16'h0,_buf_data_T_1[15:0]};
              buf_xcpt_pf_inst <=io_imem_bits_xcpt_pf_inst;
              buf_xcpt_gf_inst <=io_imem_bits_xcpt_gf_inst;
              buf_xcpt_ae_inst <=io_imem_bits_xcpt_ae_inst;
              buf_replay <=io_imem_bits_replay;
            end 
       end
  
  RVCExpander exp(.io_in(inst),.io_out_bits(io_inst_0_bits_inst_bits),.io_out_rd(io_inst_0_bits_inst_rd),.io_out_rs1(io_inst_0_bits_inst_rs1),.io_out_rs2(io_inst_0_bits_inst_rs2),.io_rvc(_exp_io_rvc)); 
  assign io_imem_ready=io_inst_0_ready&_nBufValid_T&(_nICReady_T>=_nIC_T_2|~(_nBufValid_T_6[1])); 
  assign io_pc=nBufValid ? buf_pc:io_imem_bits_pc; 
  assign io_inst_0_valid=_valid_T_1[0]&full_insn; 
  assign io_inst_0_bits_xcpt0_pf_inst=_bufMask_T_1[0] ? buf_xcpt_pf_inst:io_imem_bits_xcpt_pf_inst; 
  assign io_inst_0_bits_xcpt0_gf_inst=_bufMask_T_1[0] ? buf_xcpt_gf_inst:io_imem_bits_xcpt_gf_inst; 
  assign io_inst_0_bits_xcpt0_ae_inst=_bufMask_T_1[0] ? buf_xcpt_ae_inst:io_imem_bits_xcpt_ae_inst; 
  assign io_inst_0_bits_xcpt1_pf_inst=_io_inst_0_bits_xcpt1_T_5[2]; 
  assign io_inst_0_bits_xcpt1_gf_inst=_io_inst_0_bits_xcpt1_T_5[1]; 
  assign io_inst_0_bits_xcpt1_ae_inst=_io_inst_0_bits_xcpt1_T_5[0]; 
  assign io_inst_0_bits_replay=ic_replay[0]|~_exp_io_rvc&ic_replay[1]; 
  assign io_inst_0_bits_rvc=_exp_io_rvc; 
  assign io_inst_0_bits_raw=inst; 
endmodule
 
module CSRFile (
  input clock,
  input reset,
  input io_ungated_clock,
  input io_interrupts_debug,
  input io_interrupts_mtip,
  input io_interrupts_msip,
  input io_interrupts_meip,
  input io_hartid,
  input [11:0] io_rw_addr,
  input [2:0] io_rw_cmd,
  output [63:0] io_rw_rdata,
  input [63:0] io_rw_wdata,
  input [31:0] io_decode_0_inst,
  output io_decode_0_read_illegal,
  output io_decode_0_write_illegal,
  output io_decode_0_write_flush,
  output io_decode_0_system_illegal,
  output io_decode_0_virtual_access_illegal,
  output io_decode_0_virtual_system_illegal,
  output io_csr_stall,
  output io_eret,
  output io_singleStep,
  output io_status_debug,
  output io_status_wfi,
  output [31:0] io_status_isa,
  output io_status_dv,
  output io_status_v,
  output [33:0] io_evec,
  input io_exception,
  input io_retire,
  input [63:0] io_cause,
  input [33:0] io_pc,
  input [33:0] io_tval,
  input io_gva,
  output [63:0] io_time,
  output io_interrupt,
  output [63:0] io_interrupt_cause,
  output io_bp_0_control_action,
  output [1:0] io_bp_0_control_tmatch,
  output io_bp_0_control_x,
  output io_bp_0_control_w,
  output io_bp_0_control_r,
  output [32:0] io_bp_0_address,
  output io_pmp_cfg_l_0,
  output io_pmp_cfg_l_1,
  output io_pmp_cfg_l_2,
  output io_pmp_cfg_l_3,
  output io_pmp_cfg_l_4,
  output io_pmp_cfg_l_5,
  output io_pmp_cfg_l_6,
  output io_pmp_cfg_l_7,
  output [1:0] io_pmp_cfg_a_0,
  output [1:0] io_pmp_cfg_a_1,
  output [1:0] io_pmp_cfg_a_2,
  output [1:0] io_pmp_cfg_a_3,
  output [1:0] io_pmp_cfg_a_4,
  output [1:0] io_pmp_cfg_a_5,
  output [1:0] io_pmp_cfg_a_6,
  output [1:0] io_pmp_cfg_a_7,
  output io_pmp_cfg_x_0,
  output io_pmp_cfg_x_1,
  output io_pmp_cfg_x_2,
  output io_pmp_cfg_x_3,
  output io_pmp_cfg_x_4,
  output io_pmp_cfg_x_5,
  output io_pmp_cfg_x_6,
  output io_pmp_cfg_x_7,
  output io_pmp_cfg_w_0,
  output io_pmp_cfg_w_1,
  output io_pmp_cfg_w_2,
  output io_pmp_cfg_w_3,
  output io_pmp_cfg_w_4,
  output io_pmp_cfg_w_5,
  output io_pmp_cfg_w_6,
  output io_pmp_cfg_w_7,
  output io_pmp_cfg_r_0,
  output io_pmp_cfg_r_1,
  output io_pmp_cfg_r_2,
  output io_pmp_cfg_r_3,
  output io_pmp_cfg_r_4,
  output io_pmp_cfg_r_5,
  output io_pmp_cfg_r_6,
  output io_pmp_cfg_r_7,
  output [29:0] io_pmp_addr_0,
  output [29:0] io_pmp_addr_1,
  output [29:0] io_pmp_addr_2,
  output [29:0] io_pmp_addr_3,
  output [29:0] io_pmp_addr_4,
  output [29:0] io_pmp_addr_5,
  output [29:0] io_pmp_addr_6,
  output [29:0] io_pmp_addr_7,
  output [31:0] io_pmp_mask_0,
  output [31:0] io_pmp_mask_1,
  output [31:0] io_pmp_mask_2,
  output [31:0] io_pmp_mask_3,
  output [31:0] io_pmp_mask_4,
  output [31:0] io_pmp_mask_5,
  output [31:0] io_pmp_mask_6,
  output [31:0] io_pmp_mask_7,
  output io_inhibit_cycle,
  input [31:0] io_inst_0,
  output io_trace_valid_0,
  output [33:0] io_trace_iaddr_0,
  output [31:0] io_trace_insn_0,
  output io_trace_exception_0,
  output [63:0] io_customCSRs_0_value) ; 
   wire [63:0] _io_rw_rdata_T_262 ;  
   reg io_status_cease_r ;  
   wire io_singleStep_0 ;  
   reg reg_mstatus_v ;  
   reg reg_mstatus_mpv ;  
   reg reg_mstatus_gva ;  
   reg [1:0] reg_mstatus_mpp ;  
   reg reg_mstatus_mpie ;  
   reg reg_mstatus_mie ;  
   reg reg_dcsr_ebreakm ;  
   reg [2:0] reg_dcsr_cause ;  
   reg reg_dcsr_v ;  
   reg reg_dcsr_step ;  
   reg reg_debug ;  
   reg [33:0] reg_dpc ;  
   reg [63:0] reg_dscratch0 ;  
   reg reg_singleStepped ;  
   reg reg_bp_0_control_dmode ;  
   reg reg_bp_0_control_action ;  
   reg [1:0] reg_bp_0_control_tmatch ;  
   reg reg_bp_0_control_x ;  
   reg reg_bp_0_control_w ;  
   reg reg_bp_0_control_r ;  
   reg [32:0] reg_bp_0_address ;  
   reg reg_pmp_cfg_l_0 ;  
   reg reg_pmp_cfg_l_1 ;  
   reg reg_pmp_cfg_l_2 ;  
   reg reg_pmp_cfg_l_3 ;  
   reg reg_pmp_cfg_l_4 ;  
   reg reg_pmp_cfg_l_5 ;  
   reg reg_pmp_cfg_l_6 ;  
   reg reg_pmp_cfg_l_7 ;  
   reg [1:0] reg_pmp_cfg_a_0 ;  
   reg [1:0] reg_pmp_cfg_a_1 ;  
   reg [1:0] reg_pmp_cfg_a_2 ;  
   reg [1:0] reg_pmp_cfg_a_3 ;  
   reg [1:0] reg_pmp_cfg_a_4 ;  
   reg [1:0] reg_pmp_cfg_a_5 ;  
   reg [1:0] reg_pmp_cfg_a_6 ;  
   reg [1:0] reg_pmp_cfg_a_7 ;  
   reg reg_pmp_cfg_x_0 ;  
   reg reg_pmp_cfg_x_1 ;  
   reg reg_pmp_cfg_x_2 ;  
   reg reg_pmp_cfg_x_3 ;  
   reg reg_pmp_cfg_x_4 ;  
   reg reg_pmp_cfg_x_5 ;  
   reg reg_pmp_cfg_x_6 ;  
   reg reg_pmp_cfg_x_7 ;  
   reg reg_pmp_cfg_w_0 ;  
   reg reg_pmp_cfg_w_1 ;  
   reg reg_pmp_cfg_w_2 ;  
   reg reg_pmp_cfg_w_3 ;  
   reg reg_pmp_cfg_w_4 ;  
   reg reg_pmp_cfg_w_5 ;  
   reg reg_pmp_cfg_w_6 ;  
   reg reg_pmp_cfg_w_7 ;  
   reg reg_pmp_cfg_r_0 ;  
   reg reg_pmp_cfg_r_1 ;  
   reg reg_pmp_cfg_r_2 ;  
   reg reg_pmp_cfg_r_3 ;  
   reg reg_pmp_cfg_r_4 ;  
   reg reg_pmp_cfg_r_5 ;  
   reg reg_pmp_cfg_r_6 ;  
   reg reg_pmp_cfg_r_7 ;  
   reg [29:0] reg_pmp_addr_0 ;  
   reg [29:0] reg_pmp_addr_1 ;  
   reg [29:0] reg_pmp_addr_2 ;  
   reg [29:0] reg_pmp_addr_3 ;  
   reg [29:0] reg_pmp_addr_4 ;  
   reg [29:0] reg_pmp_addr_5 ;  
   reg [29:0] reg_pmp_addr_6 ;  
   reg [29:0] reg_pmp_addr_7 ;  
   reg [63:0] reg_mie ;  
   reg [33:0] reg_mepc ;  
   reg [63:0] reg_mcause ;  
   reg [33:0] reg_mtval ;  
   reg [63:0] reg_mscratch ;  
   reg [31:0] reg_mtvec ;  
   reg reg_wfi ;  
   reg [2:0] reg_mcountinhibit ;  
   reg [5:0] small_0 ;  
   reg [57:0] large_0 ;  
   wire [63:0] value={large_0,small_0} ;  
   reg [5:0] small_1 ;  
   reg [57:0] large_1 ;  
   wire [63:0] io_time_0={large_1,small_1} ;  
   wire [15:0] read_mip={4'h0,io_interrupts_meip,3'h0,io_interrupts_mtip,3'h0,io_interrupts_msip,3'h0} ;  
   wire [15:0] _GEN=reg_mie[15:0]&read_mip ;  
   wire [15:0] m_interrupts=reg_mstatus_mie ? _GEN:16'h0 ;  
   wire [29:0] _GEN_0={reg_pmp_addr_0[28:0],reg_pmp_cfg_a_0[0]} ;  
   wire [29:0] _GEN_1={reg_pmp_addr_1[28:0],reg_pmp_cfg_a_1[0]} ;  
   wire [29:0] _GEN_2={reg_pmp_addr_2[28:0],reg_pmp_cfg_a_2[0]} ;  
   wire [29:0] _GEN_3={reg_pmp_addr_3[28:0],reg_pmp_cfg_a_3[0]} ;  
   wire [29:0] _GEN_4={reg_pmp_addr_4[28:0],reg_pmp_cfg_a_4[0]} ;  
   wire [29:0] _GEN_5={reg_pmp_addr_5[28:0],reg_pmp_cfg_a_5[0]} ;  
   wire [29:0] _GEN_6={reg_pmp_addr_6[28:0],reg_pmp_cfg_a_6[0]} ;  
   wire [29:0] _GEN_7={reg_pmp_addr_7[28:0],reg_pmp_cfg_a_7[0]} ;  
   reg [63:0] reg_misa ;  
   wire [31:0] _read_mtvec_T_5=reg_mtvec&{24'hFFFFFF,~(reg_mtvec[0] ? 8'hFE:8'h2)} ;  
   wire [33:0] _io_evec_T_20=~reg_mepc ;  
   wire [1:0] _GEN_8={~(reg_misa[2]),1'h1} ;  
   wire [33:0] _GEN_9=~{_io_evec_T_20[33:2],_io_evec_T_20[1:0]|_GEN_8} ;  
   wire [33:0] _io_evec_T_10=~reg_dpc ;  
   wire [33:0] _GEN_10=~{_io_evec_T_10[33:2],_io_evec_T_10[1:0]|_GEN_8} ;  
   reg [63:0] reg_custom_0 ;  
   wire [11:0] decoded_decoded_invInputs=~io_rw_addr ;  
   wire [11:0] _decoded_decoded_T={decoded_decoded_invInputs[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_2={io_rw_addr[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_4={decoded_decoded_invInputs[0],decoded_decoded_invInputs[1],io_rw_addr[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_6={io_rw_addr[0],decoded_decoded_invInputs[1],io_rw_addr[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [10:0] _decoded_decoded_T_8={decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],io_rw_addr[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_68={decoded_decoded_invInputs[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],io_rw_addr[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_70={io_rw_addr[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],io_rw_addr[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_72={decoded_decoded_invInputs[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],io_rw_addr[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_74={io_rw_addr[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],io_rw_addr[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [10:0] _decoded_decoded_T_78={decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_82={decoded_decoded_invInputs[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_84={io_rw_addr[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_86={decoded_decoded_invInputs[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_88={io_rw_addr[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_90={decoded_decoded_invInputs[0],decoded_decoded_invInputs[1],io_rw_addr[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_92={io_rw_addr[0],decoded_decoded_invInputs[1],io_rw_addr[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_94={decoded_decoded_invInputs[0],io_rw_addr[1],io_rw_addr[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_96={io_rw_addr[0],io_rw_addr[1],io_rw_addr[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_116={io_rw_addr[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_118={decoded_decoded_invInputs[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_122={decoded_decoded_invInputs[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],decoded_decoded_invInputs[11]} ;  
   wire [11:0] _decoded_decoded_T_124={io_rw_addr[0],decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],decoded_decoded_invInputs[11]} ;  
   wire [10:0] _decoded_decoded_T_126={io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],io_rw_addr[5],decoded_decoded_invInputs[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],decoded_decoded_invInputs[11]} ;  
   wire [5:0] _decoded_decoded_T_128={io_rw_addr[6],io_rw_addr[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],decoded_decoded_invInputs[11]} ;  
   wire [10:0] _decoded_decoded_T_130={decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],io_rw_addr[11]} ;  
   wire [11:0] _decoded_decoded_T_132={decoded_decoded_invInputs[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],io_rw_addr[11]} ;  
   wire [63:0] _wdata_T_2=(io_rw_cmd[1] ? _io_rw_rdata_T_262:64'h0)|io_rw_wdata ;  
   wire [63:0] _wdata_T_6=~((&(io_rw_cmd[1:0])) ? io_rw_wdata:64'h0) ;  
   wire system_insn=io_rw_cmd==3'h4 ;  
   wire [11:0] _GEN_11=~io_rw_addr ;  
   wire insn_call=system_insn&(&{_GEN_11[0],_GEN_11[1],_GEN_11[2],_GEN_11[3],_GEN_11[4],_GEN_11[5],_GEN_11[6],_GEN_11[7],_GEN_11[8],_GEN_11[9],_GEN_11[10],_GEN_11[11]}) ;  
   wire insn_break=system_insn&(&{io_rw_addr[0],_GEN_11[1],_GEN_11[2],_GEN_11[3],_GEN_11[4],_GEN_11[5],_GEN_11[6],_GEN_11[7],_GEN_11[8],_GEN_11[9],_GEN_11[10],_GEN_11[11]}) ;  
   wire insn_ret=system_insn&(|{&{_GEN_11[2],_GEN_11[3],_GEN_11[4],_GEN_11[5],_GEN_11[6],_GEN_11[7],io_rw_addr[8],io_rw_addr[9],_GEN_11[10],_GEN_11[11]},&{io_rw_addr[10],_GEN_11[11]}}) ;  
   wire [9:0] decoded_invInputs_1=~(io_decode_0_inst[31:22]) ;  
   wire [31:0] _GEN_12={27'h0,io_decode_0_inst[24:20]} ;  
   wire [31:0] _io_decode_0_virtual_access_illegal_T_3=32'h0>>_GEN_12 ;  
   wire [31:0] _io_decode_0_virtual_access_illegal_T_6=32'h0>>_GEN_12 ;  
   wire csr_exists=io_decode_0_inst[31:20]==12'h7A0|io_decode_0_inst[31:20]==12'h7A1|io_decode_0_inst[31:20]==12'h7A2|io_decode_0_inst[31:20]==12'h7A3|io_decode_0_inst[31:20]==12'h301|io_decode_0_inst[31:20]==12'h300|io_decode_0_inst[31:20]==12'h305|io_decode_0_inst[31:20]==12'h344|io_decode_0_inst[31:20]==12'h304|io_decode_0_inst[31:20]==12'h340|io_decode_0_inst[31:20]==12'h341|io_decode_0_inst[31:20]==12'h343|io_decode_0_inst[31:20]==12'h342|io_decode_0_inst[31:20]==12'hF14|io_decode_0_inst[31:20]==12'h7B0|io_decode_0_inst[31:20]==12'h7B1|io_decode_0_inst[31:20]==12'h7B2|io_decode_0_inst[31:20]==12'h320|io_decode_0_inst[31:20]==12'hB00|io_decode_0_inst[31:20]==12'hB02|io_decode_0_inst[31:20]==12'h323|io_decode_0_inst[31:20]==12'hB03|io_decode_0_inst[31:20]==12'hC03|io_decode_0_inst[31:20]==12'h324|io_decode_0_inst[31:20]==12'hB04|io_decode_0_inst[31:20]==12'hC04|io_decode_0_inst[31:20]==12'h325|io_decode_0_inst[31:20]==12'hB05|io_decode_0_inst[31:20]==12'hC05|io_decode_0_inst[31:20]==12'h326|io_decode_0_inst[31:20]==12'hB06|io_decode_0_inst[31:20]==12'hC06|io_decode_0_inst[31:20]==12'h327|io_decode_0_inst[31:20]==12'hB07|io_decode_0_inst[31:20]==12'hC07|io_decode_0_inst[31:20]==12'h328|io_decode_0_inst[31:20]==12'hB08|io_decode_0_inst[31:20]==12'hC08|io_decode_0_inst[31:20]==12'h329|io_decode_0_inst[31:20]==12'hB09|io_decode_0_inst[31:20]==12'hC09|io_decode_0_inst[31:20]==12'h32A|io_decode_0_inst[31:20]==12'hB0A|io_decode_0_inst[31:20]==12'hC0A|io_decode_0_inst[31:20]==12'h32B|io_decode_0_inst[31:20]==12'hB0B|io_decode_0_inst[31:20]==12'hC0B|io_decode_0_inst[31:20]==12'h32C|io_decode_0_inst[31:20]==12'hB0C|io_decode_0_inst[31:20]==12'hC0C|io_decode_0_inst[31:20]==12'h32D|io_decode_0_inst[31:20]==12'hB0D|io_decode_0_inst[31:20]==12'hC0D|io_decode_0_inst[31:20]==12'h32E|io_decode_0_inst[31:20]==12'hB0E|io_decode_0_inst[31:20]==12'hC0E|io_decode_0_inst[31:20]==12'h32F|io_decode_0_inst[31:20]==12'hB0F|io_decode_0_inst[31:20]==12'hC0F|io_decode_0_inst[31:20]==12'h330|io_decode_0_inst[31:20]==12'hB10|io_decode_0_inst[31:20]==12'hC10|io_decode_0_inst[31:20]==12'h331|io_decode_0_inst[31:20]==12'hB11|io_decode_0_inst[31:20]==12'hC11|io_decode_0_inst[31:20]==12'h332|io_decode_0_inst[31:20]==12'hB12|io_decode_0_inst[31:20]==12'hC12|io_decode_0_inst[31:20]==12'h333|io_decode_0_inst[31:20]==12'hB13|io_decode_0_inst[31:20]==12'hC13|io_decode_0_inst[31:20]==12'h334|io_decode_0_inst[31:20]==12'hB14|io_decode_0_inst[31:20]==12'hC14|io_decode_0_inst[31:20]==12'h335|io_decode_0_inst[31:20]==12'hB15|io_decode_0_inst[31:20]==12'hC15|io_decode_0_inst[31:20]==12'h336|io_decode_0_inst[31:20]==12'hB16|io_decode_0_inst[31:20]==12'hC16|io_decode_0_inst[31:20]==12'h337|io_decode_0_inst[31:20]==12'hB17|io_decode_0_inst[31:20]==12'hC17|io_decode_0_inst[31:20]==12'h338|io_decode_0_inst[31:20]==12'hB18|io_decode_0_inst[31:20]==12'hC18|io_decode_0_inst[31:20]==12'h339|io_decode_0_inst[31:20]==12'hB19|io_decode_0_inst[31:20]==12'hC19|io_decode_0_inst[31:20]==12'h33A|io_decode_0_inst[31:20]==12'hB1A|io_decode_0_inst[31:20]==12'hC1A|io_decode_0_inst[31:20]==12'h33B|io_decode_0_inst[31:20]==12'hB1B|io_decode_0_inst[31:20]==12'hC1B|io_decode_0_inst[31:20]==12'h33C|io_decode_0_inst[31:20]==12'hB1C|io_decode_0_inst[31:20]==12'hC1C|io_decode_0_inst[31:20]==12'h33D|io_decode_0_inst[31:20]==12'hB1D|io_decode_0_inst[31:20]==12'hC1D|io_decode_0_inst[31:20]==12'h33E|io_decode_0_inst[31:20]==12'hB1E|io_decode_0_inst[31:20]==12'hC1E|io_decode_0_inst[31:20]==12'h33F|io_decode_0_inst[31:20]==12'hB1F|io_decode_0_inst[31:20]==12'hC1F|io_decode_0_inst[31:20]==12'hC00|io_decode_0_inst[31:20]==12'hC02|io_decode_0_inst[31:20]==12'h3A0|io_decode_0_inst[31:20]==12'h3A2|io_decode_0_inst[31:20]==12'h3B0|io_decode_0_inst[31:20]==12'h3B1|io_decode_0_inst[31:20]==12'h3B2|io_decode_0_inst[31:20]==12'h3B3|io_decode_0_inst[31:20]==12'h3B4|io_decode_0_inst[31:20]==12'h3B5|io_decode_0_inst[31:20]==12'h3B6|io_decode_0_inst[31:20]==12'h3B7|io_decode_0_inst[31:20]==12'h3B8|io_decode_0_inst[31:20]==12'h3B9|io_decode_0_inst[31:20]==12'h3BA|io_decode_0_inst[31:20]==12'h3BB|io_decode_0_inst[31:20]==12'h3BC|io_decode_0_inst[31:20]==12'h3BD|io_decode_0_inst[31:20]==12'h3BE|io_decode_0_inst[31:20]==12'h3BF|io_decode_0_inst[31:20]==12'h7C1|io_decode_0_inst[31:20]==12'hF12|io_decode_0_inst[31:20]==12'hF11|io_decode_0_inst[31:20]==12'hF13|io_decode_0_inst[31:20]==12'hF15 ;  
   wire [5:0] io_decode_0_read_illegal_invInputs=~(io_decode_0_inst[31:26]) ;  
   wire [11:0] io_decode_0_write_flush_addr_m={io_decode_0_inst[31:30],io_decode_0_inst[29:20]|10'h300} ;  
   wire [63:0] cause=insn_call ? {60'h0,{3'h1,~reg_mstatus_v}-4'h8}:insn_break ? 64'h3:io_cause ;  
   wire _causeIsDebugTrigger_T_2=cause[7:0]==8'hE ;  
   wire causeIsDebugInt=cause[63]&_causeIsDebugTrigger_T_2 ;  
   wire causeIsDebugTrigger=~(cause[63])&_causeIsDebugTrigger_T_2 ;  
   wire trapToDebug=reg_singleStepped|causeIsDebugInt|causeIsDebugTrigger|~(cause[63])&insn_break&reg_dcsr_ebreakm|reg_debug ;  
   wire _exception_T=insn_call|insn_break ;  
  assign io_singleStep_0=reg_dcsr_step&~reg_debug; 
   wire exception=_exception_T|io_exception ;  
   wire [2:0] _GEN_13={1'h0,{1'h0,insn_ret}+{1'h0,insn_call}}+{1'h0,{1'h0,insn_break}+{1'h0,io_exception}} ;  
  always @( posedge clock)
       begin 
         if (~reset&(|(_GEN_13[2:1])))
            begin 
              if (1)$display("Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:1010 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1.U, \"these conditions must be mutually exclusive\")\n");
              if (1)$display("");
            end 
         if (~reset&~(~reg_singleStepped|~io_retire))
            begin 
              if (1)$display("Assertion failed\n    at CSR.scala:1019 assert(!reg_singleStepped || io.retire === 0.U)\n");
              if (1)$display("");
            end 
       end
  
   wire _GEN_14=io_rw_addr[10]&io_rw_addr[7] ;  
   wire io_csr_stall_0=reg_wfi|io_status_cease_r ;  
   wire [63:0] _io_rw_rdata_T_137=((&_decoded_decoded_T_116) ? {4'h2,reg_bp_0_control_dmode,46'h40000000000,reg_bp_0_control_action,3'h0,reg_bp_0_control_tmatch,4'h8,reg_bp_0_control_x,reg_bp_0_control_w,reg_bp_0_control_r}:64'h0)|((&_decoded_decoded_T_118) ? {{31{reg_bp_0_address[32]}},reg_bp_0_address}:64'h0)|((&_decoded_decoded_T_2) ? reg_misa:64'h0)|((&_decoded_decoded_T) ? {24'h0,reg_mstatus_mpv,reg_mstatus_gva,25'h0,reg_mstatus_mpp,3'h0,reg_mstatus_mpie,3'h0,reg_mstatus_mie,3'h0}:64'h0)|((&_decoded_decoded_T_6) ? {32'h0,_read_mtvec_T_5}:64'h0) ;  
   wire [63:0] _io_rw_rdata_T_143={_io_rw_rdata_T_137[63:16],_io_rw_rdata_T_137[15:0]|((&{io_rw_addr[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],io_rw_addr[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],decoded_decoded_invInputs[10],decoded_decoded_invInputs[11]}) ? read_mip:16'h0)}|((&_decoded_decoded_T_4) ? reg_mie:64'h0)|((&_decoded_decoded_T_68) ? reg_mscratch:64'h0)|((&_decoded_decoded_T_70) ? {{30{_GEN_9[33]}},_GEN_9}:64'h0)|((&_decoded_decoded_T_74) ? {{30{reg_mtval[33]}},reg_mtval}:64'h0)|((&_decoded_decoded_T_72) ? reg_mcause:64'h0) ;  
   wire [63:0] _io_rw_rdata_T_147={_io_rw_rdata_T_143[63:32],{_io_rw_rdata_T_143[31:1],_io_rw_rdata_T_143[0]|(&{decoded_decoded_invInputs[0],decoded_decoded_invInputs[1],io_rw_addr[2],decoded_decoded_invInputs[3],io_rw_addr[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],io_rw_addr[11]})&io_hartid}|((&_decoded_decoded_T_122) ? {16'h4000,reg_dcsr_ebreakm,6'h0,reg_dcsr_cause,reg_dcsr_v,2'h0,reg_dcsr_step,2'h3}:32'h0)}|((&_decoded_decoded_T_124) ? {{30{_GEN_10[33]}},_GEN_10}:64'h0)|((&_decoded_decoded_T_126) ? reg_dscratch0:64'h0) ;  
   wire [63:0] _io_rw_rdata_T_241={_io_rw_rdata_T_147[63:3],_io_rw_rdata_T_147[2:0]|((&_decoded_decoded_T_8) ? reg_mcountinhibit:3'h0)}|((&_decoded_decoded_T_130) ? io_time_0:64'h0)|((&_decoded_decoded_T_132) ? value:64'h0)|((&{decoded_decoded_invInputs[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],decoded_decoded_invInputs[8],decoded_decoded_invInputs[9],io_rw_addr[10],io_rw_addr[11]}) ? io_time_0:64'h0)|((&{decoded_decoded_invInputs[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],decoded_decoded_invInputs[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],decoded_decoded_invInputs[8],decoded_decoded_invInputs[9],io_rw_addr[10],io_rw_addr[11]}) ? value:64'h0)|((&_decoded_decoded_T_78) ? {reg_pmp_cfg_l_7,2'h0,reg_pmp_cfg_a_7,reg_pmp_cfg_x_7,reg_pmp_cfg_w_7,reg_pmp_cfg_r_7,reg_pmp_cfg_l_6,2'h0,reg_pmp_cfg_a_6,reg_pmp_cfg_x_6,reg_pmp_cfg_w_6,reg_pmp_cfg_r_6,reg_pmp_cfg_l_5,2'h0,reg_pmp_cfg_a_5,reg_pmp_cfg_x_5,reg_pmp_cfg_w_5,reg_pmp_cfg_r_5,reg_pmp_cfg_l_4,2'h0,reg_pmp_cfg_a_4,reg_pmp_cfg_x_4,reg_pmp_cfg_w_4,reg_pmp_cfg_r_4,reg_pmp_cfg_l_3,2'h0,reg_pmp_cfg_a_3,reg_pmp_cfg_x_3,reg_pmp_cfg_w_3,reg_pmp_cfg_r_3,reg_pmp_cfg_l_2,2'h0,reg_pmp_cfg_a_2,reg_pmp_cfg_x_2,reg_pmp_cfg_w_2,reg_pmp_cfg_r_2,reg_pmp_cfg_l_1,2'h0,reg_pmp_cfg_a_1,reg_pmp_cfg_x_1,reg_pmp_cfg_w_1,reg_pmp_cfg_r_1,reg_pmp_cfg_l_0,2'h0,reg_pmp_cfg_a_0,reg_pmp_cfg_x_0,reg_pmp_cfg_w_0,reg_pmp_cfg_r_0}:64'h0) ;  
   wire [29:0] _GEN_15=_io_rw_rdata_T_241[29:0]|((&_decoded_decoded_T_82) ? reg_pmp_addr_0:30'h0)|((&_decoded_decoded_T_84) ? reg_pmp_addr_1:30'h0)|((&_decoded_decoded_T_86) ? reg_pmp_addr_2:30'h0)|((&_decoded_decoded_T_88) ? reg_pmp_addr_3:30'h0)|((&_decoded_decoded_T_90) ? reg_pmp_addr_4:30'h0)|((&_decoded_decoded_T_92) ? reg_pmp_addr_5:30'h0)|((&_decoded_decoded_T_94) ? reg_pmp_addr_6:30'h0)|((&_decoded_decoded_T_96) ? reg_pmp_addr_7:30'h0) ;  
  assign _io_rw_rdata_T_262=((&_decoded_decoded_T_128) ? reg_custom_0:64'h0)|((&{io_rw_addr[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],io_rw_addr[11]}) ? 64'h20181004:64'h0)|{_io_rw_rdata_T_241[63:30],_GEN_15[29:1],_GEN_15[0]|(&{decoded_decoded_invInputs[0],io_rw_addr[1],decoded_decoded_invInputs[2],decoded_decoded_invInputs[3],io_rw_addr[4],decoded_decoded_invInputs[5],decoded_decoded_invInputs[6],decoded_decoded_invInputs[7],io_rw_addr[8],io_rw_addr[9],io_rw_addr[10],io_rw_addr[11]})}; 
   wire _csr_wen_T_4=io_rw_cmd==3'h6|(&io_rw_cmd)|io_rw_cmd==3'h5 ;  
   wire [5:0] _GEN_16=_wdata_T_2[5:0]&_wdata_T_6[5:0] ;  
   wire [47:0] _newBPC_T_8=((io_rw_cmd[1] ? {reg_bp_0_control_dmode,46'h40000000000,reg_bp_0_control_action}:48'h0)|io_rw_wdata[59:12])&~((&(io_rw_cmd[1:0])) ? io_rw_wdata[59:12]:48'h0) ;  
   wire dMode=_newBPC_T_8[47]&reg_debug ;  
   wire [6:0] nextSmall={1'h0,small_0}+{6'h0,io_retire} ;  
   wire _GEN_17=~insn_ret|_GEN_14 ;  
   wire [31:0] _new_dcsr_WIRE=_wdata_T_2[31:0]&_wdata_T_6[31:0] ;  
   wire [63:0] wdata=_wdata_T_2&_wdata_T_6 ;  
   wire [33:0] epc={io_pc[33:1],1'h0} ;  
   wire _GEN_18=exception&trapToDebug&~reg_debug ;  
   wire _GEN_19=~exception|trapToDebug ;  
   wire [33:0] _GEN_20={wdata[33:1],1'h0} ;  
   wire _GEN_21=~reg_bp_0_control_dmode|reg_debug ;  
   wire _GEN_22=_csr_wen_T_4&_GEN_21&(&_decoded_decoded_T_116) ;  
   wire [7:0] _newCfg_WIRE=_wdata_T_2[7:0]&_wdata_T_6[7:0] ;  
   wire _GEN_23=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_0 ;  
   wire [29:0] _GEN_24=_wdata_T_2[29:0]&_wdata_T_6[29:0] ;  
   wire [7:0] _newCfg_WIRE_1=_wdata_T_2[15:8]&_wdata_T_6[15:8] ;  
   wire _GEN_25=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_1 ;  
   wire [7:0] _newCfg_WIRE_2=_wdata_T_2[23:16]&_wdata_T_6[23:16] ;  
   wire _GEN_26=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_2 ;  
   wire [7:0] _newCfg_WIRE_3=_wdata_T_2[31:24]&_wdata_T_6[31:24] ;  
   wire _GEN_27=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_3 ;  
   wire [7:0] _newCfg_WIRE_4=_wdata_T_2[39:32]&_wdata_T_6[39:32] ;  
   wire _GEN_28=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_4 ;  
   wire [7:0] _newCfg_WIRE_5=_wdata_T_2[47:40]&_wdata_T_6[47:40] ;  
   wire _GEN_29=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_5 ;  
   wire [7:0] _newCfg_WIRE_6=_wdata_T_2[55:48]&_wdata_T_6[55:48] ;  
   wire _GEN_30=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_6 ;  
   wire _GEN_31=reg_pmp_cfg_l_7&~(reg_pmp_cfg_a_7[1])&reg_pmp_cfg_a_7[0] ;  
   wire [7:0] _newCfg_T_49=_wdata_T_2[63:56]&_wdata_T_6[63:56] ;  
   wire _GEN_32=_csr_wen_T_4&(&_decoded_decoded_T_78)&~reg_pmp_cfg_l_7 ;  
   wire [63:0] _reg_misa_T=~wdata ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              reg_mstatus_v <=1'h0;
              reg_mstatus_mpv <=1'h0;
              reg_mstatus_gva <=1'h0;
              reg_mstatus_mpp <=2'h3;
              reg_mstatus_mpie <=1'h0;
              reg_mstatus_mie <=1'h0;
              reg_dcsr_ebreakm <=1'h0;
              reg_dcsr_cause <=3'h0;
              reg_dcsr_v <=1'h0;
              reg_dcsr_step <=1'h0;
              reg_debug <=1'h0;
              reg_bp_0_control_dmode <=1'h0;
              reg_bp_0_control_action <=1'h0;
              reg_bp_0_control_x <=1'h0;
              reg_bp_0_control_w <=1'h0;
              reg_bp_0_control_r <=1'h0;
              reg_pmp_cfg_l_0 <=1'h0;
              reg_pmp_cfg_l_1 <=1'h0;
              reg_pmp_cfg_l_2 <=1'h0;
              reg_pmp_cfg_l_3 <=1'h0;
              reg_pmp_cfg_l_4 <=1'h0;
              reg_pmp_cfg_l_5 <=1'h0;
              reg_pmp_cfg_l_6 <=1'h0;
              reg_pmp_cfg_l_7 <=1'h0;
              reg_pmp_cfg_a_0 <=2'h0;
              reg_pmp_cfg_a_1 <=2'h0;
              reg_pmp_cfg_a_2 <=2'h0;
              reg_pmp_cfg_a_3 <=2'h0;
              reg_pmp_cfg_a_4 <=2'h0;
              reg_pmp_cfg_a_5 <=2'h0;
              reg_pmp_cfg_a_6 <=2'h0;
              reg_pmp_cfg_a_7 <=2'h0;
              reg_mcause <=64'h0;
              reg_mtvec <=32'h0;
              reg_mcountinhibit <=3'h0;
              small_0 <=6'h0;
              large_0 <=58'h0;
              reg_misa <=64'h8000000000801105;
              reg_custom_0 <=64'h208;
              io_status_cease_r <=1'h0;
            end 
          else 
            begin 
              reg_mstatus_v <=~insn_ret&(~exception|trapToDebug&reg_debug)&reg_mstatus_v;
              reg_mstatus_mpv <=_GEN_17&(_GEN_19 ? reg_mstatus_mpv:reg_mstatus_v);
              if (_GEN_19)
                 begin 
                 end 
               else 
                 reg_mstatus_gva <=io_gva;
              if (_GEN_17&_GEN_19)
                 begin 
                 end 
               else 
                 reg_mstatus_mpp <=2'h3;
              if (_csr_wen_T_4&(&_decoded_decoded_T))
                 begin 
                   reg_mstatus_mpie <=wdata[7];
                   reg_mstatus_mie <=wdata[3];
                 end 
               else 
                 begin 
                   reg_mstatus_mpie <=insn_ret&~_GEN_14|(_GEN_19 ? reg_mstatus_mpie:reg_mstatus_mie);
                   if (_GEN_17)
                      reg_mstatus_mie <=_GEN_19&reg_mstatus_mie;
                    else 
                      reg_mstatus_mie <=reg_mstatus_mpie;
                 end 
              if (_csr_wen_T_4&(&_decoded_decoded_T_122))
                 begin 
                   reg_dcsr_ebreakm <=_new_dcsr_WIRE[15];
                   reg_dcsr_step <=_new_dcsr_WIRE[2];
                 end 
              if (_GEN_18)
                 begin 
                   reg_dcsr_cause <=reg_singleStepped ? 3'h4:{1'h0,causeIsDebugInt ? 2'h3:causeIsDebugTrigger ? 2'h2:2'h1};
                   reg_dcsr_v <=reg_mstatus_v;
                 end 
              reg_debug <=~(insn_ret&_GEN_14)&(_GEN_18|reg_debug);
              if (_GEN_22)
                 begin 
                   reg_bp_0_control_dmode <=dMode;
                   reg_bp_0_control_action <=dMode&_newBPC_T_8[0];
                   reg_bp_0_control_x <=wdata[2];
                   reg_bp_0_control_w <=wdata[1];
                   reg_bp_0_control_r <=wdata[0];
                 end 
              if (_GEN_23)
                 begin 
                   reg_pmp_cfg_l_0 <=_newCfg_WIRE[7];
                   reg_pmp_cfg_a_0 <=_newCfg_WIRE[4:3];
                 end 
              if (_GEN_25)
                 begin 
                   reg_pmp_cfg_l_1 <=_newCfg_WIRE_1[7];
                   reg_pmp_cfg_a_1 <=_newCfg_WIRE_1[4:3];
                 end 
              if (_GEN_26)
                 begin 
                   reg_pmp_cfg_l_2 <=_newCfg_WIRE_2[7];
                   reg_pmp_cfg_a_2 <=_newCfg_WIRE_2[4:3];
                 end 
              if (_GEN_27)
                 begin 
                   reg_pmp_cfg_l_3 <=_newCfg_WIRE_3[7];
                   reg_pmp_cfg_a_3 <=_newCfg_WIRE_3[4:3];
                 end 
              if (_GEN_28)
                 begin 
                   reg_pmp_cfg_l_4 <=_newCfg_WIRE_4[7];
                   reg_pmp_cfg_a_4 <=_newCfg_WIRE_4[4:3];
                 end 
              if (_GEN_29)
                 begin 
                   reg_pmp_cfg_l_5 <=_newCfg_WIRE_5[7];
                   reg_pmp_cfg_a_5 <=_newCfg_WIRE_5[4:3];
                 end 
              if (_GEN_30)
                 begin 
                   reg_pmp_cfg_l_6 <=_newCfg_WIRE_6[7];
                   reg_pmp_cfg_a_6 <=_newCfg_WIRE_6[4:3];
                 end 
              if (_GEN_32)
                 begin 
                   reg_pmp_cfg_l_7 <=_newCfg_T_49[7];
                   reg_pmp_cfg_a_7 <=_newCfg_T_49[4:3];
                 end 
              if (_csr_wen_T_4&(&_decoded_decoded_T_72))
                 reg_mcause <=wdata&64'h800000000000000F;
               else 
                 if (_GEN_19)
                    begin 
                    end 
                  else 
                    reg_mcause <=cause;
              if (_csr_wen_T_4&(&_decoded_decoded_T_6))
                 reg_mtvec <=_new_dcsr_WIRE;
              if (_csr_wen_T_4&(&_decoded_decoded_T_8))
                 reg_mcountinhibit <=_wdata_T_2[2:0]&_wdata_T_6[2:0]&3'h5;
              if (_csr_wen_T_4&(&_decoded_decoded_T_132))
                 begin 
                   small_0 <=_GEN_16;
                   large_0 <=_wdata_T_2[63:6]&_wdata_T_6[63:6];
                 end 
               else 
                 begin 
                   if (reg_mcountinhibit[2])
                      begin 
                      end 
                    else 
                      small_0 <=nextSmall[5:0];
                   if (nextSmall[6]&~(reg_mcountinhibit[2]))
                      large_0 <=large_0+58'h1;
                 end 
              if (_csr_wen_T_4&(&_decoded_decoded_T_2)&(~(io_pc[1])|_wdata_T_2[2]&_wdata_T_6[2]))
                 reg_misa <=~{_reg_misa_T[63:4],_reg_misa_T[3:0]|{~(_wdata_T_2[5]&_wdata_T_6[5]),3'h0}}&64'h1005|reg_misa&64'hFFFFFFFFFFFFEFFA;
              if (_csr_wen_T_4&(&_decoded_decoded_T_128))
                 reg_custom_0 <=wdata&64'h208|reg_custom_0&64'hFFFFFFFFFFFFFDF7;
              io_status_cease_r <=system_insn&(&{io_rw_addr[2],_GEN_11[3],_GEN_11[4],_GEN_11[5],_GEN_11[6],_GEN_11[7],io_rw_addr[8],io_rw_addr[9],_GEN_11[10],_GEN_11[11]})|io_status_cease_r;
            end 
         if (_csr_wen_T_4&(&_decoded_decoded_T_124))
            reg_dpc <=_GEN_20;
          else 
            if (_GEN_18)
               reg_dpc <=epc;
         if (_csr_wen_T_4&(&_decoded_decoded_T_126))
            reg_dscratch0 <=wdata;
         reg_singleStepped <=io_singleStep_0&(io_retire|exception|reg_singleStepped);
         if (_GEN_22)
            reg_bp_0_control_tmatch <=wdata[8:7];
         if (_csr_wen_T_4&_GEN_21&(&_decoded_decoded_T_118))
            reg_bp_0_address <=_wdata_T_2[32:0]&_wdata_T_6[32:0];
         if (_GEN_23)
            begin 
              reg_pmp_cfg_x_0 <=_newCfg_WIRE[2];
              reg_pmp_cfg_w_0 <=_newCfg_WIRE[1]&_newCfg_WIRE[0];
              reg_pmp_cfg_r_0 <=_newCfg_WIRE[0];
            end 
         if (_GEN_25)
            begin 
              reg_pmp_cfg_x_1 <=_newCfg_WIRE_1[2];
              reg_pmp_cfg_w_1 <=_newCfg_WIRE_1[1]&_newCfg_WIRE_1[0];
              reg_pmp_cfg_r_1 <=_newCfg_WIRE_1[0];
            end 
         if (_GEN_26)
            begin 
              reg_pmp_cfg_x_2 <=_newCfg_WIRE_2[2];
              reg_pmp_cfg_w_2 <=_newCfg_WIRE_2[1]&_newCfg_WIRE_2[0];
              reg_pmp_cfg_r_2 <=_newCfg_WIRE_2[0];
            end 
         if (_GEN_27)
            begin 
              reg_pmp_cfg_x_3 <=_newCfg_WIRE_3[2];
              reg_pmp_cfg_w_3 <=_newCfg_WIRE_3[1]&_newCfg_WIRE_3[0];
              reg_pmp_cfg_r_3 <=_newCfg_WIRE_3[0];
            end 
         if (_GEN_28)
            begin 
              reg_pmp_cfg_x_4 <=_newCfg_WIRE_4[2];
              reg_pmp_cfg_w_4 <=_newCfg_WIRE_4[1]&_newCfg_WIRE_4[0];
              reg_pmp_cfg_r_4 <=_newCfg_WIRE_4[0];
            end 
         if (_GEN_29)
            begin 
              reg_pmp_cfg_x_5 <=_newCfg_WIRE_5[2];
              reg_pmp_cfg_w_5 <=_newCfg_WIRE_5[1]&_newCfg_WIRE_5[0];
              reg_pmp_cfg_r_5 <=_newCfg_WIRE_5[0];
            end 
         if (_GEN_30)
            begin 
              reg_pmp_cfg_x_6 <=_newCfg_WIRE_6[2];
              reg_pmp_cfg_w_6 <=_newCfg_WIRE_6[1]&_newCfg_WIRE_6[0];
              reg_pmp_cfg_r_6 <=_newCfg_WIRE_6[0];
            end 
         if (_GEN_32)
            begin 
              reg_pmp_cfg_x_7 <=_newCfg_T_49[2];
              reg_pmp_cfg_w_7 <=_newCfg_T_49[1]&_newCfg_T_49[0];
              reg_pmp_cfg_r_7 <=_newCfg_T_49[0];
            end 
         if (_csr_wen_T_4&(&_decoded_decoded_T_82)&~(reg_pmp_cfg_l_0|reg_pmp_cfg_l_1&~(reg_pmp_cfg_a_1[1])&reg_pmp_cfg_a_1[0]))
            reg_pmp_addr_0 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_84)&~(reg_pmp_cfg_l_1|reg_pmp_cfg_l_2&~(reg_pmp_cfg_a_2[1])&reg_pmp_cfg_a_2[0]))
            reg_pmp_addr_1 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_86)&~(reg_pmp_cfg_l_2|reg_pmp_cfg_l_3&~(reg_pmp_cfg_a_3[1])&reg_pmp_cfg_a_3[0]))
            reg_pmp_addr_2 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_88)&~(reg_pmp_cfg_l_3|reg_pmp_cfg_l_4&~(reg_pmp_cfg_a_4[1])&reg_pmp_cfg_a_4[0]))
            reg_pmp_addr_3 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_90)&~(reg_pmp_cfg_l_4|reg_pmp_cfg_l_5&~(reg_pmp_cfg_a_5[1])&reg_pmp_cfg_a_5[0]))
            reg_pmp_addr_4 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_92)&~(reg_pmp_cfg_l_5|reg_pmp_cfg_l_6&~(reg_pmp_cfg_a_6[1])&reg_pmp_cfg_a_6[0]))
            reg_pmp_addr_5 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_94)&~(reg_pmp_cfg_l_6|_GEN_31))
            reg_pmp_addr_6 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_96)&~(reg_pmp_cfg_l_7|_GEN_31))
            reg_pmp_addr_7 <=_GEN_24;
         if (_csr_wen_T_4&(&_decoded_decoded_T_4))
            reg_mie <={48'h0,_wdata_T_2[15:0]&_wdata_T_6[15:0]&16'h888};
         if (_csr_wen_T_4&(&_decoded_decoded_T_70))
            reg_mepc <=_GEN_20;
          else 
            if (_GEN_19)
               begin 
               end 
             else 
               reg_mepc <=epc;
         if (_csr_wen_T_4&(&_decoded_decoded_T_74))
            reg_mtval <=_wdata_T_2[33:0]&_wdata_T_6[33:0];
          else 
            if (_GEN_19)
               begin 
               end 
             else 
               reg_mtval <=insn_break ? epc:io_tval;
         if (_csr_wen_T_4&(&_decoded_decoded_T_68))
            reg_mscratch <=wdata;
       end
  
   wire [6:0] nextSmall_1={1'h0,small_1}+{6'h0,~io_csr_stall_0} ;  
  always @( posedge io_ungated_clock)
       begin 
         if (reset)
            begin 
              reg_wfi <=1'h0;
              small_1 <=6'h0;
              large_1 <=58'h0;
            end 
          else 
            begin 
              reg_wfi <=~((|{_GEN[11],_GEN[7],_GEN[3]})|io_interrupts_debug|exception)&(system_insn&(&{io_rw_addr[8],_GEN_11[9],_GEN_11[10],_GEN_11[11]})&~io_singleStep_0&~reg_debug|reg_wfi);
              if (_csr_wen_T_4&(&_decoded_decoded_T_130))
                 begin 
                   small_1 <=_GEN_16;
                   large_1 <=_wdata_T_2[63:6]&_wdata_T_6[63:6];
                 end 
               else 
                 begin 
                   if (reg_mcountinhibit[0])
                      begin 
                      end 
                    else 
                      small_1 <=nextSmall_1[5:0];
                   if (nextSmall_1[6]&~(reg_mcountinhibit[0]))
                      large_1 <=large_1+58'h1;
                 end 
            end 
       end
  
  assign io_rw_rdata=_io_rw_rdata_T_262; 
  assign io_decode_0_read_illegal=~csr_exists|(&{io_decode_0_inst[24],io_decode_0_inst[25],io_decode_0_read_illegal_invInputs[0],io_decode_0_inst[27],io_decode_0_inst[28],io_decode_0_inst[29],io_decode_0_inst[30],io_decode_0_read_illegal_invInputs[5]})&~reg_debug; 
  assign io_decode_0_write_illegal=&(io_decode_0_inst[31:30]); 
  assign io_decode_0_write_flush=~(io_decode_0_write_flush_addr_m>12'h33F&io_decode_0_write_flush_addr_m<12'h344); 
  assign io_decode_0_system_illegal=(|{&{decoded_invInputs_1[0],decoded_invInputs_1[1],decoded_invInputs_1[2],decoded_invInputs_1[3],decoded_invInputs_1[4],decoded_invInputs_1[5],io_decode_0_inst[28],io_decode_0_inst[29],decoded_invInputs_1[8],decoded_invInputs_1[9]},&{io_decode_0_inst[30],decoded_invInputs_1[9]}})&io_decode_0_inst[30]&io_decode_0_inst[27]&~reg_debug; 
  assign io_decode_0_virtual_access_illegal=reg_mstatus_v&csr_exists&(io_decode_0_inst[29:28]==2'h2|(io_decode_0_inst[31:20]>12'hBFF&io_decode_0_inst[31:20]<12'hC20|io_decode_0_inst[31:20]>12'hC7F&io_decode_0_inst[31:20]<12'hCA0)&_io_decode_0_virtual_access_illegal_T_3[0]&~(_io_decode_0_virtual_access_illegal_T_6[0])); 
  assign io_decode_0_virtual_system_illegal=1'h0; 
  assign io_csr_stall=io_csr_stall_0; 
  assign io_eret=_exception_T|insn_ret; 
  assign io_singleStep=io_singleStep_0; 
  assign io_status_debug=reg_debug; 
  assign io_status_wfi=reg_wfi; 
  assign io_status_isa=reg_misa[31:0]; 
  assign io_status_dv=reg_mstatus_v; 
  assign io_status_v=reg_mstatus_v; 
  assign io_evec=insn_ret ? (_GEN_14 ? ~{_io_evec_T_10[33:2],_io_evec_T_10[1:0]|{~(reg_misa[2]),1'h1}}:~{_io_evec_T_20[33:2],_io_evec_T_20[1:0]|{~(reg_misa[2]),1'h1}}):trapToDebug ? {22'h0,reg_debug ? {8'h80,~insn_break,3'h0}:12'h800}:{2'h0,_read_mtvec_T_5[0]&cause[63]&cause[7:6]==2'h0 ? {_read_mtvec_T_5[31:8],cause[5:0]}:_read_mtvec_T_5[31:2],2'h0}; 
  assign io_time=io_time_0; 
  assign io_interrupt=((io_interrupts_debug|m_interrupts[15]|m_interrupts[14]|m_interrupts[13]|m_interrupts[12]|m_interrupts[11]|m_interrupts[3]|m_interrupts[7]|m_interrupts[9]|m_interrupts[1]|m_interrupts[5]|m_interrupts[10]|m_interrupts[2]|m_interrupts[6]|m_interrupts[8]|m_interrupts[0]|m_interrupts[4])&~io_singleStep_0|reg_singleStepped)&~(reg_debug|io_status_cease_r); 
  assign io_interrupt_cause={60'h0,io_interrupts_debug ? 4'hE:m_interrupts[15] ? 4'hF:m_interrupts[14] ? 4'hE:m_interrupts[13] ? 4'hD:m_interrupts[12] ? 4'hC:m_interrupts[11] ? 4'hB:m_interrupts[3] ? 4'h3:m_interrupts[7] ? 4'h7:m_interrupts[9] ? 4'h9:m_interrupts[1] ? 4'h1:m_interrupts[5] ? 4'h5:m_interrupts[10] ? 4'hA:m_interrupts[2] ? 4'h2:m_interrupts[6] ? 4'h6:m_interrupts[8] ? 4'h8:{1'h0,~(m_interrupts[0]),2'h0}}-64'h8000000000000000; 
  assign io_bp_0_control_action=reg_bp_0_control_action; 
  assign io_bp_0_control_tmatch=reg_bp_0_control_tmatch; 
  assign io_bp_0_control_x=reg_bp_0_control_x; 
  assign io_bp_0_control_w=reg_bp_0_control_w; 
  assign io_bp_0_control_r=reg_bp_0_control_r; 
  assign io_bp_0_address=reg_bp_0_address; 
  assign io_pmp_cfg_l_0=reg_pmp_cfg_l_0; 
  assign io_pmp_cfg_l_1=reg_pmp_cfg_l_1; 
  assign io_pmp_cfg_l_2=reg_pmp_cfg_l_2; 
  assign io_pmp_cfg_l_3=reg_pmp_cfg_l_3; 
  assign io_pmp_cfg_l_4=reg_pmp_cfg_l_4; 
  assign io_pmp_cfg_l_5=reg_pmp_cfg_l_5; 
  assign io_pmp_cfg_l_6=reg_pmp_cfg_l_6; 
  assign io_pmp_cfg_l_7=reg_pmp_cfg_l_7; 
  assign io_pmp_cfg_a_0=reg_pmp_cfg_a_0; 
  assign io_pmp_cfg_a_1=reg_pmp_cfg_a_1; 
  assign io_pmp_cfg_a_2=reg_pmp_cfg_a_2; 
  assign io_pmp_cfg_a_3=reg_pmp_cfg_a_3; 
  assign io_pmp_cfg_a_4=reg_pmp_cfg_a_4; 
  assign io_pmp_cfg_a_5=reg_pmp_cfg_a_5; 
  assign io_pmp_cfg_a_6=reg_pmp_cfg_a_6; 
  assign io_pmp_cfg_a_7=reg_pmp_cfg_a_7; 
  assign io_pmp_cfg_x_0=reg_pmp_cfg_x_0; 
  assign io_pmp_cfg_x_1=reg_pmp_cfg_x_1; 
  assign io_pmp_cfg_x_2=reg_pmp_cfg_x_2; 
  assign io_pmp_cfg_x_3=reg_pmp_cfg_x_3; 
  assign io_pmp_cfg_x_4=reg_pmp_cfg_x_4; 
  assign io_pmp_cfg_x_5=reg_pmp_cfg_x_5; 
  assign io_pmp_cfg_x_6=reg_pmp_cfg_x_6; 
  assign io_pmp_cfg_x_7=reg_pmp_cfg_x_7; 
  assign io_pmp_cfg_w_0=reg_pmp_cfg_w_0; 
  assign io_pmp_cfg_w_1=reg_pmp_cfg_w_1; 
  assign io_pmp_cfg_w_2=reg_pmp_cfg_w_2; 
  assign io_pmp_cfg_w_3=reg_pmp_cfg_w_3; 
  assign io_pmp_cfg_w_4=reg_pmp_cfg_w_4; 
  assign io_pmp_cfg_w_5=reg_pmp_cfg_w_5; 
  assign io_pmp_cfg_w_6=reg_pmp_cfg_w_6; 
  assign io_pmp_cfg_w_7=reg_pmp_cfg_w_7; 
  assign io_pmp_cfg_r_0=reg_pmp_cfg_r_0; 
  assign io_pmp_cfg_r_1=reg_pmp_cfg_r_1; 
  assign io_pmp_cfg_r_2=reg_pmp_cfg_r_2; 
  assign io_pmp_cfg_r_3=reg_pmp_cfg_r_3; 
  assign io_pmp_cfg_r_4=reg_pmp_cfg_r_4; 
  assign io_pmp_cfg_r_5=reg_pmp_cfg_r_5; 
  assign io_pmp_cfg_r_6=reg_pmp_cfg_r_6; 
  assign io_pmp_cfg_r_7=reg_pmp_cfg_r_7; 
  assign io_pmp_addr_0=reg_pmp_addr_0; 
  assign io_pmp_addr_1=reg_pmp_addr_1; 
  assign io_pmp_addr_2=reg_pmp_addr_2; 
  assign io_pmp_addr_3=reg_pmp_addr_3; 
  assign io_pmp_addr_4=reg_pmp_addr_4; 
  assign io_pmp_addr_5=reg_pmp_addr_5; 
  assign io_pmp_addr_6=reg_pmp_addr_6; 
  assign io_pmp_addr_7=reg_pmp_addr_7; 
  assign io_pmp_mask_0={_GEN_0&~(_GEN_0+30'h1),2'h3}; 
  assign io_pmp_mask_1={_GEN_1&~(_GEN_1+30'h1),2'h3}; 
  assign io_pmp_mask_2={_GEN_2&~(_GEN_2+30'h1),2'h3}; 
  assign io_pmp_mask_3={_GEN_3&~(_GEN_3+30'h1),2'h3}; 
  assign io_pmp_mask_4={_GEN_4&~(_GEN_4+30'h1),2'h3}; 
  assign io_pmp_mask_5={_GEN_5&~(_GEN_5+30'h1),2'h3}; 
  assign io_pmp_mask_6={_GEN_6&~(_GEN_6+30'h1),2'h3}; 
  assign io_pmp_mask_7={_GEN_7&~(_GEN_7+30'h1),2'h3}; 
  assign io_inhibit_cycle=reg_mcountinhibit[0]; 
  assign io_trace_valid_0=io_retire|exception; 
  assign io_trace_iaddr_0=io_pc; 
  assign io_trace_insn_0=io_inst_0; 
  assign io_trace_exception_0=exception; 
  assign io_customCSRs_0_value=reg_custom_0; 
endmodule
 
module BreakpointUnit (
  input io_status_debug,
  input io_bp_0_control_action,
  input [1:0] io_bp_0_control_tmatch,
  input io_bp_0_control_x,
  input io_bp_0_control_w,
  input io_bp_0_control_r,
  input [32:0] io_bp_0_address,
  input [32:0] io_pc,
  input [32:0] io_ea,
  output io_xcpt_if,
  output io_xcpt_ld,
  output io_xcpt_st,
  output io_debug_if,
  output io_debug_ld,
  output io_debug_st) ; 
   wire _w_T_2=io_ea>=io_bp_0_address ;  
   wire [32:0] _w_T_5=~io_ea ;  
   wire _r_T_8=io_bp_0_control_tmatch[0]&io_bp_0_address[0] ;  
   wire _r_T_10=_r_T_8&io_bp_0_address[1] ;  
   wire [32:0] _x_T_15=~io_bp_0_address ;  
   wire _r_T_18=io_bp_0_control_tmatch[0]&io_bp_0_address[0] ;  
   wire _r_T_20=_r_T_18&io_bp_0_address[1] ;  
   wire r=~io_status_debug&io_bp_0_control_r&(io_bp_0_control_tmatch[1] ? _w_T_2^io_bp_0_control_tmatch[0]:{_w_T_5[32:4],_w_T_5[3:0]|{_r_T_10&io_bp_0_address[2],_r_T_10,_r_T_8,io_bp_0_control_tmatch[0]}}=={_x_T_15[32:4],_x_T_15[3:0]|{_r_T_20&io_bp_0_address[2],_r_T_20,_r_T_18,io_bp_0_control_tmatch[0]}}) ;  
   wire _w_T_8=io_bp_0_control_tmatch[0]&io_bp_0_address[0] ;  
   wire _w_T_10=_w_T_8&io_bp_0_address[1] ;  
   wire _w_T_18=io_bp_0_control_tmatch[0]&io_bp_0_address[0] ;  
   wire _w_T_20=_w_T_18&io_bp_0_address[1] ;  
   wire w=~io_status_debug&io_bp_0_control_w&(io_bp_0_control_tmatch[1] ? _w_T_2^io_bp_0_control_tmatch[0]:{_w_T_5[32:4],_w_T_5[3:0]|{_w_T_10&io_bp_0_address[2],_w_T_10,_w_T_8,io_bp_0_control_tmatch[0]}}=={_x_T_15[32:4],_x_T_15[3:0]|{_w_T_20&io_bp_0_address[2],_w_T_20,_w_T_18,io_bp_0_control_tmatch[0]}}) ;  
   wire [32:0] _x_T_5=~io_pc ;  
   wire _x_T_8=io_bp_0_control_tmatch[0]&io_bp_0_address[0] ;  
   wire _x_T_10=_x_T_8&io_bp_0_address[1] ;  
   wire _x_T_18=io_bp_0_control_tmatch[0]&io_bp_0_address[0] ;  
   wire _x_T_20=_x_T_18&io_bp_0_address[1] ;  
   wire x=~io_status_debug&io_bp_0_control_x&(io_bp_0_control_tmatch[1] ? io_pc>=io_bp_0_address^io_bp_0_control_tmatch[0]:{_x_T_5[32:4],_x_T_5[3:0]|{_x_T_10&io_bp_0_address[2],_x_T_10,_x_T_8,io_bp_0_control_tmatch[0]}}=={_x_T_15[32:4],_x_T_15[3:0]|{_x_T_20&io_bp_0_address[2],_x_T_20,_x_T_18,io_bp_0_control_tmatch[0]}}) ;  
  assign io_xcpt_if=x&~io_bp_0_control_action; 
  assign io_xcpt_ld=r&~io_bp_0_control_action; 
  assign io_xcpt_st=w&~io_bp_0_control_action; 
  assign io_debug_if=x&io_bp_0_control_action; 
  assign io_debug_ld=r&io_bp_0_control_action; 
  assign io_debug_st=w&io_bp_0_control_action; 
endmodule
 
module ALU (
  input io_dw,
  input [3:0] io_fn,
  input [63:0] io_in2,
  input [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output io_cmp_out) ; 
   wire [63:0] in2_inv={64{io_fn[3]}}^io_in2 ;  
   wire [63:0] in1_xor_in2=io_in1^in2_inv ;  
   wire [63:0] _io_adder_out_T_3=io_in1+in2_inv+{63'h0,io_fn[3]} ;  
   wire slt=io_in1[63]==io_in2[63] ? _io_adder_out_T_3[63]:io_fn[1] ? io_in2[63]:io_in1[63] ;  
   wire [31:0] shin_hi=io_dw ? io_in1[63:32]:{32{io_fn[3]&io_in1[31]}} ;  
   wire _shout_T=io_fn==4'h5 ;  
   wire _shout_T_1=io_fn==4'hB ;  
   wire [31:0] _GEN={io_in1[31:16],16'h0}|shin_hi&32'hFFFF ;  
   wire [31:0] _GEN_0={{io_in1[15:0],_GEN[31:24]}&24'hFF00FF,8'h0}|_GEN&32'hFF00FF ;  
   wire [31:0] _GEN_1={{io_in1[7:0],_GEN_0[31:12]}&28'hF0F0F0F,4'h0}|_GEN_0&32'hF0F0F0F ;  
   wire [45:0] _GEN_2={io_in1[3:0],_GEN_1,_GEN_0[7:4],_GEN[11:8],_GEN[15:14]}&46'h333333333333 ;  
   wire [31:0] _GEN_3=_GEN_2[45:14]|_GEN_1&32'h33333333 ;  
   wire [1:0] _GEN_4=_GEN_2[11:10]|_GEN_0[5:4] ;  
   wire [7:0] _GEN_5={_GEN_2[5:0],2'h0}|{_GEN[15:12],shin_hi[19:16]}&8'h33 ;  
   wire [54:0] _GEN_6={io_in1[1:0],_GEN_3,_GEN_1[3:2],_GEN_4,_GEN_0[7:6],_GEN[9:8],_GEN_5,shin_hi[19:18],shin_hi[21:20],shin_hi[23]}&55'h55555555555555 ;  
   wire [63:0] shin=_shout_T|_shout_T_1 ? {shin_hi,io_in1[31:0]}:{io_in1[0],_GEN_6[54:23]|_GEN_3&32'h55555555,_GEN_3[1],_GEN_6[21]|_GEN_1[2],{_GEN_1[3],1'h0}|_GEN_4&2'h1,_GEN_6[18:15]|{_GEN_0[7:6],_GEN[9:8]}&4'h5,_GEN_6[14:7]|_GEN_5&8'h55,_GEN_5[1],_GEN_6[5]|shin_hi[18],shin_hi[19],shin_hi[20],{_GEN_6[2:0],1'h0}|{shin_hi[23:22],shin_hi[25:24]}&4'h5,shin_hi[25],shin_hi[26],shin_hi[27],shin_hi[28],shin_hi[29],shin_hi[30],shin_hi[31]} ;  
   wire [64:0] _shout_r_T_5=$signed($signed({io_fn[3]&shin[63],shin})>>>{59'h0,io_in2[5]&io_dw,io_in2[4:0]}) ;  
   wire [15:0] _GEN_7={{_shout_r_T_5[23:16],_shout_r_T_5[31:28]}&12'hF0F,4'h0}|{_shout_r_T_5[31:24],_shout_r_T_5[39:32]}&16'hF0F ;  
   wire [37:0] _GEN_8={_shout_r_T_5[11:8],_shout_r_T_5[15:12],_shout_r_T_5[19:16],_GEN_7,_shout_r_T_5[39:36],_shout_r_T_5[43:40],_shout_r_T_5[47:46]}&38'h3333333333 ;  
   wire [7:0] _GEN_9=_GEN_8[37:30]|{_shout_r_T_5[15:12],_shout_r_T_5[19:16]}&8'h33 ;  
   wire [15:0] _GEN_10=_GEN_8[29:14]|_GEN_7&16'h3333 ;  
   wire [1:0] _GEN_11=_GEN_8[11:10]|_shout_r_T_5[37:36] ;  
   wire [7:0] _GEN_12={_GEN_8[5:0],2'h0}|{_shout_r_T_5[47:44],_shout_r_T_5[51:48]}&8'h33 ;  
   wire [50:0] _GEN_13={_shout_r_T_5[5:4],_shout_r_T_5[7:6],_shout_r_T_5[9:8],_GEN_9,_GEN_10,_GEN_7[3:2],_GEN_11,_shout_r_T_5[39:38],_shout_r_T_5[41:40],_GEN_12,_shout_r_T_5[51:50],_shout_r_T_5[53:52],_shout_r_T_5[55]}&51'h5555555555555 ;  
   wire _logic_T_4=io_fn==4'h6 ;  
   wire [63:0] out=io_fn==4'h0|io_fn==4'hA ? _io_adder_out_T_3:{63'h0,io_fn>4'hB&slt}|(io_fn==4'h4|_logic_T_4 ? in1_xor_in2:64'h0)|(_logic_T_4|io_fn==4'h7 ? io_in1&io_in2:64'h0)|(_shout_T|_shout_T_1 ? _shout_r_T_5[63:0]:64'h0)|(io_fn==4'h1 ? {_shout_r_T_5[0],_shout_r_T_5[1],_shout_r_T_5[2],_shout_r_T_5[3],_shout_r_T_5[4],_GEN_13[50:47]|{_shout_r_T_5[7:6],_shout_r_T_5[9:8]}&4'h5,_GEN_13[46:39]|_GEN_9&8'h55,_GEN_13[38:23]|_GEN_10&16'h5555,_GEN_10[1],_GEN_13[21]|_GEN_7[2],{_GEN_7[3],1'h0}|_GEN_11&2'h1,_GEN_13[18:15]|{_shout_r_T_5[39:38],_shout_r_T_5[41:40]}&4'h5,_GEN_13[14:7]|_GEN_12&8'h55,_GEN_12[1],_GEN_13[5]|_shout_r_T_5[50],_shout_r_T_5[51],_shout_r_T_5[52],{_GEN_13[2:0],1'h0}|{_shout_r_T_5[55:54],_shout_r_T_5[57:56]}&4'h5,_shout_r_T_5[57],_shout_r_T_5[58],_shout_r_T_5[59],_shout_r_T_5[60],_shout_r_T_5[61],_shout_r_T_5[62],_shout_r_T_5[63]}:64'h0) ;  
  assign io_out=io_dw ? out:{{32{out[31]}},out[31:0]}; 
  assign io_adder_out=_io_adder_out_T_3; 
  assign io_cmp_out=io_fn[0]^(io_fn[3] ? slt:in1_xor_in2==64'h0); 
endmodule
 
module MulDiv (
  input clock,
  input reset,
  output io_req_ready,
  input io_req_valid,
  input [3:0] io_req_bits_fn,
  input io_req_bits_dw,
  input [63:0] io_req_bits_in1,
  input [63:0] io_req_bits_in2,
  input [4:0] io_req_bits_tag,
  input io_kill,
  input io_resp_ready,
  output io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0] io_resp_bits_tag) ; 
   reg [2:0] state ;  
   reg req_dw ;  
   reg [4:0] req_tag ;  
   reg [6:0] count ;  
   reg neg_out ;  
   reg isHi ;  
   reg resHi ;  
   reg [64:0] divisor ;  
   reg [129:0] remainder ;  
   wire [63:0] result=resHi ? remainder[128:65]:remainder[63:0] ;  
   wire [31:0] loOut=req_dw|state[0] ? result[31:0]:result[63:32] ;  
   wire io_resp_valid_0=state==3'h6|(&state) ;  
   wire io_req_ready_0=state==3'h0 ;  
   wire [65:0] _prod_T_4={{65{remainder[64]}},remainder[0]}*{divisor[64],divisor}+{remainder[129],remainder[129:65]} ;  
   wire [64:0] _subtractor_T_1=remainder[128:64]-divisor ;  
   wire [2:0] decoded_invInputs=~(io_req_bits_fn[2:0]) ;  
   wire [1:0] _decoded_T_2={decoded_invInputs[1],decoded_invInputs[2]} ;  
   wire lhs_sign=(|{decoded_invInputs[0],&_decoded_T_2})&(io_req_bits_dw ? io_req_bits_in1[63]:io_req_bits_in1[31]) ;  
   wire rhs_sign=(|{&_decoded_T_2,&{decoded_invInputs[0],io_req_bits_fn[2]}})&(io_req_bits_dw ? io_req_bits_in2[63]:io_req_bits_in2[31]) ;  
   wire _GEN=state==3'h1 ;  
   wire _GEN_0=state==3'h5 ;  
   wire _GEN_1=state==3'h2 ;  
   wire _GEN_2=_GEN_1&count==7'h3F ;  
   wire _GEN_3=state==3'h3 ;  
   wire _GEN_4=count==7'h40 ;  
   wire _GEN_5=io_req_ready_0&io_req_valid ;  
   wire [1:0] _decoded_orMatrixOutputs_T_4={&{io_req_bits_fn[0],decoded_invInputs[2]},io_req_bits_fn[1]} ;  
  always @( posedge clock)
       begin 
         if (reset)
            state <=3'h0;
          else 
            if (_GEN_5)
               state <=decoded_invInputs[2] ? 3'h2:{1'h0,~(lhs_sign|rhs_sign),1'h1};
             else 
               if (io_resp_ready&io_resp_valid_0|io_kill)
                  state <=3'h0;
                else 
                  if (_GEN_3&_GEN_4)
                     state <={1'h1,~neg_out,1'h1};
                   else 
                     if (_GEN_2)
                        state <=3'h6;
                      else 
                        if (_GEN_0)
                           state <=3'h7;
                         else 
                           if (_GEN)
                              state <=3'h3;
         if (_GEN_5)
            begin 
              req_dw <=io_req_bits_dw;
              req_tag <=io_req_bits_tag;
              count <={1'h0,decoded_invInputs[2]&~io_req_bits_dw,5'h0};
              neg_out <=(|_decoded_orMatrixOutputs_T_4) ? lhs_sign:lhs_sign!=rhs_sign;
              isHi <=|_decoded_orMatrixOutputs_T_4;
              divisor <={rhs_sign,io_req_bits_dw ? io_req_bits_in2[63:32]:{32{rhs_sign}},io_req_bits_in2[31:0]};
              remainder <={66'h0,io_req_bits_dw ? io_req_bits_in1[63:32]:{32{lhs_sign}},io_req_bits_in1[31:0]};
            end 
          else 
            begin 
              if (_GEN_3)
                 begin 
                   count <=count+7'h1;
                   remainder <={1'h0,_subtractor_T_1[64] ? remainder[127:64]:_subtractor_T_1[63:0],remainder[63:0],~(_subtractor_T_1[64])};
                 end 
               else 
                 if (_GEN_1)
                    begin 
                      count <=count+7'h1;
                      remainder <={_prod_T_4[65:1],count==7'h3E&neg_out,_prod_T_4[0],remainder[63:1]};
                    end 
                  else 
                    if (_GEN_0|_GEN&remainder[63])
                       remainder <={66'h0,64'h0-result};
              neg_out <=~(_GEN_3&count==7'h0&~(_subtractor_T_1[64])&~isHi)&neg_out;
              if (_GEN&divisor[63])
                 divisor <=_subtractor_T_1;
            end 
         resHi <=~_GEN_5&(_GEN_3&_GEN_4|_GEN_2 ? isHi:~_GEN_0&resHi);
       end
  
  assign io_req_ready=io_req_ready_0; 
  assign io_resp_valid=io_resp_valid_0; 
  assign io_resp_bits_data={req_dw ? result[63:32]:{32{loOut[31]}},loOut}; 
  assign io_resp_bits_tag=req_tag; 
endmodule
 
module PlusArgTimeout (
  input clock,
  input reset,
  input [31:0] io_count) ; 
   wire [31:0] _plusarg_reader_out ;  
  always @( posedge clock)
       begin 
         if ((|_plusarg_reader_out)&~reset&io_count>=_plusarg_reader_out)
            begin 
              if (1)$display("Assertion failed: Timeout exceeded: Kill the emulation after INT rdtime cycles. Off if 0.\n    at PlusArg.scala:64 assert (io.count < max, s\"Timeout exceeded: $docstring\")\n");
              if (1)$display("");
            end 
       end
  
endmodule
 
module rf_31x64 (
  input [4:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [63:0] R0_data,
  input [4:0] R1_addr,
  input R1_en,
  input R1_clk,
  output [63:0] R1_data,
  input [4:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [63:0] W0_data) ; 
   reg [63:0] Memory[0:30] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:64'bx; 
  assign R1_data=R1_en ? Memory[R1_addr]:64'bx; 
endmodule
 
module Rocket (
  input clock,
  input reset,
  input io_hartid,
  input io_interrupts_debug,
  input io_interrupts_mtip,
  input io_interrupts_msip,
  input io_interrupts_meip,
  output io_imem_might_request,
  output io_imem_req_valid,
  output [33:0] io_imem_req_bits_pc,
  output io_imem_req_bits_speculative,
  output io_imem_resp_ready,
  input io_imem_resp_valid,
  input [33:0] io_imem_resp_bits_pc,
  input [31:0] io_imem_resp_bits_data,
  input io_imem_resp_bits_xcpt_pf_inst,
  input io_imem_resp_bits_xcpt_gf_inst,
  input io_imem_resp_bits_xcpt_ae_inst,
  input io_imem_resp_bits_replay,
  output io_imem_btb_update_valid,
  output io_imem_bht_update_valid,
  output io_imem_flush_icache,
  input io_dmem_req_ready,
  output io_dmem_req_valid,
  output [33:0] io_dmem_req_bits_addr,
  output [5:0] io_dmem_req_bits_tag,
  output [4:0] io_dmem_req_bits_cmd,
  output [1:0] io_dmem_req_bits_size,
  output io_dmem_req_bits_signed,
  output io_dmem_req_bits_dv,
  output io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data_data,
  input io_dmem_s2_nack,
  input io_dmem_resp_valid,
  input [5:0] io_dmem_resp_bits_tag,
  input [63:0] io_dmem_resp_bits_data,
  input io_dmem_resp_bits_replay,
  input io_dmem_resp_bits_has_data,
  input [63:0] io_dmem_resp_bits_data_word_bypass,
  input io_dmem_replay_next,
  input io_dmem_s2_xcpt_ma_ld,
  input io_dmem_s2_xcpt_ma_st,
  input io_dmem_s2_xcpt_pf_ld,
  input io_dmem_s2_xcpt_pf_st,
  input io_dmem_s2_xcpt_ae_ld,
  input io_dmem_s2_xcpt_ae_st,
  input io_dmem_ordered,
  input io_dmem_perf_release,
  input io_dmem_perf_grant,
  output io_ptw_status_debug,
  output io_ptw_pmp_cfg_l_0,
  output io_ptw_pmp_cfg_l_1,
  output io_ptw_pmp_cfg_l_2,
  output io_ptw_pmp_cfg_l_3,
  output io_ptw_pmp_cfg_l_4,
  output io_ptw_pmp_cfg_l_5,
  output io_ptw_pmp_cfg_l_6,
  output io_ptw_pmp_cfg_l_7,
  output [1:0] io_ptw_pmp_cfg_a_0,
  output [1:0] io_ptw_pmp_cfg_a_1,
  output [1:0] io_ptw_pmp_cfg_a_2,
  output [1:0] io_ptw_pmp_cfg_a_3,
  output [1:0] io_ptw_pmp_cfg_a_4,
  output [1:0] io_ptw_pmp_cfg_a_5,
  output [1:0] io_ptw_pmp_cfg_a_6,
  output [1:0] io_ptw_pmp_cfg_a_7,
  output io_ptw_pmp_cfg_x_0,
  output io_ptw_pmp_cfg_x_1,
  output io_ptw_pmp_cfg_x_2,
  output io_ptw_pmp_cfg_x_3,
  output io_ptw_pmp_cfg_x_4,
  output io_ptw_pmp_cfg_x_5,
  output io_ptw_pmp_cfg_x_6,
  output io_ptw_pmp_cfg_x_7,
  output io_ptw_pmp_cfg_w_0,
  output io_ptw_pmp_cfg_w_1,
  output io_ptw_pmp_cfg_w_2,
  output io_ptw_pmp_cfg_w_3,
  output io_ptw_pmp_cfg_w_4,
  output io_ptw_pmp_cfg_w_5,
  output io_ptw_pmp_cfg_w_6,
  output io_ptw_pmp_cfg_w_7,
  output io_ptw_pmp_cfg_r_0,
  output io_ptw_pmp_cfg_r_1,
  output io_ptw_pmp_cfg_r_2,
  output io_ptw_pmp_cfg_r_3,
  output io_ptw_pmp_cfg_r_4,
  output io_ptw_pmp_cfg_r_5,
  output io_ptw_pmp_cfg_r_6,
  output io_ptw_pmp_cfg_r_7,
  output [29:0] io_ptw_pmp_addr_0,
  output [29:0] io_ptw_pmp_addr_1,
  output [29:0] io_ptw_pmp_addr_2,
  output [29:0] io_ptw_pmp_addr_3,
  output [29:0] io_ptw_pmp_addr_4,
  output [29:0] io_ptw_pmp_addr_5,
  output [29:0] io_ptw_pmp_addr_6,
  output [29:0] io_ptw_pmp_addr_7,
  output [31:0] io_ptw_pmp_mask_0,
  output [31:0] io_ptw_pmp_mask_1,
  output [31:0] io_ptw_pmp_mask_2,
  output [31:0] io_ptw_pmp_mask_3,
  output [31:0] io_ptw_pmp_mask_4,
  output [31:0] io_ptw_pmp_mask_5,
  output [31:0] io_ptw_pmp_mask_6,
  output [31:0] io_ptw_pmp_mask_7,
  output [63:0] io_ptw_customCSRs_csrs_0_value,
  output io_wfi) ; 
   wire io_dmem_req_valid_0 ;  
   wire div_io_resp_ready ;  
   wire take_pc_wb ;  
   wire take_pc_mem ;  
   wire _div_io_req_ready ;  
   wire _div_io_resp_valid ;  
   wire [63:0] _div_io_resp_bits_data ;  
   wire [4:0] _div_io_resp_bits_tag ;  
   wire [63:0] _alu_io_out ;  
   wire [63:0] _alu_io_adder_out ;  
   wire _alu_io_cmp_out ;  
   wire _bpu_io_xcpt_if ;  
   wire _bpu_io_xcpt_ld ;  
   wire _bpu_io_xcpt_st ;  
   wire _bpu_io_debug_if ;  
   wire _bpu_io_debug_ld ;  
   wire _bpu_io_debug_st ;  
   wire [63:0] _csr_io_rw_rdata ;  
   wire _csr_io_decode_0_read_illegal ;  
   wire _csr_io_decode_0_write_illegal ;  
   wire _csr_io_decode_0_write_flush ;  
   wire _csr_io_decode_0_system_illegal ;  
   wire _csr_io_decode_0_virtual_access_illegal ;  
   wire _csr_io_decode_0_virtual_system_illegal ;  
   wire _csr_io_csr_stall ;  
   wire _csr_io_eret ;  
   wire _csr_io_singleStep ;  
   wire _csr_io_status_debug ;  
   wire [31:0] _csr_io_status_isa ;  
   wire _csr_io_status_dv ;  
   wire _csr_io_status_v ;  
   wire [33:0] _csr_io_evec ;  
   wire [63:0] _csr_io_time ;  
   wire _csr_io_interrupt ;  
   wire [63:0] _csr_io_interrupt_cause ;  
   wire _csr_io_bp_0_control_action ;  
   wire [1:0] _csr_io_bp_0_control_tmatch ;  
   wire _csr_io_bp_0_control_x ;  
   wire _csr_io_bp_0_control_w ;  
   wire _csr_io_bp_0_control_r ;  
   wire [32:0] _csr_io_bp_0_address ;  
   wire _csr_io_inhibit_cycle ;  
   wire _csr_io_trace_valid_0 ;  
   wire [33:0] _csr_io_trace_iaddr_0 ;  
   wire [31:0] _csr_io_trace_insn_0 ;  
   wire _csr_io_trace_exception_0 ;  
   wire [63:0] _csr_io_customCSRs_0_value ;  
   wire [63:0] _rf_ext_R0_data ;  
   wire [63:0] _rf_ext_R1_data ;  
   wire [33:0] _ibuf_io_pc ;  
   wire _ibuf_io_inst_0_valid ;  
   wire _ibuf_io_inst_0_bits_xcpt0_pf_inst ;  
   wire _ibuf_io_inst_0_bits_xcpt0_gf_inst ;  
   wire _ibuf_io_inst_0_bits_xcpt0_ae_inst ;  
   wire _ibuf_io_inst_0_bits_xcpt1_pf_inst ;  
   wire _ibuf_io_inst_0_bits_xcpt1_gf_inst ;  
   wire _ibuf_io_inst_0_bits_xcpt1_ae_inst ;  
   wire _ibuf_io_inst_0_bits_replay ;  
   wire _ibuf_io_inst_0_bits_rvc ;  
   wire [31:0] _ibuf_io_inst_0_bits_inst_bits ;  
   wire [4:0] _ibuf_io_inst_0_bits_inst_rd ;  
   wire [4:0] _ibuf_io_inst_0_bits_inst_rs1 ;  
   wire [4:0] _ibuf_io_inst_0_bits_inst_rs2 ;  
   wire [31:0] _ibuf_io_inst_0_bits_raw ;  
   reg id_reg_pause ;  
   reg imem_might_request_reg ;  
   reg ex_ctrl_fp ;  
   reg ex_ctrl_rocc ;  
   reg ex_ctrl_branch ;  
   reg ex_ctrl_jal ;  
   reg ex_ctrl_jalr ;  
   reg ex_ctrl_rxs2 ;  
   reg ex_ctrl_rxs1 ;  
   reg [1:0] ex_ctrl_sel_alu2 ;  
   reg [1:0] ex_ctrl_sel_alu1 ;  
   reg [2:0] ex_ctrl_sel_imm ;  
   reg ex_ctrl_alu_dw ;  
   reg [3:0] ex_ctrl_alu_fn ;  
   reg ex_ctrl_mem ;  
   reg [4:0] ex_ctrl_mem_cmd ;  
   reg ex_ctrl_rfs1 ;  
   reg ex_ctrl_rfs2 ;  
   reg ex_ctrl_wfd ;  
   reg ex_ctrl_mul ;  
   reg ex_ctrl_div ;  
   reg ex_ctrl_wxd ;  
   reg [2:0] ex_ctrl_csr ;  
   reg ex_ctrl_fence_i ;  
   reg mem_ctrl_fp ;  
   reg mem_ctrl_rocc ;  
   reg mem_ctrl_branch ;  
   reg mem_ctrl_jal ;  
   reg mem_ctrl_jalr ;  
   reg mem_ctrl_rxs2 ;  
   reg mem_ctrl_rxs1 ;  
   reg mem_ctrl_mem ;  
   reg mem_ctrl_rfs1 ;  
   reg mem_ctrl_rfs2 ;  
   reg mem_ctrl_wfd ;  
   reg mem_ctrl_mul ;  
   reg mem_ctrl_div ;  
   reg mem_ctrl_wxd ;  
   reg [2:0] mem_ctrl_csr ;  
   reg mem_ctrl_fence_i ;  
   reg wb_ctrl_rocc ;  
   reg wb_ctrl_rxs2 ;  
   reg wb_ctrl_rxs1 ;  
   reg wb_ctrl_mem ;  
   reg wb_ctrl_rfs1 ;  
   reg wb_ctrl_rfs2 ;  
   reg wb_ctrl_wfd ;  
   reg wb_ctrl_div ;  
   reg wb_ctrl_wxd ;  
   reg [2:0] wb_ctrl_csr ;  
   reg wb_ctrl_fence_i ;  
   reg ex_reg_xcpt_interrupt ;  
   reg ex_reg_valid ;  
   reg ex_reg_rvc ;  
   reg ex_reg_xcpt ;  
   reg ex_reg_flush_pipe ;  
   reg ex_reg_load_use ;  
   reg [63:0] ex_reg_cause ;  
   reg ex_reg_replay ;  
   reg [33:0] ex_reg_pc ;  
   reg [1:0] ex_reg_mem_size ;  
   reg [31:0] ex_reg_inst ;  
   reg [31:0] ex_reg_raw_inst ;  
   reg mem_reg_xcpt_interrupt ;  
   reg mem_reg_valid ;  
   reg mem_reg_rvc ;  
   reg mem_reg_xcpt ;  
   reg mem_reg_replay ;  
   reg mem_reg_flush_pipe ;  
   reg [63:0] mem_reg_cause ;  
   reg mem_mem_cmd_bh ;  
   reg mem_reg_load ;  
   reg mem_reg_store ;  
   reg [33:0] mem_reg_pc ;  
   reg [31:0] mem_reg_inst ;  
   reg mem_reg_hls_or_dv ;  
   reg [31:0] mem_reg_raw_inst ;  
   reg [63:0] mem_reg_wdata ;  
   reg [63:0] mem_reg_rs2 ;  
   reg mem_br_taken ;  
   reg wb_reg_valid ;  
   reg wb_reg_xcpt ;  
   reg wb_reg_replay ;  
   reg wb_reg_flush_pipe ;  
   reg [63:0] wb_reg_cause ;  
   reg [33:0] wb_reg_pc ;  
   reg wb_reg_hls_or_dv ;  
   reg [31:0] wb_reg_inst ;  
   reg [31:0] wb_reg_raw_inst ;  
   reg [63:0] wb_reg_wdata ;  
   wire ibuf_io_kill=take_pc_wb|take_pc_mem ;  
   wire [29:0] id_ctrl_decoder_decoded_invInputs=~(_ibuf_io_inst_0_bits_inst_bits[31:2]) ;  
   wire [6:0] _id_ctrl_decoder_decoded_T={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_4={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[11]} ;  
   wire [6:0] _id_ctrl_decoder_decoded_T_6={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_8={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [8:0] _id_ctrl_decoder_decoded_T_12={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [5:0] _id_ctrl_decoder_decoded_T_14={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[4]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_18={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [14:0] _id_ctrl_decoder_decoded_T_22={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [12:0] _id_ctrl_decoder_decoded_T_26={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [14:0] _id_ctrl_decoder_decoded_T_28={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [8:0] _id_ctrl_decoder_decoded_T_36={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [9:0] _id_ctrl_decoder_decoded_T_38={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [6:0] _id_ctrl_decoder_decoded_T_40={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6]} ;  
   wire [9:0] _id_ctrl_decoder_decoded_T_46={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [13:0] _id_ctrl_decoder_decoded_T_48={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [14:0] _id_ctrl_decoder_decoded_T_52={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[3],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [8:0] _id_ctrl_decoder_decoded_T_60={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_62={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[12]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_64={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13]} ;  
   wire [10:0] _id_ctrl_decoder_decoded_T_68={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_74={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[13]} ;  
   wire [8:0] _id_ctrl_decoder_decoded_T_76={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_86={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[14]} ;  
   wire [14:0] _id_ctrl_decoder_decoded_T_88={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [14:0] _id_ctrl_decoder_decoded_T_92={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[3],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [14:0] _id_ctrl_decoder_decoded_T_98={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [13:0] _id_ctrl_decoder_decoded_T_130={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[14],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [12:0] _id_ctrl_decoder_decoded_T_136={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],_ibuf_io_inst_0_bits_inst_bits[27],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [16:0] _id_ctrl_decoder_decoded_T_138={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[18],id_ctrl_decoder_decoded_invInputs[19],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[25],_ibuf_io_inst_0_bits_inst_bits[28],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [18:0] _id_ctrl_decoder_decoded_T_140={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[18],id_ctrl_decoder_decoded_invInputs[19],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[25],_ibuf_io_inst_0_bits_inst_bits[28],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T={&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_138} ;  
   wire [21:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_8={&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_8,&_id_ctrl_decoder_decoded_T_12,&_id_ctrl_decoder_decoded_T_14,&_id_ctrl_decoder_decoded_T_22,&_id_ctrl_decoder_decoded_T_26,&_id_ctrl_decoder_decoded_T_28,&_id_ctrl_decoder_decoded_T_38,&_id_ctrl_decoder_decoded_T_40,&_id_ctrl_decoder_decoded_T_48,&_id_ctrl_decoder_decoded_T_52,&_id_ctrl_decoder_decoded_T_62,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_74,&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_92,&_id_ctrl_decoder_decoded_T_98,&_id_ctrl_decoder_decoded_T_130,&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_138} ;  
   wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_10={&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_130} ;  
   wire [5:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_19={&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10]},&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_6,&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_140} ;  
   wire [20:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_45={&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_6,&_id_ctrl_decoder_decoded_T_12,&_id_ctrl_decoder_decoded_T_22,&_id_ctrl_decoder_decoded_T_26,&_id_ctrl_decoder_decoded_T_28,&_id_ctrl_decoder_decoded_T_36,&_id_ctrl_decoder_decoded_T_48,&_id_ctrl_decoder_decoded_T_52,&_id_ctrl_decoder_decoded_T_60,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_76,&_id_ctrl_decoder_decoded_T_86,&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_92,&_id_ctrl_decoder_decoded_T_98,&_id_ctrl_decoder_decoded_T_130,&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_138} ;  
   wire [11:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_47={&_id_ctrl_decoder_decoded_T_18,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]},&_id_ctrl_decoder_decoded_T_22,&_id_ctrl_decoder_decoded_T_26,&_id_ctrl_decoder_decoded_T_28,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_86,&_id_ctrl_decoder_decoded_T_98,&_id_ctrl_decoder_decoded_T_130,&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_138} ;  
   reg id_reg_fence ;  
   wire id_mem_busy=~io_dmem_ordered|io_dmem_req_valid_0 ;  
   wire _io_rocc_cmd_valid_T=wb_reg_valid&wb_ctrl_rocc ;  
   wire _dcache_kill_mem_T=mem_reg_valid&mem_ctrl_wxd ;  
   wire _fp_data_hazard_ex_T_1=ex_reg_inst[11:7]==_ibuf_io_inst_0_bits_inst_rs1 ;  
   wire _fp_data_hazard_mem_T_1=mem_reg_inst[11:7]==_ibuf_io_inst_0_bits_inst_rs1 ;  
   wire _fp_data_hazard_ex_T_3=ex_reg_inst[11:7]==_ibuf_io_inst_0_bits_inst_rs2 ;  
   wire _fp_data_hazard_mem_T_3=mem_reg_inst[11:7]==_ibuf_io_inst_0_bits_inst_rs2 ;  
   reg ex_reg_rs_bypass_0 ;  
   reg ex_reg_rs_bypass_1 ;  
   reg [1:0] ex_reg_rs_lsb_0 ;  
   reg [1:0] ex_reg_rs_lsb_1 ;  
   reg [61:0] ex_reg_rs_msb_0 ;  
   reg [61:0] ex_reg_rs_msb_1 ;  
   reg [63:0] casez_tmp ;  
  always @(*)
       begin 
         casez (ex_reg_rs_lsb_0)
          2 'b00:
             casez_tmp =64'h0;
          2 'b01:
             casez_tmp =mem_reg_wdata;
          2 'b10:
             casez_tmp =wb_reg_wdata;
          default :
             casez_tmp =io_dmem_resp_bits_data_word_bypass;
         endcase 
       end
  
   wire [63:0] ex_rs_0=ex_reg_rs_bypass_0 ? casez_tmp:{ex_reg_rs_msb_0,ex_reg_rs_lsb_0} ;  
   reg [63:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (ex_reg_rs_lsb_1)
          2 'b00:
             casez_tmp_0 =64'h0;
          2 'b01:
             casez_tmp_0 =mem_reg_wdata;
          2 'b10:
             casez_tmp_0 =wb_reg_wdata;
          default :
             casez_tmp_0 =io_dmem_resp_bits_data_word_bypass;
         endcase 
       end
  
   wire [63:0] ex_rs_1=ex_reg_rs_bypass_1 ? casez_tmp_0:{ex_reg_rs_msb_1,ex_reg_rs_lsb_1} ;  
   reg [63:0] casez_tmp_1 ;  
   wire [3:0] _ex_op2_T_1=ex_reg_rvc ? 4'h2:4'h4 ;  
   wire _ex_imm_b0_T_4=ex_ctrl_sel_imm==3'h5 ;  
   wire ex_imm_sign=~_ex_imm_b0_T_4&ex_reg_inst[31] ;  
   wire _ex_imm_b4_1_T=ex_ctrl_sel_imm==3'h2 ;  
   wire _ex_imm_b4_1_T_2=ex_ctrl_sel_imm==3'h1 ;  
   wire _ex_imm_b0_T=ex_ctrl_sel_imm==3'h0 ;  
  always @(*)
       begin 
         casez (ex_ctrl_sel_alu2)
          2 'b00:
             casez_tmp_1 =64'h0;
          2 'b01:
             casez_tmp_1 ={{60{_ex_op2_T_1[3]}},_ex_op2_T_1};
          2 'b10:
             casez_tmp_1 =ex_rs_1;
          default :
             casez_tmp_1 ={{33{ex_imm_sign}},_ex_imm_b4_1_T ? ex_reg_inst[30:20]:{11{ex_imm_sign}},ex_ctrl_sel_imm!=3'h2&ex_ctrl_sel_imm!=3'h3 ? {8{ex_imm_sign}}:ex_reg_inst[19:12],~(_ex_imm_b4_1_T|_ex_imm_b0_T_4)&(ex_ctrl_sel_imm==3'h3 ? ex_reg_inst[20]:_ex_imm_b4_1_T_2 ? ex_reg_inst[7]:ex_imm_sign),_ex_imm_b4_1_T|_ex_imm_b0_T_4 ? 6'h0:ex_reg_inst[30:25],_ex_imm_b4_1_T ? 4'h0:_ex_imm_b0_T|_ex_imm_b4_1_T_2 ? ex_reg_inst[11:8]:_ex_imm_b0_T_4 ? ex_reg_inst[19:16]:ex_reg_inst[24:21],_ex_imm_b0_T ? ex_reg_inst[7]:ex_ctrl_sel_imm==3'h4 ? ex_reg_inst[20]:_ex_imm_b0_T_4&ex_reg_inst[15]};
         endcase 
       end
  
   wire div_io_req_valid=ex_reg_valid&ex_ctrl_div ;  
   wire ex_pc_valid=ex_reg_valid|ex_reg_replay|ex_reg_xcpt_interrupt ;  
   wire wb_dcache_miss=wb_ctrl_mem&~io_dmem_resp_valid ;  
   wire _mem_cfi_taken_T=mem_ctrl_branch&mem_br_taken ;  
   wire [3:0] _mem_br_target_T_6=mem_reg_rvc ? 4'h2:4'h4 ;  
   wire [31:0] _mem_br_target_T_8=_mem_cfi_taken_T ? {{20{mem_reg_inst[31]}},mem_reg_inst[7],mem_reg_inst[30:25],mem_reg_inst[11:8],1'h0}:mem_ctrl_jal ? {{12{mem_reg_inst[31]}},mem_reg_inst[19:12],mem_reg_inst[20],mem_reg_inst[30:21],1'h0}:{{28{_mem_br_target_T_6[3]}},_mem_br_target_T_6} ;  
   wire [33:0] _mem_br_target_T_9=mem_reg_pc+{{2{_mem_br_target_T_8[31]}},_mem_br_target_T_8} ;  
   wire [33:0] _mem_npc_T_4=mem_ctrl_jalr ? {mem_reg_wdata[63:33]==31'h0|(&(mem_reg_wdata[63:33])) ? mem_reg_wdata[33]:~(mem_reg_wdata[32]),mem_reg_wdata[32:0]}:_mem_br_target_T_9 ;  
   wire [33:0] mem_npc=_mem_npc_T_4&34'h3FFFFFFFE ;  
   wire mem_cfi_taken=_mem_cfi_taken_T|mem_ctrl_jalr|mem_ctrl_jal ;  
  assign take_pc_mem=mem_reg_valid&~mem_reg_xcpt&mem_cfi_taken; 
   reg [63:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (ex_ctrl_rocc ? 2'h3:ex_reg_mem_size)
          2 'b00:
             casez_tmp_2 ={2{{2{{2{ex_rs_1[7:0]}}}}}};
          2 'b01:
             casez_tmp_2 ={2{{2{ex_rs_1[15:0]}}}};
          2 'b10:
             casez_tmp_2 ={2{ex_rs_1[31:0]}};
          default :
             casez_tmp_2 =ex_rs_1;
         endcase 
       end
  
   wire mem_debug_breakpoint=mem_reg_load&_bpu_io_debug_ld|mem_reg_store&_bpu_io_debug_st ;  
   wire mem_ldst_xcpt=mem_debug_breakpoint|mem_reg_load&_bpu_io_xcpt_ld|mem_reg_store&_bpu_io_xcpt_st ;  
   wire dcache_kill_mem=_dcache_kill_mem_T&io_dmem_replay_next ;  
   wire killm_common=dcache_kill_mem|take_pc_wb|mem_reg_xcpt|~mem_reg_valid ;  
   reg div_io_kill_REG ;  
   wire _GEN=wb_reg_valid&wb_ctrl_mem ;  
   wire _GEN_0=_GEN&io_dmem_s2_xcpt_pf_st ;  
   wire _GEN_1=_GEN&io_dmem_s2_xcpt_pf_ld ;  
   wire _GEN_2=_GEN&io_dmem_s2_xcpt_ae_st ;  
   wire _GEN_3=_GEN&io_dmem_s2_xcpt_ae_ld ;  
   wire _GEN_4=_GEN&io_dmem_s2_xcpt_ma_st ;  
   wire wb_xcpt=wb_reg_xcpt|_GEN_0|_GEN_1|_GEN_2|_GEN_3|_GEN_4|_GEN&io_dmem_s2_xcpt_ma_ld ;  
   wire wb_wxd=wb_reg_valid&wb_ctrl_wxd ;  
   wire wb_set_sboard=wb_ctrl_div|wb_dcache_miss|wb_ctrl_rocc ;  
   wire replay_wb_common=io_dmem_s2_nack|wb_reg_replay ;  
   wire _replay_wb_T=replay_wb_common|_io_rocc_cmd_valid_T ;  
  assign take_pc_wb=_replay_wb_T|wb_xcpt|_csr_io_eret|wb_reg_flush_pipe; 
   wire dmem_resp_valid=io_dmem_resp_valid&io_dmem_resp_bits_has_data ;  
   wire _GEN_5=dmem_resp_valid&io_dmem_resp_bits_replay&~(io_dmem_resp_bits_tag[0]) ;  
  assign div_io_resp_ready=~_GEN_5&~wb_wxd; 
   wire [4:0] ll_waddr=_GEN_5 ? io_dmem_resp_bits_tag[5:1]:_div_io_resp_bits_tag ;  
   wire ll_wen=_GEN_5|div_io_resp_ready&_div_io_resp_valid ;  
   wire wb_valid=wb_reg_valid&~_replay_wb_T&~wb_xcpt ;  
   wire wb_wen=wb_valid&wb_ctrl_wxd ;  
   wire rf_wen=wb_wen|ll_wen ;  
   wire [4:0] rf_waddr=ll_wen ? ll_waddr:wb_reg_inst[11:7] ;  
   wire [63:0] rf_wdata=dmem_resp_valid&~(io_dmem_resp_bits_tag[0]) ? io_dmem_resp_bits_data:ll_wen ? _div_io_resp_bits_data:(|wb_ctrl_csr) ? _csr_io_rw_rdata:wb_reg_wdata ;  
   wire [63:0] id_rs_0=rf_wen&(|rf_waddr)&rf_waddr==_ibuf_io_inst_0_bits_inst_rs1 ? rf_wdata:_rf_ext_R1_data ;  
   wire [63:0] id_rs_1=rf_wen&(|rf_waddr)&rf_waddr==_ibuf_io_inst_0_bits_inst_rs2 ? rf_wdata:_rf_ext_R0_data ;  
   wire _csr_io_htval_htval_valid_imem_T=wb_reg_cause==64'h14 ;  
   wire tval_any_addr=~wb_reg_xcpt|wb_reg_cause==64'h3|wb_reg_cause==64'h1|wb_reg_cause==64'hC|_csr_io_htval_htval_valid_imem_T ;  
   wire _GEN_6=(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_45)&(|_ibuf_io_inst_0_bits_inst_rs1) ;  
   wire _GEN_7=(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_47)&(|_ibuf_io_inst_0_bits_inst_rs2) ;  
   wire _GEN_8=(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_8)&(|_ibuf_io_inst_0_bits_inst_rd) ;  
   reg [31:0] _r ;  
   wire [31:0] r={_r[31:1],1'h0} ;  
   wire [31:0] _id_sboard_hazard_T=r>>_ibuf_io_inst_0_bits_inst_rs1 ;  
   wire [31:0] _id_sboard_hazard_T_7=r>>_ibuf_io_inst_0_bits_inst_rs2 ;  
   wire [31:0] _id_sboard_hazard_T_14=r>>_ibuf_io_inst_0_bits_inst_rd ;  
   wire data_hazard_mem=mem_ctrl_wxd&(_GEN_6&_fp_data_hazard_mem_T_1|_GEN_7&_fp_data_hazard_mem_T_3|_GEN_8&_ibuf_io_inst_0_bits_inst_rd==mem_reg_inst[11:7]) ;  
   reg dcache_blocked_blocked ;  
   reg rocc_blocked ;  
   wire _ctrl_stalld_T_28=ex_reg_valid&ex_ctrl_wxd&(_GEN_6&_fp_data_hazard_ex_T_1|_GEN_7&_fp_data_hazard_ex_T_3|_GEN_8&_ibuf_io_inst_0_bits_inst_rd==ex_reg_inst[11:7])&((|ex_ctrl_csr)|ex_ctrl_jalr|ex_ctrl_mem|ex_ctrl_mul|ex_ctrl_div|ex_ctrl_fp|ex_ctrl_rocc)|mem_reg_valid&data_hazard_mem&((|mem_ctrl_csr)|mem_ctrl_mem&mem_mem_cmd_bh|mem_ctrl_mul|mem_ctrl_div|mem_ctrl_fp|mem_ctrl_rocc)|wb_reg_valid&wb_ctrl_wxd&(_GEN_6&_ibuf_io_inst_0_bits_inst_rs1==wb_reg_inst[11:7]|_GEN_7&_ibuf_io_inst_0_bits_inst_rs2==wb_reg_inst[11:7]|_GEN_8&_ibuf_io_inst_0_bits_inst_rd==wb_reg_inst[11:7])&wb_set_sboard|_GEN_6&_id_sboard_hazard_T[0]&~(ll_wen&ll_waddr==_ibuf_io_inst_0_bits_inst_rs1)|_GEN_7&_id_sboard_hazard_T_7[0]&~(ll_wen&ll_waddr==_ibuf_io_inst_0_bits_inst_rs2)|_GEN_8&_id_sboard_hazard_T_14[0]&~(ll_wen&ll_waddr==_ibuf_io_inst_0_bits_inst_rd)|_csr_io_singleStep&(ex_reg_valid|mem_reg_valid|wb_reg_valid)|(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_19)&dcache_blocked_blocked&~io_dmem_perf_grant|(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_10)&(~(_div_io_req_ready|_div_io_resp_valid&~wb_wxd)|div_io_req_valid)|id_mem_busy&((|_id_ctrl_decoder_decoded_orMatrixOutputs_T)&_ibuf_io_inst_0_bits_inst_bits[25]|(&_id_ctrl_decoder_decoded_T_46)|id_reg_fence&(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_19))|_csr_io_csr_stall|id_reg_pause ;  
   wire ctrl_killd=~_ibuf_io_inst_0_valid|_ibuf_io_inst_0_bits_replay|ibuf_io_kill|_ctrl_stalld_T_28|_csr_io_interrupt ;  
  assign io_dmem_req_valid_0=ex_reg_valid&ex_ctrl_mem; 
   reg [63:0] coreMonitorBundle_rd0val_REG ;  
   reg [63:0] coreMonitorBundle_rd0val_REG_1 ;  
   reg [63:0] coreMonitorBundle_rd1val_REG ;  
   reg [63:0] coreMonitorBundle_rd1val_REG_1 ;  
   wire coreMonitorBundle_wrenx=wb_wen&~wb_set_sboard ;  
   wire _GEN_9=wb_ctrl_rxs1|wb_ctrl_rfs1 ;  
   wire _GEN_10=wb_ctrl_rxs2|wb_ctrl_rfs2 ;  
  always @( posedge clock)
       begin 
         if (~reset&wb_reg_xcpt&_csr_io_htval_htval_valid_imem_T)
            begin 
              if (1)$display("Assertion failed\n    at RocketCore.scala:718 assert(!htval_valid_imem || io.imem.gpa.valid)\n");
              if (1)$display("");
            end 
         if ((1)&_csr_io_trace_valid_0&~reset)
            begin $fwrite(32'h80000001,"C%d: %d [%d] pc=[%x] W[r%d=%x][%d] R[r%d=%x] R[r%d=%x] inst=[%x] DASM(%x)\n",io_hartid,_csr_io_time[31:0],_csr_io_trace_valid_0&~_csr_io_trace_exception_0,{{30{_csr_io_trace_iaddr_0[33]}},_csr_io_trace_iaddr_0},wb_ctrl_wxd|wb_ctrl_wfd ? wb_reg_inst[11:7]:5'h0,coreMonitorBundle_wrenx ? rf_wdata:64'h0,coreMonitorBundle_wrenx,_GEN_9 ? wb_reg_inst[19:15]:5'h0,_GEN_9 ? coreMonitorBundle_rd0val_REG_1:64'h0,_GEN_10 ? wb_reg_inst[24:20]:5'h0,_GEN_10 ? coreMonitorBundle_rd1val_REG_1:64'h0,_csr_io_trace_insn_0,_csr_io_trace_insn_0);
            end 
       end
  
   wire [7:0] _id_ctrl_decoder_decoded_T_32={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[11]} ;  
   wire [14:0] _id_ctrl_decoder_decoded_T_50={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [15:0] _id_ctrl_decoder_decoded_T_54={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[3],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [15:0] _id_ctrl_decoder_decoded_T_94={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[3],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_104={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[14]} ;  
   wire [8:0] _id_ctrl_decoder_decoded_T_108={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[14]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_114={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[14]} ;  
   wire [8:0] _id_ctrl_decoder_decoded_T_118={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[14]} ;  
   wire [13:0] _id_ctrl_decoder_decoded_T_146={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],_ibuf_io_inst_0_bits_inst_bits[27],_ibuf_io_inst_0_bits_inst_bits[28],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_16={&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_138,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],_ibuf_io_inst_0_bits_inst_bits[31]}} ;  
   wire [2:0] _GEN_11={_ibuf_io_inst_0_bits_xcpt1_pf_inst,_ibuf_io_inst_0_bits_xcpt1_gf_inst,_ibuf_io_inst_0_bits_xcpt1_ae_inst} ;  
   wire _GEN_12=_bpu_io_xcpt_if|(|{_ibuf_io_inst_0_bits_xcpt0_pf_inst,_ibuf_io_inst_0_bits_xcpt0_gf_inst,_ibuf_io_inst_0_bits_xcpt0_ae_inst}) ;  
   wire [31:0] inst=_ibuf_io_inst_0_bits_rvc ? {16'h0,_ibuf_io_inst_0_bits_raw[15:0]}:_ibuf_io_inst_0_bits_raw ;  
   wire _mem_reg_store_T_3=ex_ctrl_mem_cmd==5'h7 ;  
   wire _mem_reg_store_T_5=ex_ctrl_mem_cmd==5'h4 ;  
   wire _mem_reg_store_T_6=ex_ctrl_mem_cmd==5'h9 ;  
   wire _mem_reg_store_T_7=ex_ctrl_mem_cmd==5'hA ;  
   wire _mem_reg_store_T_8=ex_ctrl_mem_cmd==5'hB ;  
   wire _mem_reg_store_T_12=ex_ctrl_mem_cmd==5'h8 ;  
   wire _mem_reg_store_T_13=ex_ctrl_mem_cmd==5'hC ;  
   wire _mem_reg_store_T_14=ex_ctrl_mem_cmd==5'hD ;  
   wire _mem_reg_store_T_15=ex_ctrl_mem_cmd==5'hE ;  
   wire _mem_reg_store_T_16=ex_ctrl_mem_cmd==5'hF ;  
   wire [31:0] _GEN_13=r&~(ll_wen ? 32'h1<<ll_waddr:32'h0) ;  
   wire _GEN_14=wb_set_sboard&wb_wen ;  
   wire [8:0] _id_ctrl_decoder_decoded_T_10={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]} ;  
   wire [7:0] _id_ctrl_decoder_decoded_T_56={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11]} ;  
   wire [27:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_53={&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_6,&_id_ctrl_decoder_decoded_T_10,&_id_ctrl_decoder_decoded_T_12,&_id_ctrl_decoder_decoded_T_14,&_id_ctrl_decoder_decoded_T_22,&_id_ctrl_decoder_decoded_T_26,&_id_ctrl_decoder_decoded_T_28,&_id_ctrl_decoder_decoded_T_36,&_id_ctrl_decoder_decoded_T_40,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],id_ctrl_decoder_decoded_invInputs[19],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_48,&_id_ctrl_decoder_decoded_T_52,&_id_ctrl_decoder_decoded_T_56,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_74,&_id_ctrl_decoder_decoded_T_86,&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_92,&_id_ctrl_decoder_decoded_T_98,&_id_ctrl_decoder_decoded_T_130,&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_140,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],_ibuf_io_inst_0_bits_inst_bits[20],id_ctrl_decoder_decoded_invInputs[19],_ibuf_io_inst_0_bits_inst_bits[22],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],_ibuf_io_inst_0_bits_inst_bits[28],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],id_ctrl_decoder_decoded_invInputs[18],_ibuf_io_inst_0_bits_inst_bits[21],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],_ibuf_io_inst_0_bits_inst_bits[28],_ibuf_io_inst_0_bits_inst_bits[29],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],id_ctrl_decoder_decoded_invInputs[18],_ibuf_io_inst_0_bits_inst_bits[21],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],_ibuf_io_inst_0_bits_inst_bits[24],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],_ibuf_io_inst_0_bits_inst_bits[27],_ibuf_io_inst_0_bits_inst_bits[28],_ibuf_io_inst_0_bits_inst_bits[29],_ibuf_io_inst_0_bits_inst_bits[30],id_ctrl_decoder_decoded_invInputs[29]}} ;  
   wire [2:0] id_ctrl_csr={|{&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],id_ctrl_decoder_decoded_invInputs[19],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_62,&_id_ctrl_decoder_decoded_T_74,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],_ibuf_io_inst_0_bits_inst_bits[20],id_ctrl_decoder_decoded_invInputs[19],_ibuf_io_inst_0_bits_inst_bits[22],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],_ibuf_io_inst_0_bits_inst_bits[28],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],id_ctrl_decoder_decoded_invInputs[18],_ibuf_io_inst_0_bits_inst_bits[21],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],id_ctrl_decoder_decoded_invInputs[22],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],_ibuf_io_inst_0_bits_inst_bits[28],_ibuf_io_inst_0_bits_inst_bits[29],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[5],id_ctrl_decoder_decoded_invInputs[6],id_ctrl_decoder_decoded_invInputs[7],id_ctrl_decoder_decoded_invInputs[8],id_ctrl_decoder_decoded_invInputs[9],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[13],id_ctrl_decoder_decoded_invInputs[14],id_ctrl_decoder_decoded_invInputs[15],id_ctrl_decoder_decoded_invInputs[16],id_ctrl_decoder_decoded_invInputs[17],id_ctrl_decoder_decoded_invInputs[18],_ibuf_io_inst_0_bits_inst_bits[21],id_ctrl_decoder_decoded_invInputs[20],id_ctrl_decoder_decoded_invInputs[21],_ibuf_io_inst_0_bits_inst_bits[24],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],_ibuf_io_inst_0_bits_inst_bits[27],_ibuf_io_inst_0_bits_inst_bits[28],_ibuf_io_inst_0_bits_inst_bits[29],_ibuf_io_inst_0_bits_inst_bits[30],id_ctrl_decoder_decoded_invInputs[29]}},&_id_ctrl_decoder_decoded_T_74,&_id_ctrl_decoder_decoded_T_62} ;  
   wire _id_csr_ren_T=id_ctrl_csr==3'h6 ;  
   wire id_csr_en=_id_csr_ren_T|(&id_ctrl_csr)|id_ctrl_csr==3'h5 ;  
   wire id_system_insn=id_ctrl_csr==3'h4 ;  
   wire id_csr_ren=(_id_csr_ren_T|(&id_ctrl_csr))&~(|_ibuf_io_inst_0_bits_inst_rs1) ;  
   wire id_illegal_insn=~(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_53)|(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_10)&~(_csr_io_status_isa[12])|(|_id_ctrl_decoder_decoded_orMatrixOutputs_T)&~(_csr_io_status_isa[0])|_ibuf_io_inst_0_bits_rvc&~(_csr_io_status_isa[2])|id_csr_en&(_csr_io_decode_0_read_illegal|~id_csr_ren&_csr_io_decode_0_write_illegal)|~_ibuf_io_inst_0_bits_rvc&id_system_insn&_csr_io_decode_0_system_illegal ;  
   wire id_virtual_insn=(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_53)&(id_csr_en&~(~id_csr_ren&_csr_io_decode_0_write_illegal)&_csr_io_decode_0_virtual_access_illegal|~_ibuf_io_inst_0_bits_rvc&id_system_insn&_csr_io_decode_0_virtual_system_illegal) ;  
   wire id_xcpt=_csr_io_interrupt|_bpu_io_debug_if|_bpu_io_xcpt_if|_ibuf_io_inst_0_bits_xcpt0_pf_inst|_ibuf_io_inst_0_bits_xcpt0_gf_inst|_ibuf_io_inst_0_bits_xcpt0_ae_inst|_ibuf_io_inst_0_bits_xcpt1_pf_inst|_ibuf_io_inst_0_bits_xcpt1_gf_inst|_ibuf_io_inst_0_bits_xcpt1_ae_inst|id_virtual_insn|id_illegal_insn ;  
   wire _GEN_15=ex_reg_valid&ex_ctrl_wxd ;  
   wire _GEN_16=_dcache_kill_mem_T&~mem_ctrl_mem ;  
   wire id_bypass_src_1_1=_GEN_15&_fp_data_hazard_ex_T_3 ;  
   wire id_bypass_src_1_2=_GEN_16&_fp_data_hazard_mem_T_3 ;  
   wire do_bypass_1=~(|_ibuf_io_inst_0_bits_inst_rs2)|id_bypass_src_1_1|id_bypass_src_1_2|_dcache_kill_mem_T&_fp_data_hazard_mem_T_3 ;  
   wire _GEN_17=(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_47)&~do_bypass_1 ;  
   wire replay_ex=ex_reg_replay|ex_reg_valid&(ex_ctrl_mem&~io_dmem_req_ready|ex_ctrl_div&~_div_io_req_ready|wb_dcache_miss&ex_reg_load_use) ;  
   wire ctrl_killx=ibuf_io_kill|replay_ex|~ex_reg_valid ;  
   wire mem_pc_valid=mem_reg_valid|mem_reg_replay|mem_reg_xcpt_interrupt ;  
   wire _mem_npc_misaligned_T_3=~(_csr_io_status_isa[2])&_mem_npc_T_4[1] ;  
   wire _GEN_18=mem_reg_valid&mem_reg_flush_pipe ;  
   wire _GEN_19=_GEN_18|~ex_pc_valid ;  
   wire _GEN_20=ex_ctrl_jalr&_csr_io_status_debug ;  
   wire _GEN_21=mem_reg_xcpt_interrupt|mem_reg_xcpt ;  
   wire _GEN_22=mem_reg_valid&_mem_npc_misaligned_T_3 ;  
   wire mem_xcpt=_GEN_21|_GEN_22|mem_reg_valid&mem_ldst_xcpt ;  
   wire _ctrl_killm_T=killm_common|mem_xcpt ;  
   wire [15:0] _id_ctrl_decoder_decoded_T_154={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],_ibuf_io_inst_0_bits_inst_bits[30],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [15:0] _id_ctrl_decoder_decoded_T_158={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],_ibuf_io_inst_0_bits_inst_bits[30],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [15:0] _id_ctrl_decoder_decoded_T_160={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[3],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],_ibuf_io_inst_0_bits_inst_bits[30],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [15:0] _id_ctrl_decoder_decoded_T_162={_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],_ibuf_io_inst_0_bits_inst_bits[30],id_ctrl_decoder_decoded_invInputs[29]} ;  
   wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_12={&_id_ctrl_decoder_decoded_T_18,&_id_ctrl_decoder_decoded_T_146,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],_ibuf_io_inst_0_bits_inst_bits[29]}} ;  
   wire [2:0] _id_ctrl_decoder_decoded_orMatrixOutputs_T_14={&_id_ctrl_decoder_decoded_T_138,&_id_ctrl_decoder_decoded_T_146,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],_ibuf_io_inst_0_bits_inst_bits[3],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],_ibuf_io_inst_0_bits_inst_bits[30]}} ;  
   wire id_bypass_src_0_1=_GEN_15&_fp_data_hazard_ex_T_1 ;  
   wire id_bypass_src_0_2=_GEN_16&_fp_data_hazard_mem_T_1 ;  
   wire do_bypass=~(|_ibuf_io_inst_0_bits_inst_rs1)|id_bypass_src_0_1|id_bypass_src_0_2|_dcache_kill_mem_T&_fp_data_hazard_mem_T_1 ;  
   wire _GEN_23=(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_45)&~do_bypass ;  
   wire _GEN_24=id_illegal_insn|id_virtual_insn ;  
   wire [3:0] id_ctrl_alu_fn={|{&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_86,&_id_ctrl_decoder_decoded_T_154,&_id_ctrl_decoder_decoded_T_158,&_id_ctrl_decoder_decoded_T_160,&_id_ctrl_decoder_decoded_T_162},|{&_id_ctrl_decoder_decoded_T_64,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10],_ibuf_io_inst_0_bits_inst_bits[14]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_86,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[3],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_130},|{&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[13]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[13],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[14]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[14]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[14],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_154,&_id_ctrl_decoder_decoded_T_158,&_id_ctrl_decoder_decoded_T_160,&_id_ctrl_decoder_decoded_T_162},|{&_id_ctrl_decoder_decoded_T_48,&_id_ctrl_decoder_decoded_T_52,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11]},&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_92,&_id_ctrl_decoder_decoded_T_98,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],id_ctrl_decoder_decoded_invInputs[2],_ibuf_io_inst_0_bits_inst_bits[5],_ibuf_io_inst_0_bits_inst_bits[6],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[14]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[13],_ibuf_io_inst_0_bits_inst_bits[14]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]},&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],_ibuf_io_inst_0_bits_inst_bits[14],_ibuf_io_inst_0_bits_inst_bits[25],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[28],id_ctrl_decoder_decoded_invInputs[29]}}} ;  
  always @( posedge clock)
       begin 
         id_reg_pause <=~(_csr_io_time[4:0]==5'h0|_csr_io_inhibit_cycle|io_dmem_perf_release|ibuf_io_kill)&(~ctrl_killd&(&_id_ctrl_decoder_decoded_T_10)&_ibuf_io_inst_0_bits_inst_bits[23:20]==4'h0|id_reg_pause);
         imem_might_request_reg <=ex_pc_valid|mem_pc_valid|_csr_io_customCSRs_0_value[1];
         ex_ctrl_fp <=ctrl_killd&ex_ctrl_fp;
         ex_ctrl_rocc <=ctrl_killd&ex_ctrl_rocc;
         if (~ctrl_killd)
            begin 
              ex_ctrl_branch <=|{&_id_ctrl_decoder_decoded_T_32,&_id_ctrl_decoder_decoded_T_86};
              ex_ctrl_jal <=&_id_ctrl_decoder_decoded_T_40;
              ex_ctrl_jalr <=&_id_ctrl_decoder_decoded_T_38;
              ex_ctrl_rxs2 <=|_id_ctrl_decoder_decoded_orMatrixOutputs_T_47;
              ex_ctrl_rxs1 <=|_id_ctrl_decoder_decoded_orMatrixOutputs_T_45;
              ex_ctrl_sel_alu2 <=id_xcpt ? (_GEN_12 ? 2'h0:{1'h0,|_GEN_11}):{|{&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_6,&_id_ctrl_decoder_decoded_T_12,&_id_ctrl_decoder_decoded_T_14,&_id_ctrl_decoder_decoded_T_22,&_id_ctrl_decoder_decoded_T_26,&_id_ctrl_decoder_decoded_T_28,&_id_ctrl_decoder_decoded_T_32,&_id_ctrl_decoder_decoded_T_36,&_id_ctrl_decoder_decoded_T_48,&_id_ctrl_decoder_decoded_T_52,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_92,&_id_ctrl_decoder_decoded_T_98,&_id_ctrl_decoder_decoded_T_104,&_id_ctrl_decoder_decoded_T_114,&_id_ctrl_decoder_decoded_T_130},|{&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_6,&_id_ctrl_decoder_decoded_T_12,&_id_ctrl_decoder_decoded_T_14,&_id_ctrl_decoder_decoded_T_38,&_id_ctrl_decoder_decoded_T_40,&_id_ctrl_decoder_decoded_T_50,&_id_ctrl_decoder_decoded_T_54,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_94,&_id_ctrl_decoder_decoded_T_108,&_id_ctrl_decoder_decoded_T_118}};
              ex_ctrl_sel_alu1 <=id_xcpt ? (_GEN_12|(|_GEN_11) ? 2'h2:2'h1):{|{&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],_ibuf_io_inst_0_bits_inst_bits[2],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],id_ctrl_decoder_decoded_invInputs[3],id_ctrl_decoder_decoded_invInputs[4]},&_id_ctrl_decoder_decoded_T_40},|{&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_6,&_id_ctrl_decoder_decoded_T_12,&_id_ctrl_decoder_decoded_T_22,&_id_ctrl_decoder_decoded_T_26,&_id_ctrl_decoder_decoded_T_28,&_id_ctrl_decoder_decoded_T_36,&_id_ctrl_decoder_decoded_T_48,&_id_ctrl_decoder_decoded_T_52,&_id_ctrl_decoder_decoded_T_60,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_76,&_id_ctrl_decoder_decoded_T_86,&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_92,&_id_ctrl_decoder_decoded_T_98,&_id_ctrl_decoder_decoded_T_130,&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_138}};
              ex_ctrl_sel_imm <={|{&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_8,&_id_ctrl_decoder_decoded_T_12,&_id_ctrl_decoder_decoded_T_38,&_id_ctrl_decoder_decoded_T_50,&_id_ctrl_decoder_decoded_T_54,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_88,&_id_ctrl_decoder_decoded_T_94,&_id_ctrl_decoder_decoded_T_108,&_id_ctrl_decoder_decoded_T_118},|{&_id_ctrl_decoder_decoded_T_14,&_id_ctrl_decoder_decoded_T_40},|{&_id_ctrl_decoder_decoded_T_32,&_id_ctrl_decoder_decoded_T_40,&_id_ctrl_decoder_decoded_T_104,&_id_ctrl_decoder_decoded_T_114}};
              ex_ctrl_alu_dw <=id_xcpt|(|{&_id_ctrl_decoder_decoded_T,&_id_ctrl_decoder_decoded_T_4,&_id_ctrl_decoder_decoded_T_6,&_id_ctrl_decoder_decoded_T_14,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],id_ctrl_decoder_decoded_invInputs[10],id_ctrl_decoder_decoded_invInputs[11],id_ctrl_decoder_decoded_invInputs[12],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_26,&_id_ctrl_decoder_decoded_T_36,&_id_ctrl_decoder_decoded_T_40,&_id_ctrl_decoder_decoded_T_48,&_id_ctrl_decoder_decoded_T_56,&_id_ctrl_decoder_decoded_T_64,&_id_ctrl_decoder_decoded_T_68,&_id_ctrl_decoder_decoded_T_74,&_id_ctrl_decoder_decoded_T_86,&_id_ctrl_decoder_decoded_T_88,&{_ibuf_io_inst_0_bits_inst_bits[0],_ibuf_io_inst_0_bits_inst_bits[1],id_ctrl_decoder_decoded_invInputs[0],id_ctrl_decoder_decoded_invInputs[1],_ibuf_io_inst_0_bits_inst_bits[4],_ibuf_io_inst_0_bits_inst_bits[5],id_ctrl_decoder_decoded_invInputs[4],_ibuf_io_inst_0_bits_inst_bits[12],id_ctrl_decoder_decoded_invInputs[11],_ibuf_io_inst_0_bits_inst_bits[14],id_ctrl_decoder_decoded_invInputs[23],id_ctrl_decoder_decoded_invInputs[24],id_ctrl_decoder_decoded_invInputs[25],id_ctrl_decoder_decoded_invInputs[26],id_ctrl_decoder_decoded_invInputs[27],id_ctrl_decoder_decoded_invInputs[29]},&_id_ctrl_decoder_decoded_T_136,&_id_ctrl_decoder_decoded_T_138});
              ex_ctrl_alu_fn <=id_xcpt ? 4'h0:id_ctrl_alu_fn;
              ex_ctrl_mem <=|_id_ctrl_decoder_decoded_orMatrixOutputs_T_19;
              ex_ctrl_mem_cmd <={1'h0,&_id_ctrl_decoder_decoded_T_68,|_id_ctrl_decoder_decoded_orMatrixOutputs_T_16,|_id_ctrl_decoder_decoded_orMatrixOutputs_T_14,|_id_ctrl_decoder_decoded_orMatrixOutputs_T_12};
              ex_ctrl_div <=|_id_ctrl_decoder_decoded_orMatrixOutputs_T_10;
              ex_ctrl_wxd <=|_id_ctrl_decoder_decoded_orMatrixOutputs_T_8;
              ex_ctrl_csr <=id_system_insn&(|_id_ctrl_decoder_decoded_orMatrixOutputs_T_19) ? 3'h0:id_csr_ren ? 3'h2:id_ctrl_csr;
              ex_ctrl_fence_i <=&_id_ctrl_decoder_decoded_T_46;
              ex_reg_rvc <=id_xcpt&(|_GEN_11)|_ibuf_io_inst_0_bits_rvc;
              ex_reg_flush_pipe <=(&_id_ctrl_decoder_decoded_T_46)|id_system_insn|id_csr_en&~id_csr_ren&_csr_io_decode_0_write_flush;
              ex_reg_load_use <=mem_reg_valid&data_hazard_mem&mem_ctrl_mem;
              ex_reg_mem_size <={&_id_ctrl_decoder_decoded_T_68,|_id_ctrl_decoder_decoded_orMatrixOutputs_T_16,|_id_ctrl_decoder_decoded_orMatrixOutputs_T_14,|_id_ctrl_decoder_decoded_orMatrixOutputs_T_12}==4'h5 ? {|_ibuf_io_inst_0_bits_inst_rs2,|_ibuf_io_inst_0_bits_inst_rs1}:_ibuf_io_inst_0_bits_inst_bits[13:12];
              ex_reg_rs_bypass_0 <=~_GEN_24&do_bypass;
              ex_reg_rs_bypass_1 <=do_bypass_1;
              ex_reg_rs_lsb_0 <=_GEN_24 ? inst[1:0]:_GEN_23 ? id_rs_0[1:0]:(|_ibuf_io_inst_0_bits_inst_rs1) ? (id_bypass_src_0_1 ? 2'h1:{1'h1,~id_bypass_src_0_2}):2'h0;
              ex_reg_rs_lsb_1 <=_GEN_17 ? id_rs_1[1:0]:(|_ibuf_io_inst_0_bits_inst_rs2) ? (id_bypass_src_1_1 ? 2'h1:{1'h1,~id_bypass_src_1_2}):2'h0;
              if (_GEN_24)
                 ex_reg_rs_msb_0 <={32'h0,inst[31:2]};
               else 
                 if (_GEN_23)
                    ex_reg_rs_msb_0 <=id_rs_0[63:2];
            end 
         ex_ctrl_rfs1 <=ctrl_killd&ex_ctrl_rfs1;
         ex_ctrl_rfs2 <=ctrl_killd&ex_ctrl_rfs2;
         ex_ctrl_wfd <=ctrl_killd&ex_ctrl_wfd;
         ex_ctrl_mul <=ctrl_killd&ex_ctrl_mul;
         if (_GEN_19)
            begin 
            end 
          else 
            begin 
              mem_ctrl_fp <=ex_ctrl_fp;
              mem_ctrl_rocc <=ex_ctrl_rocc;
              mem_ctrl_branch <=ex_ctrl_branch;
              mem_ctrl_jal <=ex_ctrl_jal;
              mem_ctrl_jalr <=ex_ctrl_jalr;
              mem_ctrl_rxs2 <=ex_ctrl_rxs2;
              mem_ctrl_rxs1 <=ex_ctrl_rxs1;
              mem_ctrl_mem <=ex_ctrl_mem;
              mem_ctrl_rfs1 <=ex_ctrl_rfs1;
              mem_ctrl_rfs2 <=ex_ctrl_rfs2;
              mem_ctrl_wfd <=ex_ctrl_wfd;
              mem_ctrl_mul <=ex_ctrl_mul;
              mem_ctrl_div <=ex_ctrl_div;
              mem_ctrl_wxd <=ex_ctrl_wxd;
              mem_ctrl_csr <=ex_ctrl_csr;
              mem_ctrl_fence_i <=_GEN_20|ex_ctrl_fence_i;
            end 
         if (mem_pc_valid)
            begin 
              wb_ctrl_rocc <=mem_ctrl_rocc;
              wb_ctrl_rxs2 <=mem_ctrl_rxs2;
              wb_ctrl_rxs1 <=mem_ctrl_rxs1;
              wb_ctrl_mem <=mem_ctrl_mem;
              wb_ctrl_rfs1 <=mem_ctrl_rfs1;
              wb_ctrl_rfs2 <=mem_ctrl_rfs2;
              wb_ctrl_wfd <=mem_ctrl_wfd;
              wb_ctrl_div <=mem_ctrl_div;
              wb_ctrl_wxd <=mem_ctrl_wxd;
              wb_ctrl_csr <=mem_ctrl_csr;
              wb_ctrl_fence_i <=mem_ctrl_fence_i;
              wb_reg_cause <=_GEN_21 ? mem_reg_cause:{60'h0,_GEN_22 ? 4'h0:mem_debug_breakpoint ? 4'hE:4'h3};
              wb_reg_pc <=mem_reg_pc;
              wb_reg_hls_or_dv <=mem_reg_hls_or_dv;
              wb_reg_inst <=mem_reg_inst;
              wb_reg_raw_inst <=mem_reg_raw_inst;
              wb_reg_wdata <=~mem_reg_xcpt&mem_ctrl_fp&mem_ctrl_wxd ? 64'h0:~mem_reg_xcpt&(mem_ctrl_jalr^_mem_npc_misaligned_T_3) ? {{30{_mem_br_target_T_9[33]}},_mem_br_target_T_9}:mem_reg_wdata;
            end 
         ex_reg_xcpt_interrupt <=~ibuf_io_kill&_ibuf_io_inst_0_valid&_csr_io_interrupt;
         ex_reg_valid <=~ctrl_killd;
         ex_reg_xcpt <=~ctrl_killd&id_xcpt;
         if (~ctrl_killd|_csr_io_interrupt|_ibuf_io_inst_0_bits_replay)
            begin 
              ex_reg_cause <=_csr_io_interrupt ? _csr_io_interrupt_cause:{59'h0,_bpu_io_debug_if ? 5'hE:_bpu_io_xcpt_if ? 5'h3:_ibuf_io_inst_0_bits_xcpt0_pf_inst ? 5'hC:_ibuf_io_inst_0_bits_xcpt0_gf_inst ? 5'h14:_ibuf_io_inst_0_bits_xcpt0_ae_inst ? 5'h1:_ibuf_io_inst_0_bits_xcpt1_pf_inst ? 5'hC:_ibuf_io_inst_0_bits_xcpt1_gf_inst ? 5'h14:_ibuf_io_inst_0_bits_xcpt1_ae_inst ? 5'h1:id_virtual_insn ? 5'h16:5'h2};
              ex_reg_pc <=_ibuf_io_pc;
              ex_reg_inst <=_ibuf_io_inst_0_bits_inst_bits;
              ex_reg_raw_inst <=_ibuf_io_inst_0_bits_raw;
            end 
         ex_reg_replay <=~ibuf_io_kill&_ibuf_io_inst_0_valid&_ibuf_io_inst_0_bits_replay;
         mem_reg_xcpt_interrupt <=~ibuf_io_kill&ex_reg_xcpt_interrupt;
         mem_reg_valid <=~ctrl_killx;
         if (_GEN_19)
            begin 
            end 
          else 
            mem_reg_rvc <=ex_reg_rvc;
         mem_reg_xcpt <=~ctrl_killx&(ex_reg_xcpt_interrupt|ex_reg_xcpt);
         mem_reg_replay <=~ibuf_io_kill&replay_ex;
         if (_GEN_19)
            begin 
            end 
          else 
            begin 
              mem_reg_flush_pipe <=_GEN_20|ex_reg_flush_pipe;
              mem_reg_cause <=ex_reg_cause;
              mem_mem_cmd_bh <=_mem_reg_store_T_3|~(ex_reg_mem_size[1]);
              mem_reg_load <=ex_ctrl_mem&(ex_ctrl_mem_cmd==5'h0|ex_ctrl_mem_cmd==5'h10|ex_ctrl_mem_cmd==5'h6|_mem_reg_store_T_3|_mem_reg_store_T_5|_mem_reg_store_T_6|_mem_reg_store_T_7|_mem_reg_store_T_8|_mem_reg_store_T_12|_mem_reg_store_T_13|_mem_reg_store_T_14|_mem_reg_store_T_15|_mem_reg_store_T_16);
              mem_reg_store <=ex_ctrl_mem&(ex_ctrl_mem_cmd==5'h1|ex_ctrl_mem_cmd==5'h11|_mem_reg_store_T_3|_mem_reg_store_T_5|_mem_reg_store_T_6|_mem_reg_store_T_7|_mem_reg_store_T_8|_mem_reg_store_T_12|_mem_reg_store_T_13|_mem_reg_store_T_14|_mem_reg_store_T_15|_mem_reg_store_T_16);
              mem_reg_pc <=ex_reg_pc;
              mem_reg_inst <=ex_reg_inst;
              mem_reg_hls_or_dv <=_csr_io_status_dv;
              mem_reg_raw_inst <=ex_reg_raw_inst;
              mem_reg_wdata <=_alu_io_out;
            end 
         if (_GEN_18|~(ex_pc_valid&ex_ctrl_rxs2&(ex_ctrl_mem|ex_ctrl_rocc)))
            begin 
            end 
          else 
            mem_reg_rs2 <=casez_tmp_2;
         if (_GEN_19)
            begin 
            end 
          else 
            mem_br_taken <=_alu_io_cmp_out;
         wb_reg_valid <=~_ctrl_killm_T;
         wb_reg_xcpt <=mem_xcpt&~take_pc_wb;
         wb_reg_replay <=(dcache_kill_mem|mem_reg_replay)&~take_pc_wb;
         wb_reg_flush_pipe <=~_ctrl_killm_T&mem_reg_flush_pipe;
         if (~ctrl_killd&_GEN_17)
            ex_reg_rs_msb_1 <=id_rs_1[63:2];
         div_io_kill_REG <=_div_io_req_ready&div_io_req_valid;
         dcache_blocked_blocked <=~io_dmem_req_ready&~io_dmem_perf_grant&(dcache_blocked_blocked|io_dmem_req_valid_0|io_dmem_s2_nack);
         rocc_blocked <=~wb_xcpt&(_io_rocc_cmd_valid_T&~replay_wb_common|rocc_blocked);
         coreMonitorBundle_rd0val_REG <=ex_rs_0;
         coreMonitorBundle_rd0val_REG_1 <=coreMonitorBundle_rd0val_REG;
         coreMonitorBundle_rd1val_REG <=ex_rs_1;
         coreMonitorBundle_rd1val_REG_1 <=coreMonitorBundle_rd1val_REG;
         if (reset)
            begin 
              id_reg_fence <=1'h0;
              _r <=32'h0;
            end 
          else 
            begin 
              id_reg_fence <=~ctrl_killd&((&_id_ctrl_decoder_decoded_T_10)|(|_id_ctrl_decoder_decoded_orMatrixOutputs_T)&_ibuf_io_inst_0_bits_inst_bits[26])|id_mem_busy&id_reg_fence;
              if (ll_wen|_GEN_14)
                 _r <=_GEN_13|(_GEN_14 ? 32'h1<<wb_reg_inst[11:7]:32'h0);
               else 
                 if (ll_wen)
                    _r <=_GEN_13;
            end 
       end
  
  IBuf ibuf(.clock(clock),.reset(reset),.io_imem_ready(io_imem_resp_ready),.io_imem_valid(io_imem_resp_valid),.io_imem_bits_pc(io_imem_resp_bits_pc),.io_imem_bits_data(io_imem_resp_bits_data),.io_imem_bits_xcpt_pf_inst(io_imem_resp_bits_xcpt_pf_inst),.io_imem_bits_xcpt_gf_inst(io_imem_resp_bits_xcpt_gf_inst),.io_imem_bits_xcpt_ae_inst(io_imem_resp_bits_xcpt_ae_inst),.io_imem_bits_replay(io_imem_resp_bits_replay),.io_kill(ibuf_io_kill),.io_pc(_ibuf_io_pc),.io_inst_0_ready(~_ctrl_stalld_T_28),.io_inst_0_valid(_ibuf_io_inst_0_valid),.io_inst_0_bits_xcpt0_pf_inst(_ibuf_io_inst_0_bits_xcpt0_pf_inst),.io_inst_0_bits_xcpt0_gf_inst(_ibuf_io_inst_0_bits_xcpt0_gf_inst),.io_inst_0_bits_xcpt0_ae_inst(_ibuf_io_inst_0_bits_xcpt0_ae_inst),.io_inst_0_bits_xcpt1_pf_inst(_ibuf_io_inst_0_bits_xcpt1_pf_inst),.io_inst_0_bits_xcpt1_gf_inst(_ibuf_io_inst_0_bits_xcpt1_gf_inst),.io_inst_0_bits_xcpt1_ae_inst(_ibuf_io_inst_0_bits_xcpt1_ae_inst),.io_inst_0_bits_replay(_ibuf_io_inst_0_bits_replay),.io_inst_0_bits_rvc(_ibuf_io_inst_0_bits_rvc),.io_inst_0_bits_inst_bits(_ibuf_io_inst_0_bits_inst_bits),.io_inst_0_bits_inst_rd(_ibuf_io_inst_0_bits_inst_rd),.io_inst_0_bits_inst_rs1(_ibuf_io_inst_0_bits_inst_rs1),.io_inst_0_bits_inst_rs2(_ibuf_io_inst_0_bits_inst_rs2),.io_inst_0_bits_raw(_ibuf_io_inst_0_bits_raw)); 
  rf_31x64 rf_ext(.R0_addr(~_ibuf_io_inst_0_bits_inst_rs2),.R0_en(1'h1),.R0_clk(clock),.R0_data(_rf_ext_R0_data),.R1_addr(~_ibuf_io_inst_0_bits_inst_rs1),.R1_en(1'h1),.R1_clk(clock),.R1_data(_rf_ext_R1_data),.W0_addr(~rf_waddr),.W0_en(rf_wen&(|rf_waddr)),.W0_clk(clock),.W0_data(rf_wdata)); 
  CSRFile csr(.clock(clock),.reset(reset),.io_ungated_clock(clock),.io_interrupts_debug(io_interrupts_debug),.io_interrupts_mtip(io_interrupts_mtip),.io_interrupts_msip(io_interrupts_msip),.io_interrupts_meip(io_interrupts_meip),.io_hartid(io_hartid),.io_rw_addr(wb_reg_inst[31:20]),.io_rw_cmd(wb_ctrl_csr&{wb_reg_valid,2'h3}),.io_rw_rdata(_csr_io_rw_rdata),.io_rw_wdata(wb_reg_wdata),.io_decode_0_inst(_ibuf_io_inst_0_bits_inst_bits),.io_decode_0_read_illegal(_csr_io_decode_0_read_illegal),.io_decode_0_write_illegal(_csr_io_decode_0_write_illegal),.io_decode_0_write_flush(_csr_io_decode_0_write_flush),.io_decode_0_system_illegal(_csr_io_decode_0_system_illegal),.io_decode_0_virtual_access_illegal(_csr_io_decode_0_virtual_access_illegal),.io_decode_0_virtual_system_illegal(_csr_io_decode_0_virtual_system_illegal),.io_csr_stall(_csr_io_csr_stall),.io_eret(_csr_io_eret),.io_singleStep(_csr_io_singleStep),.io_status_debug(_csr_io_status_debug),.io_status_wfi(io_wfi),.io_status_isa(_csr_io_status_isa),.io_status_dv(_csr_io_status_dv),.io_status_v(_csr_io_status_v),.io_evec(_csr_io_evec),.io_exception(wb_xcpt),.io_retire(wb_valid),.io_cause(wb_reg_xcpt ? wb_reg_cause:{59'h0,_GEN_0 ? 5'hF:_GEN_1 ? 5'hD:{2'h0,_GEN_2 ? 3'h7:_GEN_3 ? 3'h5:{1'h1,_GEN_4,1'h0}}}),.io_pc(wb_reg_pc),.io_tval(wb_xcpt&(tval_any_addr|wb_reg_cause==64'h2) ? {wb_reg_wdata[63:33]==31'h0|(&(wb_reg_wdata[63:33])) ? wb_reg_wdata[33]:~(wb_reg_wdata[32]),wb_reg_wdata[32:0]}:34'h0),.io_gva(wb_xcpt&(tval_any_addr&_csr_io_status_v|~wb_reg_xcpt&wb_reg_hls_or_dv)),.io_time(_csr_io_time),.io_interrupt(_csr_io_interrupt),.io_interrupt_cause(_csr_io_interrupt_cause),.io_bp_0_control_action(_csr_io_bp_0_control_action),.io_bp_0_control_tmatch(_csr_io_bp_0_control_tmatch),.io_bp_0_control_x(_csr_io_bp_0_control_x),.io_bp_0_control_w(_csr_io_bp_0_control_w),.io_bp_0_control_r(_csr_io_bp_0_control_r),.io_bp_0_address(_csr_io_bp_0_address),.io_pmp_cfg_l_0(io_ptw_pmp_cfg_l_0),.io_pmp_cfg_l_1(io_ptw_pmp_cfg_l_1),.io_pmp_cfg_l_2(io_ptw_pmp_cfg_l_2),.io_pmp_cfg_l_3(io_ptw_pmp_cfg_l_3),.io_pmp_cfg_l_4(io_ptw_pmp_cfg_l_4),.io_pmp_cfg_l_5(io_ptw_pmp_cfg_l_5),.io_pmp_cfg_l_6(io_ptw_pmp_cfg_l_6),.io_pmp_cfg_l_7(io_ptw_pmp_cfg_l_7),.io_pmp_cfg_a_0(io_ptw_pmp_cfg_a_0),.io_pmp_cfg_a_1(io_ptw_pmp_cfg_a_1),.io_pmp_cfg_a_2(io_ptw_pmp_cfg_a_2),.io_pmp_cfg_a_3(io_ptw_pmp_cfg_a_3),.io_pmp_cfg_a_4(io_ptw_pmp_cfg_a_4),.io_pmp_cfg_a_5(io_ptw_pmp_cfg_a_5),.io_pmp_cfg_a_6(io_ptw_pmp_cfg_a_6),.io_pmp_cfg_a_7(io_ptw_pmp_cfg_a_7),.io_pmp_cfg_x_0(io_ptw_pmp_cfg_x_0),.io_pmp_cfg_x_1(io_ptw_pmp_cfg_x_1),.io_pmp_cfg_x_2(io_ptw_pmp_cfg_x_2),.io_pmp_cfg_x_3(io_ptw_pmp_cfg_x_3),.io_pmp_cfg_x_4(io_ptw_pmp_cfg_x_4),.io_pmp_cfg_x_5(io_ptw_pmp_cfg_x_5),.io_pmp_cfg_x_6(io_ptw_pmp_cfg_x_6),.io_pmp_cfg_x_7(io_ptw_pmp_cfg_x_7),.io_pmp_cfg_w_0(io_ptw_pmp_cfg_w_0),.io_pmp_cfg_w_1(io_ptw_pmp_cfg_w_1),.io_pmp_cfg_w_2(io_ptw_pmp_cfg_w_2),.io_pmp_cfg_w_3(io_ptw_pmp_cfg_w_3),.io_pmp_cfg_w_4(io_ptw_pmp_cfg_w_4),.io_pmp_cfg_w_5(io_ptw_pmp_cfg_w_5),.io_pmp_cfg_w_6(io_ptw_pmp_cfg_w_6),.io_pmp_cfg_w_7(io_ptw_pmp_cfg_w_7),.io_pmp_cfg_r_0(io_ptw_pmp_cfg_r_0),.io_pmp_cfg_r_1(io_ptw_pmp_cfg_r_1),.io_pmp_cfg_r_2(io_ptw_pmp_cfg_r_2),.io_pmp_cfg_r_3(io_ptw_pmp_cfg_r_3),.io_pmp_cfg_r_4(io_ptw_pmp_cfg_r_4),.io_pmp_cfg_r_5(io_ptw_pmp_cfg_r_5),.io_pmp_cfg_r_6(io_ptw_pmp_cfg_r_6),.io_pmp_cfg_r_7(io_ptw_pmp_cfg_r_7),.io_pmp_addr_0(io_ptw_pmp_addr_0),.io_pmp_addr_1(io_ptw_pmp_addr_1),.io_pmp_addr_2(io_ptw_pmp_addr_2),.io_pmp_addr_3(io_ptw_pmp_addr_3),.io_pmp_addr_4(io_ptw_pmp_addr_4),.io_pmp_addr_5(io_ptw_pmp_addr_5),.io_pmp_addr_6(io_ptw_pmp_addr_6),.io_pmp_addr_7(io_ptw_pmp_addr_7),.io_pmp_mask_0(io_ptw_pmp_mask_0),.io_pmp_mask_1(io_ptw_pmp_mask_1),.io_pmp_mask_2(io_ptw_pmp_mask_2),.io_pmp_mask_3(io_ptw_pmp_mask_3),.io_pmp_mask_4(io_ptw_pmp_mask_4),.io_pmp_mask_5(io_ptw_pmp_mask_5),.io_pmp_mask_6(io_ptw_pmp_mask_6),.io_pmp_mask_7(io_ptw_pmp_mask_7),.io_inhibit_cycle(_csr_io_inhibit_cycle),.io_inst_0({(&(wb_reg_raw_inst[1:0])) ? wb_reg_inst[31:16]:16'h0,wb_reg_raw_inst[15:0]}),.io_trace_valid_0(_csr_io_trace_valid_0),.io_trace_iaddr_0(_csr_io_trace_iaddr_0),.io_trace_insn_0(_csr_io_trace_insn_0),.io_trace_exception_0(_csr_io_trace_exception_0),.io_customCSRs_0_value(_csr_io_customCSRs_0_value)); 
  BreakpointUnit bpu(.io_status_debug(_csr_io_status_debug),.io_bp_0_control_action(_csr_io_bp_0_control_action),.io_bp_0_control_tmatch(_csr_io_bp_0_control_tmatch),.io_bp_0_control_x(_csr_io_bp_0_control_x),.io_bp_0_control_w(_csr_io_bp_0_control_w),.io_bp_0_control_r(_csr_io_bp_0_control_r),.io_bp_0_address(_csr_io_bp_0_address),.io_pc(_ibuf_io_pc[32:0]),.io_ea(mem_reg_wdata[32:0]),.io_xcpt_if(_bpu_io_xcpt_if),.io_xcpt_ld(_bpu_io_xcpt_ld),.io_xcpt_st(_bpu_io_xcpt_st),.io_debug_if(_bpu_io_debug_if),.io_debug_ld(_bpu_io_debug_ld),.io_debug_st(_bpu_io_debug_st)); 
  ALU alu(.io_dw(ex_ctrl_alu_dw),.io_fn(ex_ctrl_alu_fn),.io_in2(casez_tmp_1),.io_in1(ex_ctrl_sel_alu1==2'h2 ? {{30{ex_reg_pc[33]}},ex_reg_pc}:ex_ctrl_sel_alu1==2'h1 ? ex_rs_0:64'h0),.io_out(_alu_io_out),.io_adder_out(_alu_io_adder_out),.io_cmp_out(_alu_io_cmp_out)); 
  MulDiv div(.clock(clock),.reset(reset),.io_req_ready(_div_io_req_ready),.io_req_valid(div_io_req_valid),.io_req_bits_fn(ex_ctrl_alu_fn),.io_req_bits_dw(ex_ctrl_alu_dw),.io_req_bits_in1(ex_rs_0),.io_req_bits_in2(ex_rs_1),.io_req_bits_tag(ex_reg_inst[11:7]),.io_kill(killm_common&div_io_kill_REG),.io_resp_ready(div_io_resp_ready),.io_resp_valid(_div_io_resp_valid),.io_resp_bits_data(_div_io_resp_bits_data),.io_resp_bits_tag(_div_io_resp_bits_tag)); 
  PlusArgTimeout PlusArgTimeout(.clock(clock),.reset(reset),.io_count(_csr_io_time[31:0])); 
  assign io_imem_might_request=imem_might_request_reg; 
  assign io_imem_req_valid=ibuf_io_kill; 
  assign io_imem_req_bits_pc=wb_xcpt|_csr_io_eret ? _csr_io_evec:_replay_wb_T ? wb_reg_pc:mem_npc; 
  assign io_imem_req_bits_speculative=~take_pc_wb; 
  assign io_imem_btb_update_valid=mem_reg_valid&~take_pc_wb&(ex_pc_valid ? mem_npc!=ex_reg_pc:~(_ibuf_io_inst_0_valid|io_imem_resp_valid)|mem_npc!=_ibuf_io_pc)&(~(mem_ctrl_branch|mem_ctrl_jalr|mem_ctrl_jal)|mem_cfi_taken); 
  assign io_imem_bht_update_valid=mem_reg_valid&~take_pc_wb; 
  assign io_imem_flush_icache=wb_reg_valid&wb_ctrl_fence_i&~io_dmem_s2_nack; 
  assign io_dmem_req_valid=io_dmem_req_valid_0; 
  assign io_dmem_req_bits_addr={ex_rs_0[63:33]==31'h0|(&(ex_rs_0[63:33])) ? _alu_io_adder_out[33]:~(_alu_io_adder_out[32]),_alu_io_adder_out[32:0]}; 
  assign io_dmem_req_bits_tag={ex_reg_inst[11:7],ex_ctrl_fp}; 
  assign io_dmem_req_bits_cmd=ex_ctrl_mem_cmd; 
  assign io_dmem_req_bits_size=ex_reg_mem_size; 
  assign io_dmem_req_bits_signed=~(ex_reg_inst[14]); 
  assign io_dmem_req_bits_dv=_csr_io_status_dv; 
  assign io_dmem_s1_kill=killm_common|mem_ldst_xcpt; 
  assign io_dmem_s1_data_data=mem_reg_rs2; 
  assign io_ptw_status_debug=_csr_io_status_debug; 
  assign io_ptw_customCSRs_csrs_0_value=_csr_io_customCSRs_0_value; 
endmodule
 
module RocketTile (
  input clock,
  input reset,
  input auto_buffer_out_a_ready,
  output auto_buffer_out_a_valid,
  output [2:0] auto_buffer_out_a_bits_opcode,
  output [2:0] auto_buffer_out_a_bits_param,
  output [3:0] auto_buffer_out_a_bits_size,
  output [1:0] auto_buffer_out_a_bits_source,
  output [31:0] auto_buffer_out_a_bits_address,
  output [7:0] auto_buffer_out_a_bits_mask,
  output [63:0] auto_buffer_out_a_bits_data,
  output auto_buffer_out_b_ready,
  input auto_buffer_out_b_valid,
  input [2:0] auto_buffer_out_b_bits_opcode,
  input [1:0] auto_buffer_out_b_bits_param,
  input [3:0] auto_buffer_out_b_bits_size,
  input [1:0] auto_buffer_out_b_bits_source,
  input [31:0] auto_buffer_out_b_bits_address,
  input [7:0] auto_buffer_out_b_bits_mask,
  input auto_buffer_out_b_bits_corrupt,
  input auto_buffer_out_c_ready,
  output auto_buffer_out_c_valid,
  output [2:0] auto_buffer_out_c_bits_opcode,
  output [2:0] auto_buffer_out_c_bits_param,
  output [3:0] auto_buffer_out_c_bits_size,
  output [1:0] auto_buffer_out_c_bits_source,
  output [31:0] auto_buffer_out_c_bits_address,
  output [63:0] auto_buffer_out_c_bits_data,
  output auto_buffer_out_d_ready,
  input auto_buffer_out_d_valid,
  input [2:0] auto_buffer_out_d_bits_opcode,
  input [1:0] auto_buffer_out_d_bits_param,
  input [3:0] auto_buffer_out_d_bits_size,
  input [1:0] auto_buffer_out_d_bits_source,
  input [1:0] auto_buffer_out_d_bits_sink,
  input auto_buffer_out_d_bits_denied,
  input [63:0] auto_buffer_out_d_bits_data,
  input auto_buffer_out_d_bits_corrupt,
  input auto_buffer_out_e_ready,
  output auto_buffer_out_e_valid,
  output [1:0] auto_buffer_out_e_bits_sink,
  output auto_wfi_out_0,
  input auto_int_local_in_2_0,
  input auto_int_local_in_1_0,
  input auto_int_local_in_1_1,
  input auto_int_local_in_0_0,
  input auto_hartid_in) ; 
   wire _core_io_imem_might_request ;  
   wire _core_io_imem_req_valid ;  
   wire [33:0] _core_io_imem_req_bits_pc ;  
   wire _core_io_imem_req_bits_speculative ;  
   wire _core_io_imem_resp_ready ;  
   wire _core_io_imem_btb_update_valid ;  
   wire _core_io_imem_bht_update_valid ;  
   wire _core_io_imem_flush_icache ;  
   wire _core_io_dmem_req_valid ;  
   wire [33:0] _core_io_dmem_req_bits_addr ;  
   wire [5:0] _core_io_dmem_req_bits_tag ;  
   wire [4:0] _core_io_dmem_req_bits_cmd ;  
   wire [1:0] _core_io_dmem_req_bits_size ;  
   wire _core_io_dmem_req_bits_signed ;  
   wire _core_io_dmem_req_bits_dv ;  
   wire _core_io_dmem_s1_kill ;  
   wire [63:0] _core_io_dmem_s1_data_data ;  
   wire _core_io_ptw_status_debug ;  
   wire _core_io_ptw_pmp_cfg_l_0 ;  
   wire _core_io_ptw_pmp_cfg_l_1 ;  
   wire _core_io_ptw_pmp_cfg_l_2 ;  
   wire _core_io_ptw_pmp_cfg_l_3 ;  
   wire _core_io_ptw_pmp_cfg_l_4 ;  
   wire _core_io_ptw_pmp_cfg_l_5 ;  
   wire _core_io_ptw_pmp_cfg_l_6 ;  
   wire _core_io_ptw_pmp_cfg_l_7 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_0 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_1 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_2 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_3 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_4 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_5 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_6 ;  
   wire [1:0] _core_io_ptw_pmp_cfg_a_7 ;  
   wire _core_io_ptw_pmp_cfg_x_0 ;  
   wire _core_io_ptw_pmp_cfg_x_1 ;  
   wire _core_io_ptw_pmp_cfg_x_2 ;  
   wire _core_io_ptw_pmp_cfg_x_3 ;  
   wire _core_io_ptw_pmp_cfg_x_4 ;  
   wire _core_io_ptw_pmp_cfg_x_5 ;  
   wire _core_io_ptw_pmp_cfg_x_6 ;  
   wire _core_io_ptw_pmp_cfg_x_7 ;  
   wire _core_io_ptw_pmp_cfg_w_0 ;  
   wire _core_io_ptw_pmp_cfg_w_1 ;  
   wire _core_io_ptw_pmp_cfg_w_2 ;  
   wire _core_io_ptw_pmp_cfg_w_3 ;  
   wire _core_io_ptw_pmp_cfg_w_4 ;  
   wire _core_io_ptw_pmp_cfg_w_5 ;  
   wire _core_io_ptw_pmp_cfg_w_6 ;  
   wire _core_io_ptw_pmp_cfg_w_7 ;  
   wire _core_io_ptw_pmp_cfg_r_0 ;  
   wire _core_io_ptw_pmp_cfg_r_1 ;  
   wire _core_io_ptw_pmp_cfg_r_2 ;  
   wire _core_io_ptw_pmp_cfg_r_3 ;  
   wire _core_io_ptw_pmp_cfg_r_4 ;  
   wire _core_io_ptw_pmp_cfg_r_5 ;  
   wire _core_io_ptw_pmp_cfg_r_6 ;  
   wire _core_io_ptw_pmp_cfg_r_7 ;  
   wire [29:0] _core_io_ptw_pmp_addr_0 ;  
   wire [29:0] _core_io_ptw_pmp_addr_1 ;  
   wire [29:0] _core_io_ptw_pmp_addr_2 ;  
   wire [29:0] _core_io_ptw_pmp_addr_3 ;  
   wire [29:0] _core_io_ptw_pmp_addr_4 ;  
   wire [29:0] _core_io_ptw_pmp_addr_5 ;  
   wire [29:0] _core_io_ptw_pmp_addr_6 ;  
   wire [29:0] _core_io_ptw_pmp_addr_7 ;  
   wire [31:0] _core_io_ptw_pmp_mask_0 ;  
   wire [31:0] _core_io_ptw_pmp_mask_1 ;  
   wire [31:0] _core_io_ptw_pmp_mask_2 ;  
   wire [31:0] _core_io_ptw_pmp_mask_3 ;  
   wire [31:0] _core_io_ptw_pmp_mask_4 ;  
   wire [31:0] _core_io_ptw_pmp_mask_5 ;  
   wire [31:0] _core_io_ptw_pmp_mask_6 ;  
   wire [31:0] _core_io_ptw_pmp_mask_7 ;  
   wire [63:0] _core_io_ptw_customCSRs_csrs_0_value ;  
   wire _core_io_wfi ;  
   wire _ptw_io_requestor_0_status_debug ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_0 ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_1 ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_2 ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_3 ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_4 ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_5 ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_6 ;  
   wire _ptw_io_requestor_0_pmp_cfg_l_7 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_0 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_1 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_2 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_3 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_4 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_5 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_6 ;  
   wire [1:0] _ptw_io_requestor_0_pmp_cfg_a_7 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_0 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_1 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_2 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_3 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_4 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_5 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_6 ;  
   wire _ptw_io_requestor_0_pmp_cfg_w_7 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_0 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_1 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_2 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_3 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_4 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_5 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_6 ;  
   wire _ptw_io_requestor_0_pmp_cfg_r_7 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_0 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_1 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_2 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_3 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_4 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_5 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_6 ;  
   wire [29:0] _ptw_io_requestor_0_pmp_addr_7 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_0 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_1 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_2 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_3 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_4 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_5 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_6 ;  
   wire [31:0] _ptw_io_requestor_0_pmp_mask_7 ;  
   wire _ptw_io_requestor_1_status_debug ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_0 ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_1 ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_2 ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_3 ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_4 ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_5 ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_6 ;  
   wire _ptw_io_requestor_1_pmp_cfg_l_7 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_0 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_1 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_2 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_3 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_4 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_5 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_6 ;  
   wire [1:0] _ptw_io_requestor_1_pmp_cfg_a_7 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_0 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_1 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_2 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_3 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_4 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_5 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_6 ;  
   wire _ptw_io_requestor_1_pmp_cfg_x_7 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_0 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_1 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_2 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_3 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_4 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_5 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_6 ;  
   wire [29:0] _ptw_io_requestor_1_pmp_addr_7 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_0 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_1 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_2 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_3 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_4 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_5 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_6 ;  
   wire [31:0] _ptw_io_requestor_1_pmp_mask_7 ;  
   wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_0_value ;  
   wire _dcacheArb_io_requestor_0_req_ready ;  
   wire _dcacheArb_io_requestor_0_s2_nack ;  
   wire _dcacheArb_io_requestor_0_resp_valid ;  
   wire [5:0] _dcacheArb_io_requestor_0_resp_bits_tag ;  
   wire [63:0] _dcacheArb_io_requestor_0_resp_bits_data ;  
   wire _dcacheArb_io_requestor_0_resp_bits_replay ;  
   wire _dcacheArb_io_requestor_0_resp_bits_has_data ;  
   wire [63:0] _dcacheArb_io_requestor_0_resp_bits_data_word_bypass ;  
   wire _dcacheArb_io_requestor_0_replay_next ;  
   wire _dcacheArb_io_requestor_0_s2_xcpt_ma_ld ;  
   wire _dcacheArb_io_requestor_0_s2_xcpt_ma_st ;  
   wire _dcacheArb_io_requestor_0_s2_xcpt_pf_ld ;  
   wire _dcacheArb_io_requestor_0_s2_xcpt_pf_st ;  
   wire _dcacheArb_io_requestor_0_s2_xcpt_ae_ld ;  
   wire _dcacheArb_io_requestor_0_s2_xcpt_ae_st ;  
   wire _dcacheArb_io_requestor_0_ordered ;  
   wire _dcacheArb_io_requestor_0_perf_release ;  
   wire _dcacheArb_io_requestor_0_perf_grant ;  
   wire _dcacheArb_io_mem_req_valid ;  
   wire [33:0] _dcacheArb_io_mem_req_bits_addr ;  
   wire [5:0] _dcacheArb_io_mem_req_bits_tag ;  
   wire [4:0] _dcacheArb_io_mem_req_bits_cmd ;  
   wire [1:0] _dcacheArb_io_mem_req_bits_size ;  
   wire _dcacheArb_io_mem_req_bits_signed ;  
   wire _dcacheArb_io_mem_req_bits_dv ;  
   wire _dcacheArb_io_mem_s1_kill ;  
   wire [63:0] _dcacheArb_io_mem_s1_data_data ;  
   wire _frontend_auto_icache_master_out_a_valid ;  
   wire [31:0] _frontend_auto_icache_master_out_a_bits_address ;  
   wire _frontend_io_cpu_resp_valid ;  
   wire [33:0] _frontend_io_cpu_resp_bits_pc ;  
   wire [31:0] _frontend_io_cpu_resp_bits_data ;  
   wire _frontend_io_cpu_resp_bits_xcpt_pf_inst ;  
   wire _frontend_io_cpu_resp_bits_xcpt_gf_inst ;  
   wire _frontend_io_cpu_resp_bits_xcpt_ae_inst ;  
   wire _frontend_io_cpu_resp_bits_replay ;  
   wire _frontend_io_ptw_req_bits_bits_need_gpa ;  
   wire _frontend_io_ptw_req_bits_bits_stage2 ;  
   wire _dcache_auto_out_a_valid ;  
   wire [2:0] _dcache_auto_out_a_bits_opcode ;  
   wire [2:0] _dcache_auto_out_a_bits_param ;  
   wire [3:0] _dcache_auto_out_a_bits_size ;  
   wire _dcache_auto_out_a_bits_source ;  
   wire [31:0] _dcache_auto_out_a_bits_address ;  
   wire [7:0] _dcache_auto_out_a_bits_mask ;  
   wire [63:0] _dcache_auto_out_a_bits_data ;  
   wire _dcache_auto_out_b_ready ;  
   wire _dcache_auto_out_c_valid ;  
   wire [2:0] _dcache_auto_out_c_bits_opcode ;  
   wire [2:0] _dcache_auto_out_c_bits_param ;  
   wire [3:0] _dcache_auto_out_c_bits_size ;  
   wire _dcache_auto_out_c_bits_source ;  
   wire [31:0] _dcache_auto_out_c_bits_address ;  
   wire [63:0] _dcache_auto_out_c_bits_data ;  
   wire _dcache_auto_out_d_ready ;  
   wire _dcache_auto_out_e_valid ;  
   wire [1:0] _dcache_auto_out_e_bits_sink ;  
   wire _dcache_io_cpu_req_ready ;  
   wire _dcache_io_cpu_s2_nack ;  
   wire _dcache_io_cpu_resp_valid ;  
   wire [5:0] _dcache_io_cpu_resp_bits_tag ;  
   wire [63:0] _dcache_io_cpu_resp_bits_data ;  
   wire _dcache_io_cpu_resp_bits_replay ;  
   wire _dcache_io_cpu_resp_bits_has_data ;  
   wire [63:0] _dcache_io_cpu_resp_bits_data_word_bypass ;  
   wire _dcache_io_cpu_replay_next ;  
   wire _dcache_io_cpu_s2_xcpt_ma_ld ;  
   wire _dcache_io_cpu_s2_xcpt_ma_st ;  
   wire _dcache_io_cpu_s2_xcpt_pf_ld ;  
   wire _dcache_io_cpu_s2_xcpt_pf_st ;  
   wire _dcache_io_cpu_s2_xcpt_ae_ld ;  
   wire _dcache_io_cpu_s2_xcpt_ae_st ;  
   wire _dcache_io_cpu_ordered ;  
   wire _dcache_io_cpu_perf_release ;  
   wire _dcache_io_cpu_perf_grant ;  
   wire _dcache_io_ptw_req_bits_bits_need_gpa ;  
   wire _dcache_io_ptw_req_bits_bits_stage2 ;  
   wire _intXbar_auto_int_out_0 ;  
   wire _intXbar_auto_int_out_1 ;  
   wire _intXbar_auto_int_out_2 ;  
   wire _intXbar_auto_int_out_3 ;  
   wire _tlMasterXbar_auto_in_1_a_ready ;  
   wire _tlMasterXbar_auto_in_1_d_valid ;  
   wire [2:0] _tlMasterXbar_auto_in_1_d_bits_opcode ;  
   wire [3:0] _tlMasterXbar_auto_in_1_d_bits_size ;  
   wire [63:0] _tlMasterXbar_auto_in_1_d_bits_data ;  
   wire _tlMasterXbar_auto_in_1_d_bits_corrupt ;  
   wire _tlMasterXbar_auto_in_0_a_ready ;  
   wire _tlMasterXbar_auto_in_0_b_valid ;  
   wire [1:0] _tlMasterXbar_auto_in_0_b_bits_param ;  
   wire [3:0] _tlMasterXbar_auto_in_0_b_bits_size ;  
   wire _tlMasterXbar_auto_in_0_b_bits_source ;  
   wire [31:0] _tlMasterXbar_auto_in_0_b_bits_address ;  
   wire _tlMasterXbar_auto_in_0_c_ready ;  
   wire _tlMasterXbar_auto_in_0_d_valid ;  
   wire [2:0] _tlMasterXbar_auto_in_0_d_bits_opcode ;  
   wire [1:0] _tlMasterXbar_auto_in_0_d_bits_param ;  
   wire [3:0] _tlMasterXbar_auto_in_0_d_bits_size ;  
   wire _tlMasterXbar_auto_in_0_d_bits_source ;  
   wire [1:0] _tlMasterXbar_auto_in_0_d_bits_sink ;  
   wire _tlMasterXbar_auto_in_0_d_bits_denied ;  
   wire [63:0] _tlMasterXbar_auto_in_0_d_bits_data ;  
   wire _tlMasterXbar_auto_in_0_e_ready ;  
   reg wfiNodeOut_0_REG ;  
  always @( posedge clock)
       begin 
         if (reset)
            wfiNodeOut_0_REG <=1'h0;
          else 
            wfiNodeOut_0_REG <=_core_io_wfi;
       end
  
  
wire  tlMasterXbar__clock;
wire  tlMasterXbar__reset;
wire  tlMasterXbar__auto_in_1_a_ready;
wire  tlMasterXbar__auto_in_1_a_valid;
wire [31:0] tlMasterXbar__auto_in_1_a_bits_address;
wire  tlMasterXbar__auto_in_1_d_valid;
wire [2:0] tlMasterXbar__auto_in_1_d_bits_opcode;
wire [3:0] tlMasterXbar__auto_in_1_d_bits_size;
wire [63:0] tlMasterXbar__auto_in_1_d_bits_data;
wire  tlMasterXbar__auto_in_1_d_bits_corrupt;
wire  tlMasterXbar__auto_in_0_a_ready;
wire  tlMasterXbar__auto_in_0_a_valid;
wire [2:0] tlMasterXbar__auto_in_0_a_bits_opcode;
wire [2:0] tlMasterXbar__auto_in_0_a_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_a_bits_size;
wire  tlMasterXbar__auto_in_0_a_bits_source;
wire [31:0] tlMasterXbar__auto_in_0_a_bits_address;
wire [7:0] tlMasterXbar__auto_in_0_a_bits_mask;
wire [63:0] tlMasterXbar__auto_in_0_a_bits_data;
wire  tlMasterXbar__auto_in_0_b_ready;
wire  tlMasterXbar__auto_in_0_b_valid;
wire [1:0] tlMasterXbar__auto_in_0_b_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_b_bits_size;
wire  tlMasterXbar__auto_in_0_b_bits_source;
wire [31:0] tlMasterXbar__auto_in_0_b_bits_address;
wire  tlMasterXbar__auto_in_0_c_ready;
wire  tlMasterXbar__auto_in_0_c_valid;
wire [2:0] tlMasterXbar__auto_in_0_c_bits_opcode;
wire [2:0] tlMasterXbar__auto_in_0_c_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_c_bits_size;
wire  tlMasterXbar__auto_in_0_c_bits_source;
wire [31:0] tlMasterXbar__auto_in_0_c_bits_address;
wire [63:0] tlMasterXbar__auto_in_0_c_bits_data;
wire  tlMasterXbar__auto_in_0_d_ready;
wire  tlMasterXbar__auto_in_0_d_valid;
wire [2:0] tlMasterXbar__auto_in_0_d_bits_opcode;
wire [1:0] tlMasterXbar__auto_in_0_d_bits_param;
wire [3:0] tlMasterXbar__auto_in_0_d_bits_size;
wire  tlMasterXbar__auto_in_0_d_bits_source;
wire [1:0] tlMasterXbar__auto_in_0_d_bits_sink;
wire  tlMasterXbar__auto_in_0_d_bits_denied;
wire [63:0] tlMasterXbar__auto_in_0_d_bits_data;
wire  tlMasterXbar__auto_in_0_e_ready;
wire  tlMasterXbar__auto_in_0_e_valid;
wire [1:0] tlMasterXbar__auto_in_0_e_bits_sink;
wire  tlMasterXbar__auto_out_a_ready;
wire  tlMasterXbar__auto_out_a_valid;
wire [2:0] tlMasterXbar__auto_out_a_bits_opcode;
wire [2:0] tlMasterXbar__auto_out_a_bits_param;
wire [3:0] tlMasterXbar__auto_out_a_bits_size;
wire [1:0] tlMasterXbar__auto_out_a_bits_source;
wire [31:0] tlMasterXbar__auto_out_a_bits_address;
wire [7:0] tlMasterXbar__auto_out_a_bits_mask;
wire [63:0] tlMasterXbar__auto_out_a_bits_data;
wire  tlMasterXbar__auto_out_b_ready;
wire  tlMasterXbar__auto_out_b_valid;
wire [2:0] tlMasterXbar__auto_out_b_bits_opcode;
wire [1:0] tlMasterXbar__auto_out_b_bits_param;
wire [3:0] tlMasterXbar__auto_out_b_bits_size;
wire [1:0] tlMasterXbar__auto_out_b_bits_source;
wire [31:0] tlMasterXbar__auto_out_b_bits_address;
wire [7:0] tlMasterXbar__auto_out_b_bits_mask;
wire  tlMasterXbar__auto_out_b_bits_corrupt;
wire  tlMasterXbar__auto_out_c_ready;
wire  tlMasterXbar__auto_out_c_valid;
wire [2:0] tlMasterXbar__auto_out_c_bits_opcode;
wire [2:0] tlMasterXbar__auto_out_c_bits_param;
wire [3:0] tlMasterXbar__auto_out_c_bits_size;
wire [1:0] tlMasterXbar__auto_out_c_bits_source;
wire [31:0] tlMasterXbar__auto_out_c_bits_address;
wire [63:0] tlMasterXbar__auto_out_c_bits_data;
wire  tlMasterXbar__auto_out_d_ready;
wire  tlMasterXbar__auto_out_d_valid;
wire [2:0] tlMasterXbar__auto_out_d_bits_opcode;
wire [1:0] tlMasterXbar__auto_out_d_bits_param;
wire [3:0] tlMasterXbar__auto_out_d_bits_size;
wire [1:0] tlMasterXbar__auto_out_d_bits_source;
wire [1:0] tlMasterXbar__auto_out_d_bits_sink;
wire  tlMasterXbar__auto_out_d_bits_denied;
wire [63:0] tlMasterXbar__auto_out_d_bits_data;
wire  tlMasterXbar__auto_out_d_bits_corrupt;
wire  tlMasterXbar__auto_out_e_ready;
wire  tlMasterXbar__auto_out_e_valid;
wire [1:0] tlMasterXbar__auto_out_e_bits_sink;
 
   wire  tlMasterXbar__requestDOI_0_1  =  tlMasterXbar__auto_out_d_bits_source  ==2'h2; 
   wire  tlMasterXbar__portsBIO_filtered_valid_0  =  tlMasterXbar__auto_out_b_valid  &~(  tlMasterXbar__auto_out_b_bits_source  [1]); 
   wire  tlMasterXbar__portsDIO_filtered_0_valid  =  tlMasterXbar__auto_out_d_valid  &~(  tlMasterXbar__auto_out_d_bits_source  [1]); 
   wire  tlMasterXbar__portsDIO_filtered_1_valid  =  tlMasterXbar__auto_out_d_valid  &  tlMasterXbar__requestDOI_0_1  ; 
   reg[8:0]  tlMasterXbar__beatsLeft  ; 
   wire  tlMasterXbar__idle  =  tlMasterXbar__beatsLeft  ==9'h0; 
   wire[1:0]  tlMasterXbar__readys_valid  ={  tlMasterXbar__auto_in_1_a_valid  ,  tlMasterXbar__auto_in_0_a_valid  }; 
   reg[1:0]  tlMasterXbar__readys_mask  ; 
   wire[1:0]  tlMasterXbar___readys_filter_T_1  =  tlMasterXbar__readys_valid  &~  tlMasterXbar__readys_mask  ; 
   wire[1:0]  tlMasterXbar__readys_readys  =~({  tlMasterXbar__readys_mask  [1],  tlMasterXbar___readys_filter_T_1  [1]|  tlMasterXbar__readys_mask  [0]}&({  tlMasterXbar___readys_filter_T_1  [0],  tlMasterXbar__auto_in_1_a_valid  }|  tlMasterXbar___readys_filter_T_1  )); 
   wire  tlMasterXbar__winner_0  =  tlMasterXbar__readys_readys  [0]&  tlMasterXbar__auto_in_0_a_valid  ; 
   wire  tlMasterXbar__winner_1  =  tlMasterXbar__readys_readys  [1]&  tlMasterXbar__auto_in_1_a_valid  ; 
   wire  tlMasterXbar___out_0_a_valid_T  =  tlMasterXbar__auto_in_0_a_valid  |  tlMasterXbar__auto_in_1_a_valid  ; 
  always @( posedge   tlMasterXbar__clock  )
       begin 
         if (~  tlMasterXbar__reset  &~(~  tlMasterXbar__winner_0  |~  tlMasterXbar__winner_1  ))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~  tlMasterXbar__reset  &~(~  tlMasterXbar___out_0_a_valid_T  |  tlMasterXbar__winner_0  |  tlMasterXbar__winner_1  ))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg  tlMasterXbar__state_0  ; 
   reg  tlMasterXbar__state_1  ; 
   wire  tlMasterXbar__muxState_0  =  tlMasterXbar__idle   ?   tlMasterXbar__winner_0  :  tlMasterXbar__state_0  ; 
   wire  tlMasterXbar__muxState_1  =  tlMasterXbar__idle   ?   tlMasterXbar__winner_1  :  tlMasterXbar__state_1  ; 
   wire  tlMasterXbar__portsAOI_filtered_0_ready  =  tlMasterXbar__auto_out_a_ready  &(  tlMasterXbar__idle   ?   tlMasterXbar__readys_readys  [0]:  tlMasterXbar__state_0  ); 
   wire  tlMasterXbar__portsAOI_filtered_1_0_ready  =  tlMasterXbar__auto_out_a_ready  &(  tlMasterXbar__idle   ?   tlMasterXbar__readys_readys  [1]:  tlMasterXbar__state_1  ); 
   wire  tlMasterXbar__out_0_a_valid  =  tlMasterXbar__idle   ?   tlMasterXbar___out_0_a_valid_T  :  tlMasterXbar__state_0  &  tlMasterXbar__auto_in_0_a_valid  |  tlMasterXbar__state_1  &  tlMasterXbar__auto_in_1_a_valid  ; 
   wire[26:0]  tlMasterXbar___beatsAI_decode_T_1  =27'hFFF<<  tlMasterXbar__auto_in_0_a_bits_size  ; 
   wire[1:0]  tlMasterXbar___readys_mask_T  =  tlMasterXbar__readys_readys  &  tlMasterXbar__readys_valid  ; 
   wire  tlMasterXbar__latch  =  tlMasterXbar__idle  &  tlMasterXbar__auto_out_a_ready  ; 
  always @( posedge   tlMasterXbar__clock  )
       begin 
         if (  tlMasterXbar__reset  )
            begin  
               tlMasterXbar__beatsLeft   <=9'h0; 
               tlMasterXbar__readys_mask   <=2'h3; 
               tlMasterXbar__state_0   <=1'h0; 
               tlMasterXbar__state_1   <=1'h0;
            end 
          else 
            begin 
              if (  tlMasterXbar__latch  ) 
                  tlMasterXbar__beatsLeft   <=  tlMasterXbar__winner_0  &~(  tlMasterXbar__auto_in_0_a_bits_opcode  [2]) ? ~(  tlMasterXbar___beatsAI_decode_T_1  [11:3]):9'h0;
               else  
                  tlMasterXbar__beatsLeft   <=  tlMasterXbar__beatsLeft  -{8'h0,  tlMasterXbar__auto_out_a_ready  &  tlMasterXbar__out_0_a_valid  };
              if (  tlMasterXbar__latch  &(|  tlMasterXbar__readys_valid  )) 
                  tlMasterXbar__readys_mask   <=  tlMasterXbar___readys_mask_T  |{  tlMasterXbar___readys_mask_T  [0],1'h0};
              if (  tlMasterXbar__idle  )
                 begin  
                    tlMasterXbar__state_0   <=  tlMasterXbar__winner_0  ; 
                    tlMasterXbar__state_1   <=  tlMasterXbar__winner_1  ;
                 end 
            end 
       end
   
  
wire  tlMasterXbar__monitor__clock;
wire  tlMasterXbar__monitor__reset;
wire  tlMasterXbar__monitor__io_in_a_ready;
wire  tlMasterXbar__monitor__io_in_a_valid;
wire [2:0] tlMasterXbar__monitor__io_in_a_bits_opcode;
wire [2:0] tlMasterXbar__monitor__io_in_a_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_a_bits_size;
wire  tlMasterXbar__monitor__io_in_a_bits_source;
wire [31:0] tlMasterXbar__monitor__io_in_a_bits_address;
wire [7:0] tlMasterXbar__monitor__io_in_a_bits_mask;
wire  tlMasterXbar__monitor__io_in_b_ready;
wire  tlMasterXbar__monitor__io_in_b_valid;
wire [2:0] tlMasterXbar__monitor__io_in_b_bits_opcode;
wire [1:0] tlMasterXbar__monitor__io_in_b_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_b_bits_size;
wire  tlMasterXbar__monitor__io_in_b_bits_source;
wire [31:0] tlMasterXbar__monitor__io_in_b_bits_address;
wire [7:0] tlMasterXbar__monitor__io_in_b_bits_mask;
wire  tlMasterXbar__monitor__io_in_b_bits_corrupt;
wire  tlMasterXbar__monitor__io_in_c_ready;
wire  tlMasterXbar__monitor__io_in_c_valid;
wire [2:0] tlMasterXbar__monitor__io_in_c_bits_opcode;
wire [2:0] tlMasterXbar__monitor__io_in_c_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_c_bits_size;
wire  tlMasterXbar__monitor__io_in_c_bits_source;
wire [31:0] tlMasterXbar__monitor__io_in_c_bits_address;
wire  tlMasterXbar__monitor__io_in_d_ready;
wire  tlMasterXbar__monitor__io_in_d_valid;
wire [2:0] tlMasterXbar__monitor__io_in_d_bits_opcode;
wire [1:0] tlMasterXbar__monitor__io_in_d_bits_param;
wire [3:0] tlMasterXbar__monitor__io_in_d_bits_size;
wire  tlMasterXbar__monitor__io_in_d_bits_source;
wire [1:0] tlMasterXbar__monitor__io_in_d_bits_sink;
wire  tlMasterXbar__monitor__io_in_d_bits_denied;
wire  tlMasterXbar__monitor__io_in_d_bits_corrupt;
wire  tlMasterXbar__monitor__io_in_e_ready;
wire  tlMasterXbar__monitor__io_in_e_valid;
wire [1:0] tlMasterXbar__monitor__io_in_e_bits_sink;
 
   wire[31:0]  tlMasterXbar__monitor___plusarg_reader_1_out  ; 
   wire[31:0]  tlMasterXbar__monitor___plusarg_reader_out  ; 
   wire[26:0]  tlMasterXbar__monitor___GEN  ={23'h0,  tlMasterXbar__monitor__io_in_a_bits_size  }; 
   wire[26:0]  tlMasterXbar__monitor___GEN_0  ={23'h0,  tlMasterXbar__monitor__io_in_c_bits_size  }; 
   wire  tlMasterXbar__monitor___a_first_T_1  =  tlMasterXbar__monitor__io_in_a_ready  &  tlMasterXbar__monitor__io_in_a_valid  ; 
   reg[8:0]  tlMasterXbar__monitor__a_first_counter  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode  ; 
   reg[2:0]  tlMasterXbar__monitor__param  ; 
   reg[3:0]  tlMasterXbar__monitor__size  ; 
   reg  tlMasterXbar__monitor__source  ; 
   reg[31:0]  tlMasterXbar__monitor__address  ; 
   wire  tlMasterXbar__monitor___d_first_T_3  =  tlMasterXbar__monitor__io_in_d_ready  &  tlMasterXbar__monitor__io_in_d_valid  ; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode_1  ; 
   reg[1:0]  tlMasterXbar__monitor__param_1  ; 
   reg[3:0]  tlMasterXbar__monitor__size_1  ; 
   reg  tlMasterXbar__monitor__source_1  ; 
   reg[1:0]  tlMasterXbar__monitor__sink  ; 
   reg  tlMasterXbar__monitor__denied  ; 
   reg[8:0]  tlMasterXbar__monitor__b_first_counter  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode_2  ; 
   reg[1:0]  tlMasterXbar__monitor__param_2  ; 
   reg[3:0]  tlMasterXbar__monitor__size_2  ; 
   reg  tlMasterXbar__monitor__source_2  ; 
   reg[31:0]  tlMasterXbar__monitor__address_1  ; 
   wire  tlMasterXbar__monitor___c_first_T_1  =  tlMasterXbar__monitor__io_in_c_ready  &  tlMasterXbar__monitor__io_in_c_valid  ; 
   reg[8:0]  tlMasterXbar__monitor__c_first_counter  ; 
   reg[2:0]  tlMasterXbar__monitor__opcode_3  ; 
   reg[2:0]  tlMasterXbar__monitor__param_3  ; 
   reg[3:0]  tlMasterXbar__monitor__size_3  ; 
   reg  tlMasterXbar__monitor__source_3  ; 
   reg[31:0]  tlMasterXbar__monitor__address_2  ; 
   reg[1:0]  tlMasterXbar__monitor__inflight  ; 
   reg[7:0]  tlMasterXbar__monitor__inflight_opcodes  ; 
   reg[15:0]  tlMasterXbar__monitor__inflight_sizes  ; 
   reg[8:0]  tlMasterXbar__monitor__a_first_counter_1  ; 
   wire  tlMasterXbar__monitor__a_first_1  =  tlMasterXbar__monitor__a_first_counter_1  ==9'h0; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter_1  ; 
   wire  tlMasterXbar__monitor__d_first_1  =  tlMasterXbar__monitor__d_first_counter_1  ==9'h0; 
   wire[7:0]  tlMasterXbar__monitor___a_opcode_lookup_T_1  =  tlMasterXbar__monitor__inflight_opcodes  >>{5'h0,  tlMasterXbar__monitor__io_in_d_bits_source  ,2'h0}; 
   wire[1:0]  tlMasterXbar__monitor___GEN_1  ={1'h0,  tlMasterXbar__monitor__io_in_a_bits_source  }; 
   wire  tlMasterXbar__monitor___GEN_2  =  tlMasterXbar__monitor___a_first_T_1  &  tlMasterXbar__monitor__a_first_1  ; 
   wire  tlMasterXbar__monitor__d_release_ack  =  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h6; 
   wire[1:0]  tlMasterXbar__monitor___GEN_3  ={1'h0,  tlMasterXbar__monitor__io_in_d_bits_source  }; 
   reg[2:0]  tlMasterXbar__monitor__casez_tmp  ; 
  always @(*)
       begin 
         casez (  tlMasterXbar__monitor__io_in_a_bits_opcode  )
          3 'b000: 
              tlMasterXbar__monitor__casez_tmp   =3'h0;
          3 'b001: 
              tlMasterXbar__monitor__casez_tmp   =3'h0;
          3 'b010: 
              tlMasterXbar__monitor__casez_tmp   =3'h1;
          3 'b011: 
              tlMasterXbar__monitor__casez_tmp   =3'h1;
          3 'b100: 
              tlMasterXbar__monitor__casez_tmp   =3'h1;
          3 'b101: 
              tlMasterXbar__monitor__casez_tmp   =3'h2;
          3 'b110: 
              tlMasterXbar__monitor__casez_tmp   =3'h4;
          default : 
              tlMasterXbar__monitor__casez_tmp   =3'h4;
         endcase 
       end
  
   reg[2:0]  tlMasterXbar__monitor__casez_tmp_0  ; 
  always @(*)
       begin 
         casez (  tlMasterXbar__monitor__io_in_a_bits_opcode  )
          3 'b000: 
              tlMasterXbar__monitor__casez_tmp_0   =3'h0;
          3 'b001: 
              tlMasterXbar__monitor__casez_tmp_0   =3'h0;
          3 'b010: 
              tlMasterXbar__monitor__casez_tmp_0   =3'h1;
          3 'b011: 
              tlMasterXbar__monitor__casez_tmp_0   =3'h1;
          3 'b100: 
              tlMasterXbar__monitor__casez_tmp_0   =3'h1;
          3 'b101: 
              tlMasterXbar__monitor__casez_tmp_0   =3'h2;
          3 'b110: 
              tlMasterXbar__monitor__casez_tmp_0   =3'h5;
          default : 
              tlMasterXbar__monitor__casez_tmp_0   =3'h4;
         endcase 
       end
  
   reg[2:0]  tlMasterXbar__monitor__casez_tmp_1  ; 
  always @(*)
       begin 
         casez (  tlMasterXbar__monitor___a_opcode_lookup_T_1  [3:1])
          3 'b000: 
              tlMasterXbar__monitor__casez_tmp_1   =3'h0;
          3 'b001: 
              tlMasterXbar__monitor__casez_tmp_1   =3'h0;
          3 'b010: 
              tlMasterXbar__monitor__casez_tmp_1   =3'h1;
          3 'b011: 
              tlMasterXbar__monitor__casez_tmp_1   =3'h1;
          3 'b100: 
              tlMasterXbar__monitor__casez_tmp_1   =3'h1;
          3 'b101: 
              tlMasterXbar__monitor__casez_tmp_1   =3'h2;
          3 'b110: 
              tlMasterXbar__monitor__casez_tmp_1   =3'h4;
          default : 
              tlMasterXbar__monitor__casez_tmp_1   =3'h4;
         endcase 
       end
  
   reg[2:0]  tlMasterXbar__monitor__casez_tmp_2  ; 
  always @(*)
       begin 
         casez (  tlMasterXbar__monitor___a_opcode_lookup_T_1  [3:1])
          3 'b000: 
              tlMasterXbar__monitor__casez_tmp_2   =3'h0;
          3 'b001: 
              tlMasterXbar__monitor__casez_tmp_2   =3'h0;
          3 'b010: 
              tlMasterXbar__monitor__casez_tmp_2   =3'h1;
          3 'b011: 
              tlMasterXbar__monitor__casez_tmp_2   =3'h1;
          3 'b100: 
              tlMasterXbar__monitor__casez_tmp_2   =3'h1;
          3 'b101: 
              tlMasterXbar__monitor__casez_tmp_2   =3'h2;
          3 'b110: 
              tlMasterXbar__monitor__casez_tmp_2   =3'h5;
          default : 
              tlMasterXbar__monitor__casez_tmp_2   =3'h4;
         endcase 
       end
  
   reg[31:0]  tlMasterXbar__monitor__watchdog  ; 
   reg[1:0]  tlMasterXbar__monitor__inflight_1  ; 
   reg[15:0]  tlMasterXbar__monitor__inflight_sizes_1  ; 
   reg[8:0]  tlMasterXbar__monitor__c_first_counter_1  ; 
   wire  tlMasterXbar__monitor__c_first_1  =  tlMasterXbar__monitor__c_first_counter_1  ==9'h0; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter_2  ; 
   wire  tlMasterXbar__monitor__d_first_2  =  tlMasterXbar__monitor__d_first_counter_2  ==9'h0; 
   wire  tlMasterXbar__monitor___GEN_4  =  tlMasterXbar__monitor__io_in_c_bits_opcode  [2]&  tlMasterXbar__monitor__io_in_c_bits_opcode  [1]; 
   wire[1:0]  tlMasterXbar__monitor___GEN_5  ={1'h0,  tlMasterXbar__monitor__io_in_c_bits_source  }; 
   wire  tlMasterXbar__monitor___GEN_6  =  tlMasterXbar__monitor___c_first_T_1  &  tlMasterXbar__monitor__c_first_1  &  tlMasterXbar__monitor___GEN_4  ; 
   reg[31:0]  tlMasterXbar__monitor__watchdog_1  ; 
   reg[3:0]  tlMasterXbar__monitor__inflight_2  ; 
   reg[8:0]  tlMasterXbar__monitor__d_first_counter_3  ; 
   wire  tlMasterXbar__monitor__d_first_3  =  tlMasterXbar__monitor__d_first_counter_3  ==9'h0; 
   wire  tlMasterXbar__monitor___GEN_7  =  tlMasterXbar__monitor___d_first_T_3  &  tlMasterXbar__monitor__d_first_3  &  tlMasterXbar__monitor__io_in_d_bits_opcode  [2]&~(  tlMasterXbar__monitor__io_in_d_bits_opcode  [1]); 
   wire[3:0]  tlMasterXbar__monitor___GEN_8  ={2'h0,  tlMasterXbar__monitor__io_in_d_bits_sink  }; 
   wire[3:0]  tlMasterXbar__monitor__d_set  =  tlMasterXbar__monitor___GEN_7   ? 4'h1<<  tlMasterXbar__monitor___GEN_8  :4'h0; 
   wire  tlMasterXbar__monitor___GEN_9  =  tlMasterXbar__monitor__io_in_e_ready  &  tlMasterXbar__monitor__io_in_e_valid  ; 
   wire[3:0]  tlMasterXbar__monitor___GEN_10  ={2'h0,  tlMasterXbar__monitor__io_in_e_bits_sink  }; 
   wire[26:0]  tlMasterXbar__monitor___is_aligned_mask_T_1  =27'hFFF<<  tlMasterXbar__monitor___GEN  ; 
   wire[11:0]  tlMasterXbar__monitor___GEN_11  =  tlMasterXbar__monitor__io_in_a_bits_address  [11:0]&~(  tlMasterXbar__monitor___is_aligned_mask_T_1  [11:0]); 
   wire  tlMasterXbar__monitor___mask_T  =  tlMasterXbar__monitor__io_in_a_bits_size  >4'h2; 
   wire  tlMasterXbar__monitor__mask_size  =  tlMasterXbar__monitor__io_in_a_bits_size  [1:0]==2'h2; 
   wire  tlMasterXbar__monitor__mask_acc  =  tlMasterXbar__monitor___mask_T  |  tlMasterXbar__monitor__mask_size  &~(  tlMasterXbar__monitor__io_in_a_bits_address  [2]); 
   wire  tlMasterXbar__monitor__mask_acc_1  =  tlMasterXbar__monitor___mask_T  |  tlMasterXbar__monitor__mask_size  &  tlMasterXbar__monitor__io_in_a_bits_address  [2]; 
   wire  tlMasterXbar__monitor__mask_size_1  =  tlMasterXbar__monitor__io_in_a_bits_size  [1:0]==2'h1; 
   wire  tlMasterXbar__monitor__mask_eq_2  =~(  tlMasterXbar__monitor__io_in_a_bits_address  [2])&~(  tlMasterXbar__monitor__io_in_a_bits_address  [1]); 
   wire  tlMasterXbar__monitor__mask_acc_2  =  tlMasterXbar__monitor__mask_acc  |  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_2  ; 
   wire  tlMasterXbar__monitor__mask_eq_3  =~(  tlMasterXbar__monitor__io_in_a_bits_address  [2])&  tlMasterXbar__monitor__io_in_a_bits_address  [1]; 
   wire  tlMasterXbar__monitor__mask_acc_3  =  tlMasterXbar__monitor__mask_acc  |  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_3  ; 
   wire  tlMasterXbar__monitor__mask_eq_4  =  tlMasterXbar__monitor__io_in_a_bits_address  [2]&~(  tlMasterXbar__monitor__io_in_a_bits_address  [1]); 
   wire  tlMasterXbar__monitor__mask_acc_4  =  tlMasterXbar__monitor__mask_acc_1  |  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_4  ; 
   wire  tlMasterXbar__monitor__mask_eq_5  =  tlMasterXbar__monitor__io_in_a_bits_address  [2]&  tlMasterXbar__monitor__io_in_a_bits_address  [1]; 
   wire  tlMasterXbar__monitor__mask_acc_5  =  tlMasterXbar__monitor__mask_acc_1  |  tlMasterXbar__monitor__mask_size_1  &  tlMasterXbar__monitor__mask_eq_5  ; 
   wire[7:0]  tlMasterXbar__monitor__mask  ={  tlMasterXbar__monitor__mask_acc_5  |  tlMasterXbar__monitor__mask_eq_5  &  tlMasterXbar__monitor__io_in_a_bits_address  [0],  tlMasterXbar__monitor__mask_acc_5  |  tlMasterXbar__monitor__mask_eq_5  &~(  tlMasterXbar__monitor__io_in_a_bits_address  [0]),  tlMasterXbar__monitor__mask_acc_4  |  tlMasterXbar__monitor__mask_eq_4  &  tlMasterXbar__monitor__io_in_a_bits_address  [0],  tlMasterXbar__monitor__mask_acc_4  |  tlMasterXbar__monitor__mask_eq_4  &~(  tlMasterXbar__monitor__io_in_a_bits_address  [0]),  tlMasterXbar__monitor__mask_acc_3  |  tlMasterXbar__monitor__mask_eq_3  &  tlMasterXbar__monitor__io_in_a_bits_address  [0],  tlMasterXbar__monitor__mask_acc_3  |  tlMasterXbar__monitor__mask_eq_3  &~(  tlMasterXbar__monitor__io_in_a_bits_address  [0]),  tlMasterXbar__monitor__mask_acc_2  |  tlMasterXbar__monitor__mask_eq_2  &  tlMasterXbar__monitor__io_in_a_bits_address  [0],  tlMasterXbar__monitor__mask_acc_2  |  tlMasterXbar__monitor__mask_eq_2  &~(  tlMasterXbar__monitor__io_in_a_bits_address  [0])}; 
   wire  tlMasterXbar__monitor___GEN_12  =  tlMasterXbar__monitor__io_in_a_bits_size  <4'hD; 
   wire  tlMasterXbar__monitor___GEN_13  =  tlMasterXbar__monitor__io_in_a_bits_size  <4'h7; 
   wire  tlMasterXbar__monitor___GEN_14  =  tlMasterXbar__monitor__io_in_a_bits_address  [31:28]==4'h8; 
   wire  tlMasterXbar__monitor___GEN_15  =  tlMasterXbar__monitor___GEN_12  &  tlMasterXbar__monitor___GEN_13  &  tlMasterXbar__monitor___GEN_14  ; 
   wire  tlMasterXbar__monitor___GEN_16  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h6&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_17  =  tlMasterXbar__monitor__io_in_a_bits_address  [31:12]==20'h0; 
   wire  tlMasterXbar__monitor___GEN_18  ={  tlMasterXbar__monitor__io_in_a_bits_address  [31:14],~(  tlMasterXbar__monitor__io_in_a_bits_address  [13:12])}==20'h0; 
   wire  tlMasterXbar__monitor___GEN_19  ={  tlMasterXbar__monitor__io_in_a_bits_address  [31:17],~(  tlMasterXbar__monitor__io_in_a_bits_address  [16])}==16'h0; 
   wire  tlMasterXbar__monitor___GEN_20  ={  tlMasterXbar__monitor__io_in_a_bits_address  [31:26],  tlMasterXbar__monitor__io_in_a_bits_address  [25:16]^10'h200}==16'h0; 
   wire  tlMasterXbar__monitor___GEN_21  ={  tlMasterXbar__monitor__io_in_a_bits_address  [31:28],~(  tlMasterXbar__monitor__io_in_a_bits_address  [27:26])}==6'h0; 
   wire  tlMasterXbar__monitor___GEN_22  ={  tlMasterXbar__monitor__io_in_a_bits_address  [31],~(  tlMasterXbar__monitor__io_in_a_bits_address  [30:29])}==3'h0; 
   wire  tlMasterXbar__monitor___GEN_23  =  tlMasterXbar__monitor___GEN_17  |  tlMasterXbar__monitor___GEN_18  ; 
   wire  tlMasterXbar__monitor___GEN_24  =~  tlMasterXbar__monitor__io_in_a_bits_source  &  tlMasterXbar__monitor__io_in_a_bits_size  ==4'h6&  tlMasterXbar__monitor___GEN_12  &(  tlMasterXbar__monitor___GEN_23  |  tlMasterXbar__monitor___GEN_19  |  tlMasterXbar__monitor___GEN_20  |  tlMasterXbar__monitor___GEN_21  |  tlMasterXbar__monitor___GEN_22  |  tlMasterXbar__monitor___GEN_14  ); 
   wire  tlMasterXbar__monitor___GEN_25  =  tlMasterXbar__monitor__io_in_a_bits_param  >3'h2; 
   wire  tlMasterXbar__monitor___GEN_26  =  tlMasterXbar__monitor__io_in_a_bits_mask  !=8'hFF; 
   wire  tlMasterXbar__monitor___GEN_27  =  tlMasterXbar__monitor__io_in_a_valid  &(&  tlMasterXbar__monitor__io_in_a_bits_opcode  )&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_28  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h4&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_29  =  tlMasterXbar__monitor___GEN_12  &  tlMasterXbar__monitor___GEN_18  ; 
   wire  tlMasterXbar__monitor___GEN_30  =  tlMasterXbar__monitor__io_in_a_bits_mask  !=  tlMasterXbar__monitor__mask  ; 
   wire  tlMasterXbar__monitor___GEN_31  =  tlMasterXbar__monitor___GEN_12  &(  tlMasterXbar__monitor___GEN_29  |  tlMasterXbar__monitor___GEN_13  &(  tlMasterXbar__monitor___GEN_17  |  tlMasterXbar__monitor___GEN_20  |  tlMasterXbar__monitor___GEN_21  |  tlMasterXbar__monitor___GEN_14  )|  tlMasterXbar__monitor__io_in_a_bits_size  <4'h9&  tlMasterXbar__monitor___GEN_22  ); 
   wire  tlMasterXbar__monitor___GEN_32  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h0&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_33  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h1&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_34  =  tlMasterXbar__monitor___GEN_12  &  tlMasterXbar__monitor__io_in_a_bits_size  <4'h4&(  tlMasterXbar__monitor___GEN_23  |  tlMasterXbar__monitor___GEN_20  |  tlMasterXbar__monitor___GEN_21  ); 
   wire  tlMasterXbar__monitor___GEN_35  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h2&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_36  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h3&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_37  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_opcode  ==3'h5&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_38  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h6&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_39  =  tlMasterXbar__monitor__io_in_d_bits_size  <4'h3; 
   wire  tlMasterXbar__monitor___GEN_40  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h4&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_41  =  tlMasterXbar__monitor__io_in_d_bits_param  ==2'h2; 
   wire  tlMasterXbar__monitor___GEN_42  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h5&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_43  =~  tlMasterXbar__monitor__io_in_d_bits_denied  |  tlMasterXbar__monitor__io_in_d_bits_corrupt  ; 
   wire  tlMasterXbar__monitor___GEN_44  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h0&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_45  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h1&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_46  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__io_in_d_bits_opcode  ==3'h2&~  tlMasterXbar__monitor__reset  ; 
   wire[19:0]  tlMasterXbar__monitor___GEN_47  ={  tlMasterXbar__monitor__io_in_b_bits_address  [31:14],~(  tlMasterXbar__monitor__io_in_b_bits_address  [13:12])}; 
   wire[5:0]  tlMasterXbar__monitor___GEN_48  ={  tlMasterXbar__monitor__io_in_b_bits_address  [31:28],~(  tlMasterXbar__monitor__io_in_b_bits_address  [27:26])}; 
   wire[15:0]  tlMasterXbar__monitor___GEN_49  ={  tlMasterXbar__monitor__io_in_b_bits_address  [31:26],  tlMasterXbar__monitor__io_in_b_bits_address  [25:16]^10'h200}; 
   wire[15:0]  tlMasterXbar__monitor___GEN_50  ={  tlMasterXbar__monitor__io_in_b_bits_address  [31:17],~(  tlMasterXbar__monitor__io_in_b_bits_address  [16])}; 
   wire  tlMasterXbar__monitor___GEN_51  =  tlMasterXbar__monitor__io_in_b_bits_address  [31:28]!=4'h8; 
   wire[2:0]  tlMasterXbar__monitor___GEN_52  ={  tlMasterXbar__monitor__io_in_b_bits_address  [31],~(  tlMasterXbar__monitor__io_in_b_bits_address  [30:29])}; 
   wire  tlMasterXbar__monitor__address_ok  =~(|  tlMasterXbar__monitor___GEN_47  )|~(|  tlMasterXbar__monitor___GEN_48  )|~(|  tlMasterXbar__monitor___GEN_49  )|~(|(  tlMasterXbar__monitor__io_in_b_bits_address  [31:12]))|~(|  tlMasterXbar__monitor___GEN_50  )|~  tlMasterXbar__monitor___GEN_51  |~(|  tlMasterXbar__monitor___GEN_52  ); 
   wire[26:0]  tlMasterXbar__monitor___is_aligned_mask_T_4  =27'hFFF<<  tlMasterXbar__monitor__io_in_b_bits_size  ; 
   wire[11:0]  tlMasterXbar__monitor___GEN_53  =  tlMasterXbar__monitor__io_in_b_bits_address  [11:0]&~(  tlMasterXbar__monitor___is_aligned_mask_T_4  [11:0]); 
   wire  tlMasterXbar__monitor___mask_T_1  =  tlMasterXbar__monitor__io_in_b_bits_size  >4'h2; 
   wire  tlMasterXbar__monitor__mask_size_3  =  tlMasterXbar__monitor__io_in_b_bits_size  [1:0]==2'h2; 
   wire  tlMasterXbar__monitor__mask_acc_14  =  tlMasterXbar__monitor___mask_T_1  |  tlMasterXbar__monitor__mask_size_3  &~(  tlMasterXbar__monitor__io_in_b_bits_address  [2]); 
   wire  tlMasterXbar__monitor__mask_acc_15  =  tlMasterXbar__monitor___mask_T_1  |  tlMasterXbar__monitor__mask_size_3  &  tlMasterXbar__monitor__io_in_b_bits_address  [2]; 
   wire  tlMasterXbar__monitor__mask_size_4  =  tlMasterXbar__monitor__io_in_b_bits_size  [1:0]==2'h1; 
   wire  tlMasterXbar__monitor__mask_eq_16  =~(  tlMasterXbar__monitor__io_in_b_bits_address  [2])&~(  tlMasterXbar__monitor__io_in_b_bits_address  [1]); 
   wire  tlMasterXbar__monitor__mask_acc_16  =  tlMasterXbar__monitor__mask_acc_14  |  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_16  ; 
   wire  tlMasterXbar__monitor__mask_eq_17  =~(  tlMasterXbar__monitor__io_in_b_bits_address  [2])&  tlMasterXbar__monitor__io_in_b_bits_address  [1]; 
   wire  tlMasterXbar__monitor__mask_acc_17  =  tlMasterXbar__monitor__mask_acc_14  |  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_17  ; 
   wire  tlMasterXbar__monitor__mask_eq_18  =  tlMasterXbar__monitor__io_in_b_bits_address  [2]&~(  tlMasterXbar__monitor__io_in_b_bits_address  [1]); 
   wire  tlMasterXbar__monitor__mask_acc_18  =  tlMasterXbar__monitor__mask_acc_15  |  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_18  ; 
   wire  tlMasterXbar__monitor__mask_eq_19  =  tlMasterXbar__monitor__io_in_b_bits_address  [2]&  tlMasterXbar__monitor__io_in_b_bits_address  [1]; 
   wire  tlMasterXbar__monitor__mask_acc_19  =  tlMasterXbar__monitor__mask_acc_15  |  tlMasterXbar__monitor__mask_size_4  &  tlMasterXbar__monitor__mask_eq_19  ; 
   wire[7:0]  tlMasterXbar__monitor__mask_1  ={  tlMasterXbar__monitor__mask_acc_19  |  tlMasterXbar__monitor__mask_eq_19  &  tlMasterXbar__monitor__io_in_b_bits_address  [0],  tlMasterXbar__monitor__mask_acc_19  |  tlMasterXbar__monitor__mask_eq_19  &~(  tlMasterXbar__monitor__io_in_b_bits_address  [0]),  tlMasterXbar__monitor__mask_acc_18  |  tlMasterXbar__monitor__mask_eq_18  &  tlMasterXbar__monitor__io_in_b_bits_address  [0],  tlMasterXbar__monitor__mask_acc_18  |  tlMasterXbar__monitor__mask_eq_18  &~(  tlMasterXbar__monitor__io_in_b_bits_address  [0]),  tlMasterXbar__monitor__mask_acc_17  |  tlMasterXbar__monitor__mask_eq_17  &  tlMasterXbar__monitor__io_in_b_bits_address  [0],  tlMasterXbar__monitor__mask_acc_17  |  tlMasterXbar__monitor__mask_eq_17  &~(  tlMasterXbar__monitor__io_in_b_bits_address  [0]),  tlMasterXbar__monitor__mask_acc_16  |  tlMasterXbar__monitor__mask_eq_16  &  tlMasterXbar__monitor__io_in_b_bits_address  [0],  tlMasterXbar__monitor__mask_acc_16  |  tlMasterXbar__monitor__mask_eq_16  &~(  tlMasterXbar__monitor__io_in_b_bits_address  [0])}; 
   wire  tlMasterXbar__monitor___GEN_54  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h6&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_55  =  tlMasterXbar__monitor__io_in_b_bits_mask  !=  tlMasterXbar__monitor__mask_1  ; 
   wire  tlMasterXbar__monitor___GEN_56  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h4&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_57  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h0&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_58  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h1&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_59  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h2&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_60  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h3&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_61  =  tlMasterXbar__monitor__io_in_b_valid  &  tlMasterXbar__monitor__io_in_b_bits_opcode  ==3'h5&~  tlMasterXbar__monitor__reset  ; 
   wire[26:0]  tlMasterXbar__monitor___is_aligned_mask_T_7  =27'hFFF<<  tlMasterXbar__monitor___GEN_0  ; 
   wire[11:0]  tlMasterXbar__monitor___GEN_62  =  tlMasterXbar__monitor__io_in_c_bits_address  [11:0]&~(  tlMasterXbar__monitor___is_aligned_mask_T_7  [11:0]); 
   wire[19:0]  tlMasterXbar__monitor___GEN_63  ={  tlMasterXbar__monitor__io_in_c_bits_address  [31:14],~(  tlMasterXbar__monitor__io_in_c_bits_address  [13:12])}; 
   wire[5:0]  tlMasterXbar__monitor___GEN_64  ={  tlMasterXbar__monitor__io_in_c_bits_address  [31:28],~(  tlMasterXbar__monitor__io_in_c_bits_address  [27:26])}; 
   wire[15:0]  tlMasterXbar__monitor___GEN_65  ={  tlMasterXbar__monitor__io_in_c_bits_address  [31:26],  tlMasterXbar__monitor__io_in_c_bits_address  [25:16]^10'h200}; 
   wire[15:0]  tlMasterXbar__monitor___GEN_66  ={  tlMasterXbar__monitor__io_in_c_bits_address  [31:17],~(  tlMasterXbar__monitor__io_in_c_bits_address  [16])}; 
   wire  tlMasterXbar__monitor___GEN_67  =  tlMasterXbar__monitor__io_in_c_bits_address  [31:28]!=4'h8; 
   wire[2:0]  tlMasterXbar__monitor___GEN_68  ={  tlMasterXbar__monitor__io_in_c_bits_address  [31],~(  tlMasterXbar__monitor__io_in_c_bits_address  [30:29])}; 
   wire  tlMasterXbar__monitor__address_ok_1  =~(|  tlMasterXbar__monitor___GEN_63  )|~(|  tlMasterXbar__monitor___GEN_64  )|~(|  tlMasterXbar__monitor___GEN_65  )|~(|(  tlMasterXbar__monitor__io_in_c_bits_address  [31:12]))|~(|  tlMasterXbar__monitor___GEN_66  )|~  tlMasterXbar__monitor___GEN_67  |~(|  tlMasterXbar__monitor___GEN_68  ); 
   wire  tlMasterXbar__monitor___GEN_69  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h4&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_70  =  tlMasterXbar__monitor__io_in_c_bits_size  <4'h3; 
   wire  tlMasterXbar__monitor___GEN_71  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h5&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_72  =  tlMasterXbar__monitor__io_in_c_bits_size  <4'hD; 
   wire  tlMasterXbar__monitor___GEN_73  =  tlMasterXbar__monitor___GEN_72  &  tlMasterXbar__monitor__io_in_c_bits_size  <4'h7&~  tlMasterXbar__monitor___GEN_67  ; 
   wire  tlMasterXbar__monitor___GEN_74  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h6&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_75  =~  tlMasterXbar__monitor__io_in_c_bits_source  &  tlMasterXbar__monitor__io_in_c_bits_size  ==4'h6&  tlMasterXbar__monitor___GEN_72  &(~(|(  tlMasterXbar__monitor__io_in_c_bits_address  [31:12]))|~(|  tlMasterXbar__monitor___GEN_63  )|~(|  tlMasterXbar__monitor___GEN_66  )|~(|  tlMasterXbar__monitor___GEN_65  )|~(|  tlMasterXbar__monitor___GEN_64  )|~(|  tlMasterXbar__monitor___GEN_68  )|~  tlMasterXbar__monitor___GEN_67  ); 
   wire  tlMasterXbar__monitor___GEN_76  =  tlMasterXbar__monitor__io_in_c_valid  &(&  tlMasterXbar__monitor__io_in_c_bits_opcode  )&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_77  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h0&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_78  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h1&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_79  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h2&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_80  =  tlMasterXbar__monitor__io_in_a_valid  &(|  tlMasterXbar__monitor__a_first_counter  )&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_81  =  tlMasterXbar__monitor__io_in_d_valid  &(|  tlMasterXbar__monitor__d_first_counter  )&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_82  =  tlMasterXbar__monitor__io_in_b_valid  &(|  tlMasterXbar__monitor__b_first_counter  )&~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_83  =  tlMasterXbar__monitor__io_in_c_valid  &(|  tlMasterXbar__monitor__c_first_counter  )&~  tlMasterXbar__monitor__reset  ; 
   wire[15:0]  tlMasterXbar__monitor___GEN_84  ={12'h0,  tlMasterXbar__monitor__io_in_d_bits_source  ,3'h0}; 
   wire  tlMasterXbar__monitor___same_cycle_resp_T_1  =  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__a_first_1  ; 
   wire[1:0]  tlMasterXbar__monitor__a_set_wo_ready  =  tlMasterXbar__monitor___same_cycle_resp_T_1   ? 2'h1<<  tlMasterXbar__monitor___GEN_1  :2'h0; 
   wire  tlMasterXbar__monitor___GEN_85  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__d_first_1  ; 
   wire  tlMasterXbar__monitor___GEN_86  =  tlMasterXbar__monitor___GEN_85  &~  tlMasterXbar__monitor__d_release_ack  ; 
   wire  tlMasterXbar__monitor__same_cycle_resp  =  tlMasterXbar__monitor___same_cycle_resp_T_1  &  tlMasterXbar__monitor__io_in_a_bits_source  ==  tlMasterXbar__monitor__io_in_d_bits_source  ; 
   wire  tlMasterXbar__monitor___GEN_87  =  tlMasterXbar__monitor___GEN_86  &  tlMasterXbar__monitor__same_cycle_resp  &~  tlMasterXbar__monitor__reset  ; 
   wire  tlMasterXbar__monitor___GEN_88  =  tlMasterXbar__monitor___GEN_86  &~  tlMasterXbar__monitor__same_cycle_resp  &~  tlMasterXbar__monitor__reset  ; 
   wire[7:0]  tlMasterXbar__monitor___GEN_89  ={4'h0,  tlMasterXbar__monitor__io_in_d_bits_size  }; 
   wire  tlMasterXbar__monitor___same_cycle_resp_T_3  =  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__c_first_1  ; 
   wire[1:0]  tlMasterXbar__monitor__c_set_wo_ready  =  tlMasterXbar__monitor___same_cycle_resp_T_3  &  tlMasterXbar__monitor___GEN_4   ? 2'h1<<  tlMasterXbar__monitor___GEN_5  :2'h0; 
   wire  tlMasterXbar__monitor___GEN_90  =  tlMasterXbar__monitor__io_in_d_valid  &  tlMasterXbar__monitor__d_first_2  ; 
   wire  tlMasterXbar__monitor___GEN_91  =  tlMasterXbar__monitor___GEN_90  &  tlMasterXbar__monitor__d_release_ack  ; 
   wire  tlMasterXbar__monitor__same_cycle_resp_1  =  tlMasterXbar__monitor___same_cycle_resp_T_3  &  tlMasterXbar__monitor__io_in_c_bits_opcode  [2]&  tlMasterXbar__monitor__io_in_c_bits_opcode  [1]&  tlMasterXbar__monitor__io_in_c_bits_source  ==  tlMasterXbar__monitor__io_in_d_bits_source  ; 
   wire[1:0]  tlMasterXbar__monitor___GEN_92  =  tlMasterXbar__monitor__inflight  >>  tlMasterXbar__monitor___GEN_1  ; 
   wire[1:0]  tlMasterXbar__monitor___GEN_93  =  tlMasterXbar__monitor__inflight  >>  tlMasterXbar__monitor___GEN_3  ; 
   wire[15:0]  tlMasterXbar__monitor___a_size_lookup_T_1  =  tlMasterXbar__monitor__inflight_sizes  >>  tlMasterXbar__monitor___GEN_84  ; 
   wire[1:0]  tlMasterXbar__monitor___GEN_94  =  tlMasterXbar__monitor__inflight_1  >>  tlMasterXbar__monitor___GEN_5  ; 
   wire[1:0]  tlMasterXbar__monitor___GEN_95  =  tlMasterXbar__monitor__inflight_1  >>  tlMasterXbar__monitor___GEN_3  ; 
   wire[15:0]  tlMasterXbar__monitor___c_size_lookup_T_1  =  tlMasterXbar__monitor__inflight_sizes_1  >>  tlMasterXbar__monitor___GEN_84  ; 
   wire[3:0]  tlMasterXbar__monitor___GEN_96  =  tlMasterXbar__monitor__inflight_2  >>  tlMasterXbar__monitor___GEN_8  ; 
   wire[3:0]  tlMasterXbar__monitor___GEN_97  =(  tlMasterXbar__monitor__d_set  |  tlMasterXbar__monitor__inflight_2  )>>  tlMasterXbar__monitor___GEN_10  ; 
  always @( posedge   tlMasterXbar__monitor__clock  )
       begin 
         if (  tlMasterXbar__monitor___GEN_16  &~  tlMasterXbar__monitor___GEN_15  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_16  &~  tlMasterXbar__monitor___GEN_24  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_16  &~  tlMasterXbar__monitor___mask_T  )
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_16  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_16  &  tlMasterXbar__monitor___GEN_25  )
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_16  &  tlMasterXbar__monitor___GEN_26  )
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_27  &~  tlMasterXbar__monitor___GEN_15  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_27  &~  tlMasterXbar__monitor___GEN_24  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_27  &~  tlMasterXbar__monitor___mask_T  )
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_27  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_27  &  tlMasterXbar__monitor___GEN_25  )
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_27  &~(|  tlMasterXbar__monitor__io_in_a_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_27  &  tlMasterXbar__monitor___GEN_26  )
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_28  &~  tlMasterXbar__monitor___GEN_12  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_28  &~(  tlMasterXbar__monitor___GEN_29  |  tlMasterXbar__monitor___GEN_13  &(  tlMasterXbar__monitor___GEN_17  |  tlMasterXbar__monitor___GEN_19  |  tlMasterXbar__monitor___GEN_20  |  tlMasterXbar__monitor___GEN_21  |  tlMasterXbar__monitor___GEN_22  |  tlMasterXbar__monitor___GEN_14  )))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_28  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_28  &(|  tlMasterXbar__monitor__io_in_a_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_28  &  tlMasterXbar__monitor___GEN_30  )
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_32  &~  tlMasterXbar__monitor___GEN_31  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_32  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_32  &(|  tlMasterXbar__monitor__io_in_a_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_32  &  tlMasterXbar__monitor___GEN_30  )
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_33  &~  tlMasterXbar__monitor___GEN_31  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_33  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_33  &(|  tlMasterXbar__monitor__io_in_a_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_33  &(|(  tlMasterXbar__monitor__io_in_a_bits_mask  &~  tlMasterXbar__monitor__mask  )))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_35  &~  tlMasterXbar__monitor___GEN_34  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_35  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_35  &  tlMasterXbar__monitor__io_in_a_bits_param  >3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_35  &  tlMasterXbar__monitor___GEN_30  )
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_36  &~  tlMasterXbar__monitor___GEN_34  )
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_36  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_36  &  tlMasterXbar__monitor__io_in_a_bits_param  [2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_36  &  tlMasterXbar__monitor___GEN_30  )
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_37  &~(  tlMasterXbar__monitor___GEN_12  &  tlMasterXbar__monitor___GEN_29  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_37  &(|  tlMasterXbar__monitor___GEN_11  ))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_37  &(|(  tlMasterXbar__monitor__io_in_a_bits_param  [2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_37  &  tlMasterXbar__monitor___GEN_30  )
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor__io_in_d_valid  &~  tlMasterXbar__monitor__reset  &(&  tlMasterXbar__monitor__io_in_d_bits_opcode  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_38  &  tlMasterXbar__monitor___GEN_39  )
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_38  &(|  tlMasterXbar__monitor__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_38  &  tlMasterXbar__monitor__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_38  &  tlMasterXbar__monitor__io_in_d_bits_denied  )
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_40  &  tlMasterXbar__monitor___GEN_39  )
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_40  &(&  tlMasterXbar__monitor__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_40  &  tlMasterXbar__monitor___GEN_41  )
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_40  &  tlMasterXbar__monitor__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_42  &  tlMasterXbar__monitor___GEN_39  )
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_42  &(&  tlMasterXbar__monitor__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_42  &  tlMasterXbar__monitor___GEN_41  )
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_42  &~  tlMasterXbar__monitor___GEN_43  )
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_44  &(|  tlMasterXbar__monitor__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_44  &  tlMasterXbar__monitor__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_45  &(|  tlMasterXbar__monitor__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_45  &~  tlMasterXbar__monitor___GEN_43  )
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_46  &(|  tlMasterXbar__monitor__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_46  &  tlMasterXbar__monitor__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor__io_in_b_valid  &~  tlMasterXbar__monitor__reset  &(&  tlMasterXbar__monitor__io_in_b_bits_opcode  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_54  &~(~  tlMasterXbar__monitor__io_in_b_bits_source  &  tlMasterXbar__monitor__io_in_b_bits_size  ==4'h6&  tlMasterXbar__monitor__io_in_b_bits_size  <4'hD&(~(|(  tlMasterXbar__monitor__io_in_b_bits_address  [31:12]))|~(|  tlMasterXbar__monitor___GEN_47  )|~(|  tlMasterXbar__monitor___GEN_50  )|~(|  tlMasterXbar__monitor___GEN_49  )|~(|  tlMasterXbar__monitor___GEN_48  )|~(|  tlMasterXbar__monitor___GEN_52  )|~  tlMasterXbar__monitor___GEN_51  )))
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_54  &~  tlMasterXbar__monitor__address_ok  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_54  &(|  tlMasterXbar__monitor___GEN_53  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_54  &(&  tlMasterXbar__monitor__io_in_b_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_54  &  tlMasterXbar__monitor___GEN_55  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_54  &  tlMasterXbar__monitor__io_in_b_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_56  )
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_56  &~  tlMasterXbar__monitor__address_ok  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Get carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_56  &(|  tlMasterXbar__monitor___GEN_53  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel Get address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_56  &(|  tlMasterXbar__monitor__io_in_b_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel Get carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_56  &  tlMasterXbar__monitor___GEN_55  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Get contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_56  &  tlMasterXbar__monitor__io_in_b_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Get is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_57  )
            begin 
              if (1)$display("Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_57  &~  tlMasterXbar__monitor__address_ok  )
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_57  &(|  tlMasterXbar__monitor___GEN_53  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_57  &(|  tlMasterXbar__monitor__io_in_b_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_57  &  tlMasterXbar__monitor___GEN_55  )
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_58  )
            begin 
              if (1)$display("Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_58  &~  tlMasterXbar__monitor__address_ok  )
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_58  &(|  tlMasterXbar__monitor___GEN_53  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_58  &(|  tlMasterXbar__monitor__io_in_b_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_58  &(|(  tlMasterXbar__monitor__io_in_b_bits_mask  &~  tlMasterXbar__monitor__mask_1  )))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_59  )
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_59  &~  tlMasterXbar__monitor__address_ok  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_59  &(|  tlMasterXbar__monitor___GEN_53  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_59  &  tlMasterXbar__monitor___GEN_55  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_60  )
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Logical type unsupported by client (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_60  &~  tlMasterXbar__monitor__address_ok  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_60  &(|  tlMasterXbar__monitor___GEN_53  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_60  &  tlMasterXbar__monitor___GEN_55  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_61  )
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Hint type unsupported by client (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_61  &~  tlMasterXbar__monitor__address_ok  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_61  &(|  tlMasterXbar__monitor___GEN_53  ))
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_61  &  tlMasterXbar__monitor___GEN_55  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_61  &  tlMasterXbar__monitor__io_in_b_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_69  &~  tlMasterXbar__monitor__address_ok_1  )
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_69  &  tlMasterXbar__monitor___GEN_70  )
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_69  &(|  tlMasterXbar__monitor___GEN_62  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_69  &(&(  tlMasterXbar__monitor__io_in_c_bits_param  [2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_71  &~  tlMasterXbar__monitor__address_ok_1  )
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_71  &  tlMasterXbar__monitor___GEN_70  )
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_71  &(|  tlMasterXbar__monitor___GEN_62  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_71  &(&(  tlMasterXbar__monitor__io_in_c_bits_param  [2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_74  &~  tlMasterXbar__monitor___GEN_73  )
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_74  &~  tlMasterXbar__monitor___GEN_75  )
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_74  &  tlMasterXbar__monitor___GEN_70  )
            begin 
              if (1)$display("Assertion failed: 'C' channel Release smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_74  &(|  tlMasterXbar__monitor___GEN_62  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_74  &(&(  tlMasterXbar__monitor__io_in_c_bits_param  [2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_76  &~  tlMasterXbar__monitor___GEN_73  )
            begin 
              if (1)$display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_76  &~  tlMasterXbar__monitor___GEN_75  )
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_76  &  tlMasterXbar__monitor___GEN_70  )
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_76  &(|  tlMasterXbar__monitor___GEN_62  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_76  &(&(  tlMasterXbar__monitor__io_in_c_bits_param  [2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_77  &~  tlMasterXbar__monitor__address_ok_1  )
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_77  &(|  tlMasterXbar__monitor___GEN_62  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_77  &(|  tlMasterXbar__monitor__io_in_c_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_78  &~  tlMasterXbar__monitor__address_ok_1  )
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_78  &(|  tlMasterXbar__monitor___GEN_62  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_78  &(|  tlMasterXbar__monitor__io_in_c_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_79  &~  tlMasterXbar__monitor__address_ok_1  )
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_79  &(|  tlMasterXbar__monitor___GEN_62  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_79  &(|  tlMasterXbar__monitor__io_in_c_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_80  &  tlMasterXbar__monitor__io_in_a_bits_opcode  !=  tlMasterXbar__monitor__opcode  )
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_80  &  tlMasterXbar__monitor__io_in_a_bits_param  !=  tlMasterXbar__monitor__param  )
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_80  &  tlMasterXbar__monitor__io_in_a_bits_size  !=  tlMasterXbar__monitor__size  )
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_80  &  tlMasterXbar__monitor__io_in_a_bits_source  !=  tlMasterXbar__monitor__source  )
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_80  &  tlMasterXbar__monitor__io_in_a_bits_address  !=  tlMasterXbar__monitor__address  )
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_81  &  tlMasterXbar__monitor__io_in_d_bits_opcode  !=  tlMasterXbar__monitor__opcode_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_81  &  tlMasterXbar__monitor__io_in_d_bits_param  !=  tlMasterXbar__monitor__param_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_81  &  tlMasterXbar__monitor__io_in_d_bits_size  !=  tlMasterXbar__monitor__size_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_81  &  tlMasterXbar__monitor__io_in_d_bits_source  !=  tlMasterXbar__monitor__source_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_81  &  tlMasterXbar__monitor__io_in_d_bits_sink  !=  tlMasterXbar__monitor__sink  )
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_81  &  tlMasterXbar__monitor__io_in_d_bits_denied  !=  tlMasterXbar__monitor__denied  )
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_82  &  tlMasterXbar__monitor__io_in_b_bits_opcode  !=  tlMasterXbar__monitor__opcode_2  )
            begin 
              if (1)$display("Assertion failed: 'B' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_82  &  tlMasterXbar__monitor__io_in_b_bits_param  !=  tlMasterXbar__monitor__param_2  )
            begin 
              if (1)$display("Assertion failed: 'B' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_82  &  tlMasterXbar__monitor__io_in_b_bits_size  !=  tlMasterXbar__monitor__size_2  )
            begin 
              if (1)$display("Assertion failed: 'B' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_82  &  tlMasterXbar__monitor__io_in_b_bits_source  !=  tlMasterXbar__monitor__source_2  )
            begin 
              if (1)$display("Assertion failed: 'B' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_82  &  tlMasterXbar__monitor__io_in_b_bits_address  !=  tlMasterXbar__monitor__address_1  )
            begin 
              if (1)$display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_83  &  tlMasterXbar__monitor__io_in_c_bits_opcode  !=  tlMasterXbar__monitor__opcode_3  )
            begin 
              if (1)$display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_83  &  tlMasterXbar__monitor__io_in_c_bits_param  !=  tlMasterXbar__monitor__param_3  )
            begin 
              if (1)$display("Assertion failed: 'C' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_83  &  tlMasterXbar__monitor__io_in_c_bits_size  !=  tlMasterXbar__monitor__size_3  )
            begin 
              if (1)$display("Assertion failed: 'C' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_83  &  tlMasterXbar__monitor__io_in_c_bits_source  !=  tlMasterXbar__monitor__source_3  )
            begin 
              if (1)$display("Assertion failed: 'C' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_83  &  tlMasterXbar__monitor__io_in_c_bits_address  !=  tlMasterXbar__monitor__address_2  )
            begin 
              if (1)$display("Assertion failed: 'C' channel address changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_2  &~  tlMasterXbar__monitor__reset  &  tlMasterXbar__monitor___GEN_92  [0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_86  &~  tlMasterXbar__monitor__reset  &~(  tlMasterXbar__monitor___GEN_93  [0]|  tlMasterXbar__monitor__same_cycle_resp  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_87  &~(  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor__casez_tmp  |  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor__casez_tmp_0  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_87  &  tlMasterXbar__monitor__io_in_a_bits_size  !=  tlMasterXbar__monitor__io_in_d_bits_size  )
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_88  &~(  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor__casez_tmp_1  |  tlMasterXbar__monitor__io_in_d_bits_opcode  ==  tlMasterXbar__monitor__casez_tmp_2  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_88  &  tlMasterXbar__monitor___GEN_89  !={1'h0,  tlMasterXbar__monitor___a_size_lookup_T_1  [7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_85  &  tlMasterXbar__monitor__a_first_1  &  tlMasterXbar__monitor__io_in_a_valid  &  tlMasterXbar__monitor__io_in_a_bits_source  ==  tlMasterXbar__monitor__io_in_d_bits_source  &~  tlMasterXbar__monitor__d_release_ack  &~  tlMasterXbar__monitor__reset  &~(~  tlMasterXbar__monitor__io_in_d_ready  |  tlMasterXbar__monitor__io_in_a_ready  ))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~  tlMasterXbar__monitor__reset  &~(  tlMasterXbar__monitor__a_set_wo_ready  !=(  tlMasterXbar__monitor___GEN_86   ? 2'h1<<  tlMasterXbar__monitor___GEN_3  :2'h0)|  tlMasterXbar__monitor__a_set_wo_ready  ==2'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~  tlMasterXbar__monitor__reset  &~(  tlMasterXbar__monitor__inflight  ==2'h0|  tlMasterXbar__monitor___plusarg_reader_out  ==32'h0|  tlMasterXbar__monitor__watchdog  <  tlMasterXbar__monitor___plusarg_reader_out  ))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_6  &~  tlMasterXbar__monitor__reset  &  tlMasterXbar__monitor___GEN_94  [0])
            begin 
              if (1)$display("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_91  &~  tlMasterXbar__monitor__reset  &~(  tlMasterXbar__monitor___GEN_95  [0]|  tlMasterXbar__monitor__same_cycle_resp_1  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_91  &  tlMasterXbar__monitor__same_cycle_resp_1  &~  tlMasterXbar__monitor__reset  &  tlMasterXbar__monitor__io_in_d_bits_size  !=  tlMasterXbar__monitor__io_in_c_bits_size  )
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_91  &~  tlMasterXbar__monitor__same_cycle_resp_1  &~  tlMasterXbar__monitor__reset  &  tlMasterXbar__monitor___GEN_89  !={1'h0,  tlMasterXbar__monitor___c_size_lookup_T_1  [7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_90  &  tlMasterXbar__monitor__c_first_1  &  tlMasterXbar__monitor__io_in_c_valid  &  tlMasterXbar__monitor__io_in_c_bits_source  ==  tlMasterXbar__monitor__io_in_d_bits_source  &  tlMasterXbar__monitor__d_release_ack  &~(  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h4|  tlMasterXbar__monitor__io_in_c_bits_opcode  ==3'h5)&~  tlMasterXbar__monitor__reset  &~(~  tlMasterXbar__monitor__io_in_d_ready  |  tlMasterXbar__monitor__io_in_c_ready  ))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if ((|  tlMasterXbar__monitor__c_set_wo_ready  )&~  tlMasterXbar__monitor__reset  &  tlMasterXbar__monitor__c_set_wo_ready  ==(  tlMasterXbar__monitor___GEN_91   ? 2'h1<<  tlMasterXbar__monitor___GEN_3  :2'h0))
            begin 
              if (1)$display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~  tlMasterXbar__monitor__reset  &~(  tlMasterXbar__monitor__inflight_1  ==2'h0|  tlMasterXbar__monitor___plusarg_reader_1_out  ==32'h0|  tlMasterXbar__monitor__watchdog_1  <  tlMasterXbar__monitor___plusarg_reader_1_out  ))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_7  &~  tlMasterXbar__monitor__reset  &  tlMasterXbar__monitor___GEN_96  [0])
            begin 
              if (1)$display("Assertion failed: 'D' channel re-used a sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor___GEN_9  &~  tlMasterXbar__monitor__reset  &~(  tlMasterXbar__monitor___GEN_97  [0]))
            begin 
              if (1)$display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire[26:0]  tlMasterXbar__monitor___a_first_beats1_decode_T_1  =27'hFFF<<  tlMasterXbar__monitor___GEN  ; 
   wire[26:0]  tlMasterXbar__monitor___a_first_beats1_decode_T_5  =27'hFFF<<  tlMasterXbar__monitor___GEN  ; 
   wire[26:0]  tlMasterXbar__monitor___GEN_98  ={23'h0,  tlMasterXbar__monitor__io_in_d_bits_size  }; 
   wire[26:0]  tlMasterXbar__monitor___d_first_beats1_decode_T_1  =27'hFFF<<  tlMasterXbar__monitor___GEN_98  ; 
   wire[26:0]  tlMasterXbar__monitor___d_first_beats1_decode_T_5  =27'hFFF<<  tlMasterXbar__monitor___GEN_98  ; 
   wire[26:0]  tlMasterXbar__monitor___d_first_beats1_decode_T_9  =27'hFFF<<  tlMasterXbar__monitor___GEN_98  ; 
   wire[26:0]  tlMasterXbar__monitor___d_first_beats1_decode_T_13  =27'hFFF<<  tlMasterXbar__monitor___GEN_98  ; 
   wire[26:0]  tlMasterXbar__monitor___c_first_beats1_decode_T_1  =27'hFFF<<  tlMasterXbar__monitor___GEN_0  ; 
   wire[26:0]  tlMasterXbar__monitor___c_first_beats1_decode_T_5  =27'hFFF<<  tlMasterXbar__monitor___GEN_0  ; 
   wire  tlMasterXbar__monitor___GEN_99  =  tlMasterXbar__monitor___d_first_T_3  &  tlMasterXbar__monitor__d_first_1  &~  tlMasterXbar__monitor__d_release_ack  ; 
   wire[30:0]  tlMasterXbar__monitor___GEN_100  ={27'h0,  tlMasterXbar__monitor__io_in_d_bits_source  ,3'h0}; 
   wire  tlMasterXbar__monitor___GEN_101  =  tlMasterXbar__monitor___d_first_T_3  &  tlMasterXbar__monitor__d_first_2  &  tlMasterXbar__monitor__d_release_ack  ; 
   wire[30:0]  tlMasterXbar__monitor___d_opcodes_clr_T_5  =31'hF<<{28'h0,  tlMasterXbar__monitor__io_in_d_bits_source  ,2'h0}; 
   wire[18:0]  tlMasterXbar__monitor___a_opcodes_set_T_1  ={15'h0,  tlMasterXbar__monitor___GEN_2   ? {  tlMasterXbar__monitor__io_in_a_bits_opcode  ,1'h1}:4'h0}<<{16'h0,  tlMasterXbar__monitor__io_in_a_bits_source  ,2'h0}; 
   wire[30:0]  tlMasterXbar__monitor___d_sizes_clr_T_5  =31'hFF<<  tlMasterXbar__monitor___GEN_100  ; 
   wire[19:0]  tlMasterXbar__monitor___a_sizes_set_T_1  ={15'h0,  tlMasterXbar__monitor___GEN_2   ? {  tlMasterXbar__monitor__io_in_a_bits_size  ,1'h1}:5'h0}<<{16'h0,  tlMasterXbar__monitor__io_in_a_bits_source  ,3'h0}; 
   wire[30:0]  tlMasterXbar__monitor___d_sizes_clr_T_11  =31'hFF<<  tlMasterXbar__monitor___GEN_100  ; 
   wire[19:0]  tlMasterXbar__monitor___c_sizes_set_T_1  ={15'h0,  tlMasterXbar__monitor___GEN_6   ? {  tlMasterXbar__monitor__io_in_c_bits_size  ,1'h1}:5'h0}<<{16'h0,  tlMasterXbar__monitor__io_in_c_bits_source  ,3'h0}; 
   wire  tlMasterXbar__monitor__b_first_done  =  tlMasterXbar__monitor__io_in_b_ready  &  tlMasterXbar__monitor__io_in_b_valid  ; 
  always @( posedge   tlMasterXbar__monitor__clock  )
       begin 
         if (  tlMasterXbar__monitor__reset  )
            begin  
               tlMasterXbar__monitor__a_first_counter   <=9'h0; 
               tlMasterXbar__monitor__d_first_counter   <=9'h0; 
               tlMasterXbar__monitor__b_first_counter   <=9'h0; 
               tlMasterXbar__monitor__c_first_counter   <=9'h0; 
               tlMasterXbar__monitor__inflight   <=2'h0; 
               tlMasterXbar__monitor__inflight_opcodes   <=8'h0; 
               tlMasterXbar__monitor__inflight_sizes   <=16'h0; 
               tlMasterXbar__monitor__a_first_counter_1   <=9'h0; 
               tlMasterXbar__monitor__d_first_counter_1   <=9'h0; 
               tlMasterXbar__monitor__watchdog   <=32'h0; 
               tlMasterXbar__monitor__inflight_1   <=2'h0; 
               tlMasterXbar__monitor__inflight_sizes_1   <=16'h0; 
               tlMasterXbar__monitor__c_first_counter_1   <=9'h0; 
               tlMasterXbar__monitor__d_first_counter_2   <=9'h0; 
               tlMasterXbar__monitor__watchdog_1   <=32'h0; 
               tlMasterXbar__monitor__inflight_2   <=4'h0; 
               tlMasterXbar__monitor__d_first_counter_3   <=9'h0;
            end 
          else 
            begin 
              if (  tlMasterXbar__monitor___a_first_T_1  )
                 begin 
                   if (|  tlMasterXbar__monitor__a_first_counter  ) 
                       tlMasterXbar__monitor__a_first_counter   <=  tlMasterXbar__monitor__a_first_counter  -9'h1;
                    else  
                       tlMasterXbar__monitor__a_first_counter   <=  tlMasterXbar__monitor__io_in_a_bits_opcode  [2] ? 9'h0:~(  tlMasterXbar__monitor___a_first_beats1_decode_T_1  [11:3]);
                   if (  tlMasterXbar__monitor__a_first_1  ) 
                       tlMasterXbar__monitor__a_first_counter_1   <=  tlMasterXbar__monitor__io_in_a_bits_opcode  [2] ? 9'h0:~(  tlMasterXbar__monitor___a_first_beats1_decode_T_5  [11:3]);
                    else  
                       tlMasterXbar__monitor__a_first_counter_1   <=  tlMasterXbar__monitor__a_first_counter_1  -9'h1;
                 end 
              if (  tlMasterXbar__monitor___d_first_T_3  )
                 begin 
                   if (|  tlMasterXbar__monitor__d_first_counter  ) 
                       tlMasterXbar__monitor__d_first_counter   <=  tlMasterXbar__monitor__d_first_counter  -9'h1;
                    else  
                       tlMasterXbar__monitor__d_first_counter   <=  tlMasterXbar__monitor__io_in_d_bits_opcode  [0] ? ~(  tlMasterXbar__monitor___d_first_beats1_decode_T_1  [11:3]):9'h0;
                   if (  tlMasterXbar__monitor__d_first_1  ) 
                       tlMasterXbar__monitor__d_first_counter_1   <=  tlMasterXbar__monitor__io_in_d_bits_opcode  [0] ? ~(  tlMasterXbar__monitor___d_first_beats1_decode_T_5  [11:3]):9'h0;
                    else  
                       tlMasterXbar__monitor__d_first_counter_1   <=  tlMasterXbar__monitor__d_first_counter_1  -9'h1;
                   if (  tlMasterXbar__monitor__d_first_2  ) 
                       tlMasterXbar__monitor__d_first_counter_2   <=  tlMasterXbar__monitor__io_in_d_bits_opcode  [0] ? ~(  tlMasterXbar__monitor___d_first_beats1_decode_T_9  [11:3]):9'h0;
                    else  
                       tlMasterXbar__monitor__d_first_counter_2   <=  tlMasterXbar__monitor__d_first_counter_2  -9'h1;
                   if (  tlMasterXbar__monitor__d_first_3  ) 
                       tlMasterXbar__monitor__d_first_counter_3   <=  tlMasterXbar__monitor__io_in_d_bits_opcode  [0] ? ~(  tlMasterXbar__monitor___d_first_beats1_decode_T_13  [11:3]):9'h0;
                    else  
                       tlMasterXbar__monitor__d_first_counter_3   <=  tlMasterXbar__monitor__d_first_counter_3  -9'h1;
                 end 
              if (  tlMasterXbar__monitor__b_first_done  )
                 begin 
                   if (|  tlMasterXbar__monitor__b_first_counter  ) 
                       tlMasterXbar__monitor__b_first_counter   <=  tlMasterXbar__monitor__b_first_counter  -9'h1;
                    else  
                       tlMasterXbar__monitor__b_first_counter   <=9'h0;
                 end 
              if (  tlMasterXbar__monitor___c_first_T_1  )
                 begin 
                   if (|  tlMasterXbar__monitor__c_first_counter  ) 
                       tlMasterXbar__monitor__c_first_counter   <=  tlMasterXbar__monitor__c_first_counter  -9'h1;
                    else  
                       tlMasterXbar__monitor__c_first_counter   <=  tlMasterXbar__monitor__io_in_c_bits_opcode  [0] ? ~(  tlMasterXbar__monitor___c_first_beats1_decode_T_1  [11:3]):9'h0;
                   if (  tlMasterXbar__monitor__c_first_1  ) 
                       tlMasterXbar__monitor__c_first_counter_1   <=  tlMasterXbar__monitor__io_in_c_bits_opcode  [0] ? ~(  tlMasterXbar__monitor___c_first_beats1_decode_T_5  [11:3]):9'h0;
                    else  
                       tlMasterXbar__monitor__c_first_counter_1   <=  tlMasterXbar__monitor__c_first_counter_1  -9'h1;
                 end  
               tlMasterXbar__monitor__inflight   <=(  tlMasterXbar__monitor__inflight  |(  tlMasterXbar__monitor___GEN_2   ? 2'h1<<  tlMasterXbar__monitor___GEN_1  :2'h0))&~(  tlMasterXbar__monitor___GEN_99   ? 2'h1<<  tlMasterXbar__monitor___GEN_3  :2'h0); 
               tlMasterXbar__monitor__inflight_opcodes   <=(  tlMasterXbar__monitor__inflight_opcodes  |(  tlMasterXbar__monitor___GEN_2   ?   tlMasterXbar__monitor___a_opcodes_set_T_1  [7:0]:8'h0))&~(  tlMasterXbar__monitor___GEN_99   ?   tlMasterXbar__monitor___d_opcodes_clr_T_5  [7:0]:8'h0); 
               tlMasterXbar__monitor__inflight_sizes   <=(  tlMasterXbar__monitor__inflight_sizes  |(  tlMasterXbar__monitor___GEN_2   ?   tlMasterXbar__monitor___a_sizes_set_T_1  [15:0]:16'h0))&~(  tlMasterXbar__monitor___GEN_99   ?   tlMasterXbar__monitor___d_sizes_clr_T_5  [15:0]:16'h0);
              if (  tlMasterXbar__monitor___a_first_T_1  |  tlMasterXbar__monitor___d_first_T_3  ) 
                  tlMasterXbar__monitor__watchdog   <=32'h0;
               else  
                  tlMasterXbar__monitor__watchdog   <=  tlMasterXbar__monitor__watchdog  +32'h1; 
               tlMasterXbar__monitor__inflight_1   <=(  tlMasterXbar__monitor__inflight_1  |(  tlMasterXbar__monitor___GEN_6   ? 2'h1<<  tlMasterXbar__monitor___GEN_5  :2'h0))&~(  tlMasterXbar__monitor___GEN_101   ? 2'h1<<  tlMasterXbar__monitor___GEN_3  :2'h0); 
               tlMasterXbar__monitor__inflight_sizes_1   <=(  tlMasterXbar__monitor__inflight_sizes_1  |(  tlMasterXbar__monitor___GEN_6   ?   tlMasterXbar__monitor___c_sizes_set_T_1  [15:0]:16'h0))&~(  tlMasterXbar__monitor___GEN_101   ?   tlMasterXbar__monitor___d_sizes_clr_T_11  [15:0]:16'h0);
              if (  tlMasterXbar__monitor___c_first_T_1  |  tlMasterXbar__monitor___d_first_T_3  ) 
                  tlMasterXbar__monitor__watchdog_1   <=32'h0;
               else  
                  tlMasterXbar__monitor__watchdog_1   <=  tlMasterXbar__monitor__watchdog_1  +32'h1; 
               tlMasterXbar__monitor__inflight_2   <=(  tlMasterXbar__monitor__inflight_2  |  tlMasterXbar__monitor__d_set  )&~(  tlMasterXbar__monitor___GEN_9   ? 4'h1<<  tlMasterXbar__monitor___GEN_10  :4'h0);
            end 
         if (  tlMasterXbar__monitor___a_first_T_1  &~(|  tlMasterXbar__monitor__a_first_counter  ))
            begin  
               tlMasterXbar__monitor__opcode   <=  tlMasterXbar__monitor__io_in_a_bits_opcode  ; 
               tlMasterXbar__monitor__param   <=  tlMasterXbar__monitor__io_in_a_bits_param  ; 
               tlMasterXbar__monitor__size   <=  tlMasterXbar__monitor__io_in_a_bits_size  ; 
               tlMasterXbar__monitor__source   <=  tlMasterXbar__monitor__io_in_a_bits_source  ; 
               tlMasterXbar__monitor__address   <=  tlMasterXbar__monitor__io_in_a_bits_address  ;
            end 
         if (  tlMasterXbar__monitor___d_first_T_3  &~(|  tlMasterXbar__monitor__d_first_counter  ))
            begin  
               tlMasterXbar__monitor__opcode_1   <=  tlMasterXbar__monitor__io_in_d_bits_opcode  ; 
               tlMasterXbar__monitor__param_1   <=  tlMasterXbar__monitor__io_in_d_bits_param  ; 
               tlMasterXbar__monitor__size_1   <=  tlMasterXbar__monitor__io_in_d_bits_size  ; 
               tlMasterXbar__monitor__source_1   <=  tlMasterXbar__monitor__io_in_d_bits_source  ; 
               tlMasterXbar__monitor__sink   <=  tlMasterXbar__monitor__io_in_d_bits_sink  ; 
               tlMasterXbar__monitor__denied   <=  tlMasterXbar__monitor__io_in_d_bits_denied  ;
            end 
         if (  tlMasterXbar__monitor__b_first_done  &~(|  tlMasterXbar__monitor__b_first_counter  ))
            begin  
               tlMasterXbar__monitor__opcode_2   <=  tlMasterXbar__monitor__io_in_b_bits_opcode  ; 
               tlMasterXbar__monitor__param_2   <=  tlMasterXbar__monitor__io_in_b_bits_param  ; 
               tlMasterXbar__monitor__size_2   <=  tlMasterXbar__monitor__io_in_b_bits_size  ; 
               tlMasterXbar__monitor__source_2   <=  tlMasterXbar__monitor__io_in_b_bits_source  ; 
               tlMasterXbar__monitor__address_1   <=  tlMasterXbar__monitor__io_in_b_bits_address  ;
            end 
         if (  tlMasterXbar__monitor___c_first_T_1  &~(|  tlMasterXbar__monitor__c_first_counter  ))
            begin  
               tlMasterXbar__monitor__opcode_3   <=  tlMasterXbar__monitor__io_in_c_bits_opcode  ; 
               tlMasterXbar__monitor__param_3   <=  tlMasterXbar__monitor__io_in_c_bits_param  ; 
               tlMasterXbar__monitor__size_3   <=  tlMasterXbar__monitor__io_in_c_bits_size  ; 
               tlMasterXbar__monitor__source_3   <=  tlMasterXbar__monitor__io_in_c_bits_source  ; 
               tlMasterXbar__monitor__address_2   <=  tlMasterXbar__monitor__io_in_c_bits_address  ;
            end 
       end
 
assign tlMasterXbar__monitor__clock = tlMasterXbar__clock;
assign tlMasterXbar__monitor__reset = tlMasterXbar__reset;
assign tlMasterXbar__monitor__io_in_a_ready = tlMasterXbar__portsAOI_filtered_0_ready;
assign tlMasterXbar__monitor__io_in_a_valid = tlMasterXbar__auto_in_0_a_valid;
assign tlMasterXbar__monitor__io_in_a_bits_opcode = tlMasterXbar__auto_in_0_a_bits_opcode;
assign tlMasterXbar__monitor__io_in_a_bits_param = tlMasterXbar__auto_in_0_a_bits_param;
assign tlMasterXbar__monitor__io_in_a_bits_size = tlMasterXbar__auto_in_0_a_bits_size;
assign tlMasterXbar__monitor__io_in_a_bits_source = tlMasterXbar__auto_in_0_a_bits_source;
assign tlMasterXbar__monitor__io_in_a_bits_address = tlMasterXbar__auto_in_0_a_bits_address;
assign tlMasterXbar__monitor__io_in_a_bits_mask = tlMasterXbar__auto_in_0_a_bits_mask;
assign tlMasterXbar__monitor__io_in_b_ready = tlMasterXbar__auto_in_0_b_ready;
assign tlMasterXbar__monitor__io_in_b_valid = tlMasterXbar__portsBIO_filtered_valid_0;
assign tlMasterXbar__monitor__io_in_b_bits_opcode = tlMasterXbar__auto_out_b_bits_opcode;
assign tlMasterXbar__monitor__io_in_b_bits_param = tlMasterXbar__auto_out_b_bits_param;
assign tlMasterXbar__monitor__io_in_b_bits_size = tlMasterXbar__auto_out_b_bits_size;
assign tlMasterXbar__monitor__io_in_b_bits_source = tlMasterXbar__auto_out_b_bits_source[0];
assign tlMasterXbar__monitor__io_in_b_bits_address = tlMasterXbar__auto_out_b_bits_address;
assign tlMasterXbar__monitor__io_in_b_bits_mask = tlMasterXbar__auto_out_b_bits_mask;
assign tlMasterXbar__monitor__io_in_b_bits_corrupt = tlMasterXbar__auto_out_b_bits_corrupt;
assign tlMasterXbar__monitor__io_in_c_ready = tlMasterXbar__auto_out_c_ready;
assign tlMasterXbar__monitor__io_in_c_valid = tlMasterXbar__auto_in_0_c_valid;
assign tlMasterXbar__monitor__io_in_c_bits_opcode = tlMasterXbar__auto_in_0_c_bits_opcode;
assign tlMasterXbar__monitor__io_in_c_bits_param = tlMasterXbar__auto_in_0_c_bits_param;
assign tlMasterXbar__monitor__io_in_c_bits_size = tlMasterXbar__auto_in_0_c_bits_size;
assign tlMasterXbar__monitor__io_in_c_bits_source = tlMasterXbar__auto_in_0_c_bits_source;
assign tlMasterXbar__monitor__io_in_c_bits_address = tlMasterXbar__auto_in_0_c_bits_address;
assign tlMasterXbar__monitor__io_in_d_ready = tlMasterXbar__auto_in_0_d_ready;
assign tlMasterXbar__monitor__io_in_d_valid = tlMasterXbar__portsDIO_filtered_0_valid;
assign tlMasterXbar__monitor__io_in_d_bits_opcode = tlMasterXbar__auto_out_d_bits_opcode;
assign tlMasterXbar__monitor__io_in_d_bits_param = tlMasterXbar__auto_out_d_bits_param;
assign tlMasterXbar__monitor__io_in_d_bits_size = tlMasterXbar__auto_out_d_bits_size;
assign tlMasterXbar__monitor__io_in_d_bits_source = tlMasterXbar__auto_out_d_bits_source[0];
assign tlMasterXbar__monitor__io_in_d_bits_sink = tlMasterXbar__auto_out_d_bits_sink;
assign tlMasterXbar__monitor__io_in_d_bits_denied = tlMasterXbar__auto_out_d_bits_denied;
assign tlMasterXbar__monitor__io_in_d_bits_corrupt = tlMasterXbar__auto_out_d_bits_corrupt;
assign tlMasterXbar__monitor__io_in_e_ready = tlMasterXbar__auto_out_e_ready;
assign tlMasterXbar__monitor__io_in_e_valid = tlMasterXbar__auto_in_0_e_valid;
assign tlMasterXbar__monitor__io_in_e_bits_sink = tlMasterXbar__auto_in_0_e_bits_sink;
  
  
wire  tlMasterXbar__monitor_1__clock;
wire  tlMasterXbar__monitor_1__reset;
wire  tlMasterXbar__monitor_1__io_in_a_ready;
wire  tlMasterXbar__monitor_1__io_in_a_valid;
wire [31:0] tlMasterXbar__monitor_1__io_in_a_bits_address;
wire  tlMasterXbar__monitor_1__io_in_d_valid;
wire [2:0] tlMasterXbar__monitor_1__io_in_d_bits_opcode;
wire [1:0] tlMasterXbar__monitor_1__io_in_d_bits_param;
wire [3:0] tlMasterXbar__monitor_1__io_in_d_bits_size;
wire [1:0] tlMasterXbar__monitor_1__io_in_d_bits_sink;
wire  tlMasterXbar__monitor_1__io_in_d_bits_denied;
wire  tlMasterXbar__monitor_1__io_in_d_bits_corrupt;
 
   wire[31:0]  tlMasterXbar__monitor_1___plusarg_reader_1_out  ; 
   wire[31:0]  tlMasterXbar__monitor_1___plusarg_reader_out  ; 
   wire  tlMasterXbar__monitor_1___a_first_T_1  =  tlMasterXbar__monitor_1__io_in_a_ready  &  tlMasterXbar__monitor_1__io_in_a_valid  ; 
   reg[8:0]  tlMasterXbar__monitor_1__a_first_counter  ; 
   reg[31:0]  tlMasterXbar__monitor_1__address  ; 
   reg[8:0]  tlMasterXbar__monitor_1__d_first_counter  ; 
   reg[2:0]  tlMasterXbar__monitor_1__opcode_1  ; 
   reg[1:0]  tlMasterXbar__monitor_1__param_1  ; 
   reg[3:0]  tlMasterXbar__monitor_1__size_1  ; 
   reg[1:0]  tlMasterXbar__monitor_1__sink  ; 
   reg  tlMasterXbar__monitor_1__denied  ; 
   reg  tlMasterXbar__monitor_1__inflight  ; 
   reg[3:0]  tlMasterXbar__monitor_1__inflight_opcodes  ; 
   reg[7:0]  tlMasterXbar__monitor_1__inflight_sizes  ; 
   reg[8:0]  tlMasterXbar__monitor_1__a_first_counter_1  ; 
   wire  tlMasterXbar__monitor_1__a_first_1  =  tlMasterXbar__monitor_1__a_first_counter_1  ==9'h0; 
   reg[8:0]  tlMasterXbar__monitor_1__d_first_counter_1  ; 
   wire  tlMasterXbar__monitor_1__d_first_1  =  tlMasterXbar__monitor_1__d_first_counter_1  ==9'h0; 
   wire  tlMasterXbar__monitor_1__a_set  =  tlMasterXbar__monitor_1___a_first_T_1  &  tlMasterXbar__monitor_1__a_first_1  ; 
   wire  tlMasterXbar__monitor_1__d_release_ack  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h6; 
   wire  tlMasterXbar__monitor_1___GEN  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__d_first_1  ; 
   wire  tlMasterXbar__monitor_1__d_clr  =  tlMasterXbar__monitor_1___GEN  &~  tlMasterXbar__monitor_1__d_release_ack  ; 
   reg[2:0]  tlMasterXbar__monitor_1__casez_tmp  ; 
  always @(*)
       begin 
         casez (  tlMasterXbar__monitor_1__inflight_opcodes  [3:1])
          3 'b000: 
              tlMasterXbar__monitor_1__casez_tmp   =3'h0;
          3 'b001: 
              tlMasterXbar__monitor_1__casez_tmp   =3'h0;
          3 'b010: 
              tlMasterXbar__monitor_1__casez_tmp   =3'h1;
          3 'b011: 
              tlMasterXbar__monitor_1__casez_tmp   =3'h1;
          3 'b100: 
              tlMasterXbar__monitor_1__casez_tmp   =3'h1;
          3 'b101: 
              tlMasterXbar__monitor_1__casez_tmp   =3'h2;
          3 'b110: 
              tlMasterXbar__monitor_1__casez_tmp   =3'h4;
          default : 
              tlMasterXbar__monitor_1__casez_tmp   =3'h4;
         endcase 
       end
  
   reg[2:0]  tlMasterXbar__monitor_1__casez_tmp_0  ; 
  always @(*)
       begin 
         casez (  tlMasterXbar__monitor_1__inflight_opcodes  [3:1])
          3 'b000: 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h0;
          3 'b001: 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h0;
          3 'b010: 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h1;
          3 'b011: 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h1;
          3 'b100: 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h1;
          3 'b101: 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h2;
          3 'b110: 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h5;
          default : 
              tlMasterXbar__monitor_1__casez_tmp_0   =3'h4;
         endcase 
       end
  
   reg[31:0]  tlMasterXbar__monitor_1__watchdog  ; 
   reg  tlMasterXbar__monitor_1__inflight_1  ; 
   reg[7:0]  tlMasterXbar__monitor_1__inflight_sizes_1  ; 
   reg[8:0]  tlMasterXbar__monitor_1__d_first_counter_2  ; 
   wire  tlMasterXbar__monitor_1__d_first_2  =  tlMasterXbar__monitor_1__d_first_counter_2  ==9'h0; 
   wire  tlMasterXbar__monitor_1__d_clr_1  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__d_first_2  &  tlMasterXbar__monitor_1__d_release_ack  ; 
   reg[31:0]  tlMasterXbar__monitor_1__watchdog_1  ; 
   wire  tlMasterXbar__monitor_1___GEN_0  =  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_1  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h6&~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_2  =  tlMasterXbar__monitor_1__io_in_d_bits_size  <4'h3; 
   wire  tlMasterXbar__monitor_1___GEN_3  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h4&~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_4  =  tlMasterXbar__monitor_1__io_in_d_bits_param  ==2'h2; 
   wire  tlMasterXbar__monitor_1___GEN_5  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h5&~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_6  =~  tlMasterXbar__monitor_1__io_in_d_bits_denied  |  tlMasterXbar__monitor_1__io_in_d_bits_corrupt  ; 
   wire  tlMasterXbar__monitor_1___GEN_7  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h0&~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_8  =  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h1; 
   wire  tlMasterXbar__monitor_1___GEN_9  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1___GEN_8  &~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_10  =  tlMasterXbar__monitor_1__io_in_d_valid  &  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==3'h2&~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_11  =  tlMasterXbar__monitor_1__io_in_d_valid  &(|  tlMasterXbar__monitor_1__d_first_counter  )&~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1__a_set_wo_ready  =  tlMasterXbar__monitor_1__io_in_a_valid  &  tlMasterXbar__monitor_1__a_first_1  ; 
   wire  tlMasterXbar__monitor_1___GEN_12  =  tlMasterXbar__monitor_1__d_clr  &  tlMasterXbar__monitor_1__a_set_wo_ready  &~  tlMasterXbar__monitor_1__reset  ; 
   wire  tlMasterXbar__monitor_1___GEN_13  =  tlMasterXbar__monitor_1__d_clr  &~  tlMasterXbar__monitor_1__a_set_wo_ready  &~  tlMasterXbar__monitor_1__reset  ; 
   wire[7:0]  tlMasterXbar__monitor_1___GEN_14  ={4'h0,  tlMasterXbar__monitor_1__io_in_d_bits_size  }; 
   wire  tlMasterXbar__monitor_1___GEN_15  =  tlMasterXbar__monitor_1__d_clr_1  &~  tlMasterXbar__monitor_1__reset  ; 
  always @( posedge   tlMasterXbar__monitor_1__clock  )
       begin 
         if (  tlMasterXbar__monitor_1___GEN_0  &~({  tlMasterXbar__monitor_1__io_in_a_bits_address  [31:14],~(  tlMasterXbar__monitor_1__io_in_a_bits_address  [13:12])}==20'h0|  tlMasterXbar__monitor_1__io_in_a_bits_address  [31:12]==20'h0|{  tlMasterXbar__monitor_1__io_in_a_bits_address  [31:17],~(  tlMasterXbar__monitor_1__io_in_a_bits_address  [16])}==16'h0|{  tlMasterXbar__monitor_1__io_in_a_bits_address  [31:26],  tlMasterXbar__monitor_1__io_in_a_bits_address  [25:16]^10'h200}==16'h0|{  tlMasterXbar__monitor_1__io_in_a_bits_address  [31:28],~(  tlMasterXbar__monitor_1__io_in_a_bits_address  [27:26])}==6'h0|{  tlMasterXbar__monitor_1__io_in_a_bits_address  [31],~(  tlMasterXbar__monitor_1__io_in_a_bits_address  [30:29])}==3'h0|  tlMasterXbar__monitor_1__io_in_a_bits_address  [31:28]==4'h8))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_0  &(|(  tlMasterXbar__monitor_1__io_in_a_bits_address  [5:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1__io_in_d_valid  &~  tlMasterXbar__monitor_1__reset  &(&  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_1  &  tlMasterXbar__monitor_1___GEN_2  )
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_1  &(|  tlMasterXbar__monitor_1__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_1  &  tlMasterXbar__monitor_1__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_1  &  tlMasterXbar__monitor_1__io_in_d_bits_denied  )
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_3  &  tlMasterXbar__monitor_1___GEN_2  )
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_3  &(&  tlMasterXbar__monitor_1__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_3  &  tlMasterXbar__monitor_1___GEN_4  )
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_3  &  tlMasterXbar__monitor_1__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_5  &  tlMasterXbar__monitor_1___GEN_2  )
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_5  &(&  tlMasterXbar__monitor_1__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_5  &  tlMasterXbar__monitor_1___GEN_4  )
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_5  &~  tlMasterXbar__monitor_1___GEN_6  )
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_7  &(|  tlMasterXbar__monitor_1__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_7  &  tlMasterXbar__monitor_1__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_9  &(|  tlMasterXbar__monitor_1__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_9  &~  tlMasterXbar__monitor_1___GEN_6  )
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_10  &(|  tlMasterXbar__monitor_1__io_in_d_bits_param  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_10  &  tlMasterXbar__monitor_1__io_in_d_bits_corrupt  )
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1__io_in_a_valid  &(|  tlMasterXbar__monitor_1__a_first_counter  )&~  tlMasterXbar__monitor_1__reset  &  tlMasterXbar__monitor_1__io_in_a_bits_address  !=  tlMasterXbar__monitor_1__address  )
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_11  &  tlMasterXbar__monitor_1__io_in_d_bits_opcode  !=  tlMasterXbar__monitor_1__opcode_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_11  &  tlMasterXbar__monitor_1__io_in_d_bits_param  !=  tlMasterXbar__monitor_1__param_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_11  &  tlMasterXbar__monitor_1__io_in_d_bits_size  !=  tlMasterXbar__monitor_1__size_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_11  &  tlMasterXbar__monitor_1__io_in_d_bits_sink  !=  tlMasterXbar__monitor_1__sink  )
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_11  &  tlMasterXbar__monitor_1__io_in_d_bits_denied  !=  tlMasterXbar__monitor_1__denied  )
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1__a_set  &~  tlMasterXbar__monitor_1__reset  &  tlMasterXbar__monitor_1__inflight  )
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1__d_clr  &~  tlMasterXbar__monitor_1__reset  &~(  tlMasterXbar__monitor_1__inflight  |  tlMasterXbar__monitor_1__a_set_wo_ready  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_12  &~  tlMasterXbar__monitor_1___GEN_8  )
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_12  &  tlMasterXbar__monitor_1__io_in_d_bits_size  !=4'h6)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_13  &~(  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==  tlMasterXbar__monitor_1__casez_tmp  |  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ==  tlMasterXbar__monitor_1__casez_tmp_0  ))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_13  &  tlMasterXbar__monitor_1___GEN_14  !={1'h0,  tlMasterXbar__monitor_1__inflight_sizes  [7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN  &  tlMasterXbar__monitor_1__a_first_1  &  tlMasterXbar__monitor_1__io_in_a_valid  &~  tlMasterXbar__monitor_1__d_release_ack  &~  tlMasterXbar__monitor_1__reset  &~  tlMasterXbar__monitor_1__io_in_a_ready  )
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~  tlMasterXbar__monitor_1__reset  &~(  tlMasterXbar__monitor_1__a_set_wo_ready  !=  tlMasterXbar__monitor_1__d_clr  |~  tlMasterXbar__monitor_1__a_set_wo_ready  ))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~  tlMasterXbar__monitor_1__reset  &~(~  tlMasterXbar__monitor_1__inflight  |  tlMasterXbar__monitor_1___plusarg_reader_out  ==32'h0|  tlMasterXbar__monitor_1__watchdog  <  tlMasterXbar__monitor_1___plusarg_reader_out  ))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_15  &~  tlMasterXbar__monitor_1__inflight_1  )
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (  tlMasterXbar__monitor_1___GEN_15  &  tlMasterXbar__monitor_1___GEN_14  !={1'h0,  tlMasterXbar__monitor_1__inflight_sizes_1  [7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~  tlMasterXbar__monitor_1__reset  &~(~  tlMasterXbar__monitor_1__inflight_1  |  tlMasterXbar__monitor_1___plusarg_reader_1_out  ==32'h0|  tlMasterXbar__monitor_1__watchdog_1  <  tlMasterXbar__monitor_1___plusarg_reader_1_out  ))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire[26:0]  tlMasterXbar__monitor_1___GEN_16  ={23'h0,  tlMasterXbar__monitor_1__io_in_d_bits_size  }; 
   wire[26:0]  tlMasterXbar__monitor_1___d_first_beats1_decode_T_1  =27'hFFF<<  tlMasterXbar__monitor_1___GEN_16  ; 
   wire[26:0]  tlMasterXbar__monitor_1___d_first_beats1_decode_T_5  =27'hFFF<<  tlMasterXbar__monitor_1___GEN_16  ; 
   wire[26:0]  tlMasterXbar__monitor_1___d_first_beats1_decode_T_9  =27'hFFF<<  tlMasterXbar__monitor_1___GEN_16  ; 
  always @( posedge   tlMasterXbar__monitor_1__clock  )
       begin 
         if (  tlMasterXbar__monitor_1__reset  )
            begin  
               tlMasterXbar__monitor_1__a_first_counter   <=9'h0; 
               tlMasterXbar__monitor_1__d_first_counter   <=9'h0; 
               tlMasterXbar__monitor_1__inflight   <=1'h0; 
               tlMasterXbar__monitor_1__inflight_opcodes   <=4'h0; 
               tlMasterXbar__monitor_1__inflight_sizes   <=8'h0; 
               tlMasterXbar__monitor_1__a_first_counter_1   <=9'h0; 
               tlMasterXbar__monitor_1__d_first_counter_1   <=9'h0; 
               tlMasterXbar__monitor_1__watchdog   <=32'h0; 
               tlMasterXbar__monitor_1__inflight_1   <=1'h0; 
               tlMasterXbar__monitor_1__inflight_sizes_1   <=8'h0; 
               tlMasterXbar__monitor_1__d_first_counter_2   <=9'h0; 
               tlMasterXbar__monitor_1__watchdog_1   <=32'h0;
            end 
          else 
            begin 
              if (  tlMasterXbar__monitor_1___a_first_T_1  )
                 begin 
                   if (|  tlMasterXbar__monitor_1__a_first_counter  ) 
                       tlMasterXbar__monitor_1__a_first_counter   <=  tlMasterXbar__monitor_1__a_first_counter  -9'h1;
                    else  
                       tlMasterXbar__monitor_1__a_first_counter   <=9'h0;
                   if (  tlMasterXbar__monitor_1__a_first_1  ) 
                       tlMasterXbar__monitor_1__a_first_counter_1   <=9'h0;
                    else  
                       tlMasterXbar__monitor_1__a_first_counter_1   <=  tlMasterXbar__monitor_1__a_first_counter_1  -9'h1;
                 end 
              if (  tlMasterXbar__monitor_1__io_in_d_valid  )
                 begin 
                   if (|  tlMasterXbar__monitor_1__d_first_counter  ) 
                       tlMasterXbar__monitor_1__d_first_counter   <=  tlMasterXbar__monitor_1__d_first_counter  -9'h1;
                    else  
                       tlMasterXbar__monitor_1__d_first_counter   <=  tlMasterXbar__monitor_1__io_in_d_bits_opcode  [0] ? ~(  tlMasterXbar__monitor_1___d_first_beats1_decode_T_1  [11:3]):9'h0;
                   if (  tlMasterXbar__monitor_1__d_first_1  ) 
                       tlMasterXbar__monitor_1__d_first_counter_1   <=  tlMasterXbar__monitor_1__io_in_d_bits_opcode  [0] ? ~(  tlMasterXbar__monitor_1___d_first_beats1_decode_T_5  [11:3]):9'h0;
                    else  
                       tlMasterXbar__monitor_1__d_first_counter_1   <=  tlMasterXbar__monitor_1__d_first_counter_1  -9'h1;
                   if (  tlMasterXbar__monitor_1__d_first_2  ) 
                       tlMasterXbar__monitor_1__d_first_counter_2   <=  tlMasterXbar__monitor_1__io_in_d_bits_opcode  [0] ? ~(  tlMasterXbar__monitor_1___d_first_beats1_decode_T_9  [11:3]):9'h0;
                    else  
                       tlMasterXbar__monitor_1__d_first_counter_2   <=  tlMasterXbar__monitor_1__d_first_counter_2  -9'h1; 
                    tlMasterXbar__monitor_1__watchdog_1   <=32'h0;
                 end 
               else  
                  tlMasterXbar__monitor_1__watchdog_1   <=  tlMasterXbar__monitor_1__watchdog_1  +32'h1; 
               tlMasterXbar__monitor_1__inflight   <=(  tlMasterXbar__monitor_1__inflight  |  tlMasterXbar__monitor_1__a_set  )&~  tlMasterXbar__monitor_1__d_clr  ; 
               tlMasterXbar__monitor_1__inflight_opcodes   <=(  tlMasterXbar__monitor_1__inflight_opcodes  |(  tlMasterXbar__monitor_1__a_set   ? 4'h9:4'h0))&~{4{  tlMasterXbar__monitor_1__d_clr  }}; 
               tlMasterXbar__monitor_1__inflight_sizes   <=(  tlMasterXbar__monitor_1__inflight_sizes  |(  tlMasterXbar__monitor_1__a_set   ? {3'h0,  tlMasterXbar__monitor_1__a_set   ? 5'hD:5'h0}:8'h0))&~{8{  tlMasterXbar__monitor_1__d_clr  }};
              if (  tlMasterXbar__monitor_1___a_first_T_1  |  tlMasterXbar__monitor_1__io_in_d_valid  ) 
                  tlMasterXbar__monitor_1__watchdog   <=32'h0;
               else  
                  tlMasterXbar__monitor_1__watchdog   <=  tlMasterXbar__monitor_1__watchdog  +32'h1; 
               tlMasterXbar__monitor_1__inflight_1   <=  tlMasterXbar__monitor_1__inflight_1  &~  tlMasterXbar__monitor_1__d_clr_1  ; 
               tlMasterXbar__monitor_1__inflight_sizes_1   <=  tlMasterXbar__monitor_1__inflight_sizes_1  &~{8{  tlMasterXbar__monitor_1__d_clr_1  }};
            end 
         if (  tlMasterXbar__monitor_1___a_first_T_1  &~(|  tlMasterXbar__monitor_1__a_first_counter  )) 
             tlMasterXbar__monitor_1__address   <=  tlMasterXbar__monitor_1__io_in_a_bits_address  ;
         if (  tlMasterXbar__monitor_1__io_in_d_valid  &~(|  tlMasterXbar__monitor_1__d_first_counter  ))
            begin  
               tlMasterXbar__monitor_1__opcode_1   <=  tlMasterXbar__monitor_1__io_in_d_bits_opcode  ; 
               tlMasterXbar__monitor_1__param_1   <=  tlMasterXbar__monitor_1__io_in_d_bits_param  ; 
               tlMasterXbar__monitor_1__size_1   <=  tlMasterXbar__monitor_1__io_in_d_bits_size  ; 
               tlMasterXbar__monitor_1__sink   <=  tlMasterXbar__monitor_1__io_in_d_bits_sink  ; 
               tlMasterXbar__monitor_1__denied   <=  tlMasterXbar__monitor_1__io_in_d_bits_denied  ;
            end 
       end
 
assign tlMasterXbar__monitor_1__clock = tlMasterXbar__clock;
assign tlMasterXbar__monitor_1__reset = tlMasterXbar__reset;
assign tlMasterXbar__monitor_1__io_in_a_ready = tlMasterXbar__portsAOI_filtered_1_0_ready;
assign tlMasterXbar__monitor_1__io_in_a_valid = tlMasterXbar__auto_in_1_a_valid;
assign tlMasterXbar__monitor_1__io_in_a_bits_address = tlMasterXbar__auto_in_1_a_bits_address;
assign tlMasterXbar__monitor_1__io_in_d_valid = tlMasterXbar__portsDIO_filtered_1_valid;
assign tlMasterXbar__monitor_1__io_in_d_bits_opcode = tlMasterXbar__auto_out_d_bits_opcode;
assign tlMasterXbar__monitor_1__io_in_d_bits_param = tlMasterXbar__auto_out_d_bits_param;
assign tlMasterXbar__monitor_1__io_in_d_bits_size = tlMasterXbar__auto_out_d_bits_size;
assign tlMasterXbar__monitor_1__io_in_d_bits_sink = tlMasterXbar__auto_out_d_bits_sink;
assign tlMasterXbar__monitor_1__io_in_d_bits_denied = tlMasterXbar__auto_out_d_bits_denied;
assign tlMasterXbar__monitor_1__io_in_d_bits_corrupt = tlMasterXbar__auto_out_d_bits_corrupt;
 
  assign   tlMasterXbar__auto_in_1_a_ready  =  tlMasterXbar__portsAOI_filtered_1_0_ready  ; 
  assign   tlMasterXbar__auto_in_1_d_valid  =  tlMasterXbar__portsDIO_filtered_1_valid  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_opcode  =  tlMasterXbar__auto_out_d_bits_opcode  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_size  =  tlMasterXbar__auto_out_d_bits_size  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_data  =  tlMasterXbar__auto_out_d_bits_data  ; 
  assign   tlMasterXbar__auto_in_1_d_bits_corrupt  =  tlMasterXbar__auto_out_d_bits_corrupt  ; 
  assign   tlMasterXbar__auto_in_0_a_ready  =  tlMasterXbar__portsAOI_filtered_0_ready  ; 
  assign   tlMasterXbar__auto_in_0_b_valid  =  tlMasterXbar__portsBIO_filtered_valid_0  ; 
  assign   tlMasterXbar__auto_in_0_b_bits_param  =  tlMasterXbar__auto_out_b_bits_param  ; 
  assign   tlMasterXbar__auto_in_0_b_bits_size  =  tlMasterXbar__auto_out_b_bits_size  ; 
  assign   tlMasterXbar__auto_in_0_b_bits_source  =  tlMasterXbar__auto_out_b_bits_source  [0]; 
  assign   tlMasterXbar__auto_in_0_b_bits_address  =  tlMasterXbar__auto_out_b_bits_address  ; 
  assign   tlMasterXbar__auto_in_0_c_ready  =  tlMasterXbar__auto_out_c_ready  ; 
  assign   tlMasterXbar__auto_in_0_d_valid  =  tlMasterXbar__portsDIO_filtered_0_valid  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_opcode  =  tlMasterXbar__auto_out_d_bits_opcode  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_param  =  tlMasterXbar__auto_out_d_bits_param  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_size  =  tlMasterXbar__auto_out_d_bits_size  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_source  =  tlMasterXbar__auto_out_d_bits_source  [0]; 
  assign   tlMasterXbar__auto_in_0_d_bits_sink  =  tlMasterXbar__auto_out_d_bits_sink  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_denied  =  tlMasterXbar__auto_out_d_bits_denied  ; 
  assign   tlMasterXbar__auto_in_0_d_bits_data  =  tlMasterXbar__auto_out_d_bits_data  ; 
  assign   tlMasterXbar__auto_in_0_e_ready  =  tlMasterXbar__auto_out_e_ready  ; 
  assign   tlMasterXbar__auto_out_a_valid  =  tlMasterXbar__out_0_a_valid  ; 
  assign   tlMasterXbar__auto_out_a_bits_opcode  =(  tlMasterXbar__muxState_0   ?   tlMasterXbar__auto_in_0_a_bits_opcode  :3'h0)|{  tlMasterXbar__muxState_1  ,2'h0}; 
  assign   tlMasterXbar__auto_out_a_bits_param  =  tlMasterXbar__muxState_0   ?   tlMasterXbar__auto_in_0_a_bits_param  :3'h0; 
  assign   tlMasterXbar__auto_out_a_bits_size  =(  tlMasterXbar__muxState_0   ?   tlMasterXbar__auto_in_0_a_bits_size  :4'h0)|(  tlMasterXbar__muxState_1   ? 4'h6:4'h0); 
  assign   tlMasterXbar__auto_out_a_bits_source  =(  tlMasterXbar__muxState_0   ? {1'h0,  tlMasterXbar__auto_in_0_a_bits_source  }:2'h0)|{  tlMasterXbar__muxState_1  ,1'h0}; 
  assign   tlMasterXbar__auto_out_a_bits_address  =(  tlMasterXbar__muxState_0   ?   tlMasterXbar__auto_in_0_a_bits_address  :32'h0)|(  tlMasterXbar__muxState_1   ?   tlMasterXbar__auto_in_1_a_bits_address  :32'h0); 
  assign   tlMasterXbar__auto_out_a_bits_mask  =(  tlMasterXbar__muxState_0   ?   tlMasterXbar__auto_in_0_a_bits_mask  :8'h0)|{8{  tlMasterXbar__muxState_1  }}; 
  assign   tlMasterXbar__auto_out_a_bits_data  =  tlMasterXbar__muxState_0   ?   tlMasterXbar__auto_in_0_a_bits_data  :64'h0; 
  assign   tlMasterXbar__auto_out_b_ready  =~(  tlMasterXbar__auto_out_b_bits_source  [1])&  tlMasterXbar__auto_in_0_b_ready  ; 
  assign   tlMasterXbar__auto_out_c_valid  =  tlMasterXbar__auto_in_0_c_valid  ; 
  assign   tlMasterXbar__auto_out_c_bits_opcode  =  tlMasterXbar__auto_in_0_c_bits_opcode  ; 
  assign   tlMasterXbar__auto_out_c_bits_param  =  tlMasterXbar__auto_in_0_c_bits_param  ; 
  assign   tlMasterXbar__auto_out_c_bits_size  =  tlMasterXbar__auto_in_0_c_bits_size  ; 
  assign   tlMasterXbar__auto_out_c_bits_source  ={1'h0,  tlMasterXbar__auto_in_0_c_bits_source  }; 
  assign   tlMasterXbar__auto_out_c_bits_address  =  tlMasterXbar__auto_in_0_c_bits_address  ; 
  assign   tlMasterXbar__auto_out_c_bits_data  =  tlMasterXbar__auto_in_0_c_bits_data  ; 
  assign   tlMasterXbar__auto_out_d_ready  =~(  tlMasterXbar__auto_out_d_bits_source  [1])&  tlMasterXbar__auto_in_0_d_ready  |  tlMasterXbar__requestDOI_0_1  ; 
  assign   tlMasterXbar__auto_out_e_valid  =  tlMasterXbar__auto_in_0_e_valid  ; 
  assign   tlMasterXbar__auto_out_e_bits_sink  =  tlMasterXbar__auto_in_0_e_bits_sink  ;
assign tlMasterXbar__clock = clock;
assign tlMasterXbar__reset = reset;
assign _tlMasterXbar_auto_in_1_a_ready = tlMasterXbar__auto_in_1_a_ready;
assign tlMasterXbar__auto_in_1_a_valid = _frontend_auto_icache_master_out_a_valid;
assign tlMasterXbar__auto_in_1_a_bits_address = _frontend_auto_icache_master_out_a_bits_address;
assign _tlMasterXbar_auto_in_1_d_valid = tlMasterXbar__auto_in_1_d_valid;
assign _tlMasterXbar_auto_in_1_d_bits_opcode = tlMasterXbar__auto_in_1_d_bits_opcode;
assign _tlMasterXbar_auto_in_1_d_bits_size = tlMasterXbar__auto_in_1_d_bits_size;
assign _tlMasterXbar_auto_in_1_d_bits_data = tlMasterXbar__auto_in_1_d_bits_data;
assign _tlMasterXbar_auto_in_1_d_bits_corrupt = tlMasterXbar__auto_in_1_d_bits_corrupt;
assign _tlMasterXbar_auto_in_0_a_ready = tlMasterXbar__auto_in_0_a_ready;
assign tlMasterXbar__auto_in_0_a_valid = _dcache_auto_out_a_valid;
assign tlMasterXbar__auto_in_0_a_bits_opcode = _dcache_auto_out_a_bits_opcode;
assign tlMasterXbar__auto_in_0_a_bits_param = _dcache_auto_out_a_bits_param;
assign tlMasterXbar__auto_in_0_a_bits_size = _dcache_auto_out_a_bits_size;
assign tlMasterXbar__auto_in_0_a_bits_source = _dcache_auto_out_a_bits_source;
assign tlMasterXbar__auto_in_0_a_bits_address = _dcache_auto_out_a_bits_address;
assign tlMasterXbar__auto_in_0_a_bits_mask = _dcache_auto_out_a_bits_mask;
assign tlMasterXbar__auto_in_0_a_bits_data = _dcache_auto_out_a_bits_data;
assign tlMasterXbar__auto_in_0_b_ready = _dcache_auto_out_b_ready;
assign _tlMasterXbar_auto_in_0_b_valid = tlMasterXbar__auto_in_0_b_valid;
assign _tlMasterXbar_auto_in_0_b_bits_param = tlMasterXbar__auto_in_0_b_bits_param;
assign _tlMasterXbar_auto_in_0_b_bits_size = tlMasterXbar__auto_in_0_b_bits_size;
assign _tlMasterXbar_auto_in_0_b_bits_source = tlMasterXbar__auto_in_0_b_bits_source;
assign _tlMasterXbar_auto_in_0_b_bits_address = tlMasterXbar__auto_in_0_b_bits_address;
assign _tlMasterXbar_auto_in_0_c_ready = tlMasterXbar__auto_in_0_c_ready;
assign tlMasterXbar__auto_in_0_c_valid = _dcache_auto_out_c_valid;
assign tlMasterXbar__auto_in_0_c_bits_opcode = _dcache_auto_out_c_bits_opcode;
assign tlMasterXbar__auto_in_0_c_bits_param = _dcache_auto_out_c_bits_param;
assign tlMasterXbar__auto_in_0_c_bits_size = _dcache_auto_out_c_bits_size;
assign tlMasterXbar__auto_in_0_c_bits_source = _dcache_auto_out_c_bits_source;
assign tlMasterXbar__auto_in_0_c_bits_address = _dcache_auto_out_c_bits_address;
assign tlMasterXbar__auto_in_0_c_bits_data = _dcache_auto_out_c_bits_data;
assign tlMasterXbar__auto_in_0_d_ready = _dcache_auto_out_d_ready;
assign _tlMasterXbar_auto_in_0_d_valid = tlMasterXbar__auto_in_0_d_valid;
assign _tlMasterXbar_auto_in_0_d_bits_opcode = tlMasterXbar__auto_in_0_d_bits_opcode;
assign _tlMasterXbar_auto_in_0_d_bits_param = tlMasterXbar__auto_in_0_d_bits_param;
assign _tlMasterXbar_auto_in_0_d_bits_size = tlMasterXbar__auto_in_0_d_bits_size;
assign _tlMasterXbar_auto_in_0_d_bits_source = tlMasterXbar__auto_in_0_d_bits_source;
assign _tlMasterXbar_auto_in_0_d_bits_sink = tlMasterXbar__auto_in_0_d_bits_sink;
assign _tlMasterXbar_auto_in_0_d_bits_denied = tlMasterXbar__auto_in_0_d_bits_denied;
assign _tlMasterXbar_auto_in_0_d_bits_data = tlMasterXbar__auto_in_0_d_bits_data;
assign _tlMasterXbar_auto_in_0_e_ready = tlMasterXbar__auto_in_0_e_ready;
assign tlMasterXbar__auto_in_0_e_valid = _dcache_auto_out_e_valid;
assign tlMasterXbar__auto_in_0_e_bits_sink = _dcache_auto_out_e_bits_sink;
assign tlMasterXbar__auto_out_a_ready = auto_buffer_out_a_ready;
assign auto_buffer_out_a_valid = tlMasterXbar__auto_out_a_valid;
assign auto_buffer_out_a_bits_opcode = tlMasterXbar__auto_out_a_bits_opcode;
assign auto_buffer_out_a_bits_param = tlMasterXbar__auto_out_a_bits_param;
assign auto_buffer_out_a_bits_size = tlMasterXbar__auto_out_a_bits_size;
assign auto_buffer_out_a_bits_source = tlMasterXbar__auto_out_a_bits_source;
assign auto_buffer_out_a_bits_address = tlMasterXbar__auto_out_a_bits_address;
assign auto_buffer_out_a_bits_mask = tlMasterXbar__auto_out_a_bits_mask;
assign auto_buffer_out_a_bits_data = tlMasterXbar__auto_out_a_bits_data;
assign auto_buffer_out_b_ready = tlMasterXbar__auto_out_b_ready;
assign tlMasterXbar__auto_out_b_valid = auto_buffer_out_b_valid;
assign tlMasterXbar__auto_out_b_bits_opcode = auto_buffer_out_b_bits_opcode;
assign tlMasterXbar__auto_out_b_bits_param = auto_buffer_out_b_bits_param;
assign tlMasterXbar__auto_out_b_bits_size = auto_buffer_out_b_bits_size;
assign tlMasterXbar__auto_out_b_bits_source = auto_buffer_out_b_bits_source;
assign tlMasterXbar__auto_out_b_bits_address = auto_buffer_out_b_bits_address;
assign tlMasterXbar__auto_out_b_bits_mask = auto_buffer_out_b_bits_mask;
assign tlMasterXbar__auto_out_b_bits_corrupt = auto_buffer_out_b_bits_corrupt;
assign tlMasterXbar__auto_out_c_ready = auto_buffer_out_c_ready;
assign auto_buffer_out_c_valid = tlMasterXbar__auto_out_c_valid;
assign auto_buffer_out_c_bits_opcode = tlMasterXbar__auto_out_c_bits_opcode;
assign auto_buffer_out_c_bits_param = tlMasterXbar__auto_out_c_bits_param;
assign auto_buffer_out_c_bits_size = tlMasterXbar__auto_out_c_bits_size;
assign auto_buffer_out_c_bits_source = tlMasterXbar__auto_out_c_bits_source;
assign auto_buffer_out_c_bits_address = tlMasterXbar__auto_out_c_bits_address;
assign auto_buffer_out_c_bits_data = tlMasterXbar__auto_out_c_bits_data;
assign auto_buffer_out_d_ready = tlMasterXbar__auto_out_d_ready;
assign tlMasterXbar__auto_out_d_valid = auto_buffer_out_d_valid;
assign tlMasterXbar__auto_out_d_bits_opcode = auto_buffer_out_d_bits_opcode;
assign tlMasterXbar__auto_out_d_bits_param = auto_buffer_out_d_bits_param;
assign tlMasterXbar__auto_out_d_bits_size = auto_buffer_out_d_bits_size;
assign tlMasterXbar__auto_out_d_bits_source = auto_buffer_out_d_bits_source;
assign tlMasterXbar__auto_out_d_bits_sink = auto_buffer_out_d_bits_sink;
assign tlMasterXbar__auto_out_d_bits_denied = auto_buffer_out_d_bits_denied;
assign tlMasterXbar__auto_out_d_bits_data = auto_buffer_out_d_bits_data;
assign tlMasterXbar__auto_out_d_bits_corrupt = auto_buffer_out_d_bits_corrupt;
assign tlMasterXbar__auto_out_e_ready = auto_buffer_out_e_ready;
assign auto_buffer_out_e_valid = tlMasterXbar__auto_out_e_valid;
assign auto_buffer_out_e_bits_sink = tlMasterXbar__auto_out_e_bits_sink;
 
  
wire  intXbar__auto_int_in_2_0;
wire  intXbar__auto_int_in_1_0;
wire  intXbar__auto_int_in_1_1;
wire  intXbar__auto_int_in_0_0;
wire  intXbar__auto_int_out_0;
wire  intXbar__auto_int_out_1;
wire  intXbar__auto_int_out_2;
wire  intXbar__auto_int_out_3;
 
  assign   intXbar__auto_int_out_0  =  intXbar__auto_int_in_0_0  ; 
  assign   intXbar__auto_int_out_1  =  intXbar__auto_int_in_1_0  ; 
  assign   intXbar__auto_int_out_2  =  intXbar__auto_int_in_1_1  ; 
  assign   intXbar__auto_int_out_3  =  intXbar__auto_int_in_2_0  ;
assign intXbar__auto_int_in_2_0 = auto_int_local_in_2_0;
assign intXbar__auto_int_in_1_0 = auto_int_local_in_1_0;
assign intXbar__auto_int_in_1_1 = auto_int_local_in_1_1;
assign intXbar__auto_int_in_0_0 = auto_int_local_in_0_0;
assign _intXbar_auto_int_out_0 = intXbar__auto_int_out_0;
assign _intXbar_auto_int_out_1 = intXbar__auto_int_out_1;
assign _intXbar_auto_int_out_2 = intXbar__auto_int_out_2;
assign _intXbar_auto_int_out_3 = intXbar__auto_int_out_3;
 
  
wire  dcache__clock;
wire  dcache__reset;
wire  dcache__auto_out_a_ready;
wire  dcache__auto_out_a_valid;
wire [2:0] dcache__auto_out_a_bits_opcode;
wire [2:0] dcache__auto_out_a_bits_param;
wire [3:0] dcache__auto_out_a_bits_size;
wire  dcache__auto_out_a_bits_source;
wire [31:0] dcache__auto_out_a_bits_address;
wire [7:0] dcache__auto_out_a_bits_mask;
wire [63:0] dcache__auto_out_a_bits_data;
wire  dcache__auto_out_b_ready;
wire  dcache__auto_out_b_valid;
wire [1:0] dcache__auto_out_b_bits_param;
wire [3:0] dcache__auto_out_b_bits_size;
wire  dcache__auto_out_b_bits_source;
wire [31:0] dcache__auto_out_b_bits_address;
wire  dcache__auto_out_c_ready;
wire  dcache__auto_out_c_valid;
wire [2:0] dcache__auto_out_c_bits_opcode;
wire [2:0] dcache__auto_out_c_bits_param;
wire [3:0] dcache__auto_out_c_bits_size;
wire  dcache__auto_out_c_bits_source;
wire [31:0] dcache__auto_out_c_bits_address;
wire [63:0] dcache__auto_out_c_bits_data;
wire  dcache__auto_out_d_ready;
wire  dcache__auto_out_d_valid;
wire [2:0] dcache__auto_out_d_bits_opcode;
wire [1:0] dcache__auto_out_d_bits_param;
wire [3:0] dcache__auto_out_d_bits_size;
wire  dcache__auto_out_d_bits_source;
wire [1:0] dcache__auto_out_d_bits_sink;
wire  dcache__auto_out_d_bits_denied;
wire [63:0] dcache__auto_out_d_bits_data;
wire  dcache__auto_out_e_ready;
wire  dcache__auto_out_e_valid;
wire [1:0] dcache__auto_out_e_bits_sink;
wire  dcache__io_cpu_req_ready;
wire  dcache__io_cpu_req_valid;
wire [33:0] dcache__io_cpu_req_bits_addr;
wire [5:0] dcache__io_cpu_req_bits_tag;
wire [4:0] dcache__io_cpu_req_bits_cmd;
wire [1:0] dcache__io_cpu_req_bits_size;
wire  dcache__io_cpu_req_bits_signed;
wire  dcache__io_cpu_req_bits_dv;
wire  dcache__io_cpu_s1_kill;
wire [63:0] dcache__io_cpu_s1_data_data;
wire [7:0] dcache__io_cpu_s1_data_mask;
wire  dcache__io_cpu_s2_nack;
wire  dcache__io_cpu_resp_valid;
wire [33:0] dcache__io_cpu_resp_bits_addr;
wire [5:0] dcache__io_cpu_resp_bits_tag;
wire [4:0] dcache__io_cpu_resp_bits_cmd;
wire [1:0] dcache__io_cpu_resp_bits_size;
wire  dcache__io_cpu_resp_bits_signed;
wire [1:0] dcache__io_cpu_resp_bits_dprv;
wire  dcache__io_cpu_resp_bits_dv;
wire [63:0] dcache__io_cpu_resp_bits_data;
wire [7:0] dcache__io_cpu_resp_bits_mask;
wire  dcache__io_cpu_resp_bits_replay;
wire  dcache__io_cpu_resp_bits_has_data;
wire [63:0] dcache__io_cpu_resp_bits_data_word_bypass;
wire [63:0] dcache__io_cpu_resp_bits_data_raw;
wire [63:0] dcache__io_cpu_resp_bits_store_data;
wire  dcache__io_cpu_replay_next;
wire  dcache__io_cpu_s2_xcpt_ma_ld;
wire  dcache__io_cpu_s2_xcpt_ma_st;
wire  dcache__io_cpu_s2_xcpt_pf_ld;
wire  dcache__io_cpu_s2_xcpt_pf_st;
wire  dcache__io_cpu_s2_xcpt_ae_ld;
wire  dcache__io_cpu_s2_xcpt_ae_st;
wire  dcache__io_cpu_ordered;
wire  dcache__io_cpu_perf_release;
wire  dcache__io_cpu_perf_grant;
wire  dcache__io_ptw_req_bits_bits_need_gpa;
wire  dcache__io_ptw_req_bits_bits_stage2;
wire  dcache__io_ptw_status_debug;
wire  dcache__io_ptw_pmp_cfg_l_0;
wire  dcache__io_ptw_pmp_cfg_l_1;
wire  dcache__io_ptw_pmp_cfg_l_2;
wire  dcache__io_ptw_pmp_cfg_l_3;
wire  dcache__io_ptw_pmp_cfg_l_4;
wire  dcache__io_ptw_pmp_cfg_l_5;
wire  dcache__io_ptw_pmp_cfg_l_6;
wire  dcache__io_ptw_pmp_cfg_l_7;
wire [1:0] dcache__io_ptw_pmp_cfg_a_0;
wire [1:0] dcache__io_ptw_pmp_cfg_a_1;
wire [1:0] dcache__io_ptw_pmp_cfg_a_2;
wire [1:0] dcache__io_ptw_pmp_cfg_a_3;
wire [1:0] dcache__io_ptw_pmp_cfg_a_4;
wire [1:0] dcache__io_ptw_pmp_cfg_a_5;
wire [1:0] dcache__io_ptw_pmp_cfg_a_6;
wire [1:0] dcache__io_ptw_pmp_cfg_a_7;
wire  dcache__io_ptw_pmp_cfg_w_0;
wire  dcache__io_ptw_pmp_cfg_w_1;
wire  dcache__io_ptw_pmp_cfg_w_2;
wire  dcache__io_ptw_pmp_cfg_w_3;
wire  dcache__io_ptw_pmp_cfg_w_4;
wire  dcache__io_ptw_pmp_cfg_w_5;
wire  dcache__io_ptw_pmp_cfg_w_6;
wire  dcache__io_ptw_pmp_cfg_w_7;
wire  dcache__io_ptw_pmp_cfg_r_0;
wire  dcache__io_ptw_pmp_cfg_r_1;
wire  dcache__io_ptw_pmp_cfg_r_2;
wire  dcache__io_ptw_pmp_cfg_r_3;
wire  dcache__io_ptw_pmp_cfg_r_4;
wire  dcache__io_ptw_pmp_cfg_r_5;
wire  dcache__io_ptw_pmp_cfg_r_6;
wire  dcache__io_ptw_pmp_cfg_r_7;
wire [29:0] dcache__io_ptw_pmp_addr_0;
wire [29:0] dcache__io_ptw_pmp_addr_1;
wire [29:0] dcache__io_ptw_pmp_addr_2;
wire [29:0] dcache__io_ptw_pmp_addr_3;
wire [29:0] dcache__io_ptw_pmp_addr_4;
wire [29:0] dcache__io_ptw_pmp_addr_5;
wire [29:0] dcache__io_ptw_pmp_addr_6;
wire [29:0] dcache__io_ptw_pmp_addr_7;
wire [31:0] dcache__io_ptw_pmp_mask_0;
wire [31:0] dcache__io_ptw_pmp_mask_1;
wire [31:0] dcache__io_ptw_pmp_mask_2;
wire [31:0] dcache__io_ptw_pmp_mask_3;
wire [31:0] dcache__io_ptw_pmp_mask_4;
wire [31:0] dcache__io_ptw_pmp_mask_5;
wire [31:0] dcache__io_ptw_pmp_mask_6;
wire [31:0] dcache__io_ptw_pmp_mask_7;
 
   wire  dcache__io_cpu_s2_xcpt_ma_st_0  ; 
   wire  dcache__io_cpu_s2_xcpt_ma_ld_0  ; 
   wire  dcache__io_cpu_s2_xcpt_ae_st_0  ; 
   wire  dcache__io_cpu_s2_xcpt_ae_ld_0  ; 
   wire  dcache__io_cpu_s2_xcpt_pf_st_0  ; 
   wire  dcache__io_cpu_s2_xcpt_pf_ld_0  ; 
   wire[21:0]  dcache__metaArb_io_in_bits_data_7  ; 
   wire  dcache__metaArb_io_in_valid_4  ; 
   wire[11:0]  dcache__dataArb_io_in_bits_addr_2  ; 
   wire  dcache__dataArb_io_in_valid_2  ; 
   wire[3:0]  dcache__nodeOut_c_bits_size  ; 
   wire[2:0]  dcache__nodeOut_c_bits_opcode  ; 
   wire  dcache__nodeOut_c_valid  ; 
   wire[5:0]  dcache__metaArb_io_in_bits_idx_6  ; 
   wire  dcache__metaArb_io_in_valid_6  ; 
   wire  dcache__s1_nack  ; 
   wire  dcache__dataArb_io_in_bits_write_1  ; 
   wire  dcache__dataArb_io_in_valid_1  ; 
   wire  dcache__nodeOut_d_ready  ; 
   wire[21:0]  dcache__metaArb_io_in_bits_data_3  ; 
   wire  dcache__metaArb_io_in_valid_3  ; 
   wire[11:0]  dcache__dataArb_io_in_bits_addr_1  ; 
   wire[7:0]  dcache__dataArb_io_in_bits_eccMask_0  ; 
   wire[63:0]  dcache__dataArb_io_in_bits_wdata_0  ; 
   wire[11:0]  dcache___dataArb_io_in_0_bits_wordMask_wordMask_T  ; 
   wire  dcache__dataArb_io_in_valid_0  ; 
   wire  dcache__pstore_drain  ; 
   wire[21:0]  dcache__metaArb_io_in_bits_data_2  ; 
   wire[5:0]  dcache__metaArb_io_in_bits_idx_3  ; 
   wire[5:0]  dcache__metaArb_io_in_bits_idx_4  ; 
   wire  dcache__metaArb_io_in_valid_2  ; 
   reg[33:0]  dcache__s2_req_addr  ; 
   wire  dcache__readEnable  ; 
   wire  dcache__writeEnable  ; 
   wire[5:0]  dcache__metaArb_io_in_bits_idx_7  ; 
   wire[11:0]  dcache__dataArb_io_in_bits_addr_3  ; 
   wire  dcache__dataArb_io_in_valid_3  ; 
   reg[5:0]  dcache__flushCounter  ; 
   reg  dcache__resetting  ; 
   reg[33:0]  dcache__s1_tlb_req_vaddr  ; 
   wire[63:0]  dcache___amoalus_0_io_out  ; 
   wire[63:0]  dcache___data_io_resp_0  ; 
   wire[21:0]  dcache___tag_array_0_ext_RW0_rdata  ; 
   wire  dcache___tlb_pmp_io_r  ; 
   wire  dcache___tlb_pmp_io_w  ; 
   wire  dcache___GEN  =  dcache__metaArb_io_in_valid_2  |  dcache__metaArb_io_in_valid_3  ; 
   wire  dcache__metaArb_io_out_bits_write  =  dcache__resetting  |  dcache__metaArb_io_in_valid_2  |  dcache__metaArb_io_in_valid_3  |  dcache__metaArb_io_in_valid_4  ; 
   wire  dcache__metaArb__grant_T_2  =  dcache__resetting  |  dcache__metaArb_io_in_valid_2  |  dcache__metaArb_io_in_valid_3  ; 
   wire  dcache__metaArb__grant_T_3  =  dcache__metaArb__grant_T_2  |  dcache__metaArb_io_in_valid_4  ; 
   wire  dcache__metaArb__grant_T_5  =  dcache__metaArb__grant_T_3  |  dcache__metaArb_io_in_valid_6  ; 
   wire  dcache__metaArb_io_out_valid  =  dcache__metaArb__grant_T_5  |  dcache__io_cpu_req_valid  ; 
   wire  dcache__dataArb__grant_T  =  dcache__dataArb_io_in_valid_0  |  dcache__dataArb_io_in_valid_1  ; 
   wire  dcache__dataArb__grant_T_1  =  dcache__dataArb__grant_T  |  dcache__dataArb_io_in_valid_2  ; 
   wire  dcache__dataArb_io_out_valid  =  dcache__dataArb__grant_T_1  |  dcache__dataArb_io_in_valid_3  ; 
   reg  dcache__s1_valid  ; 
   reg  dcache__s1_probe  ; 
   reg[1:0]  dcache__probe_bits_param  ; 
   reg[3:0]  dcache__probe_bits_size  ; 
   reg  dcache__probe_bits_source  ; 
   reg[31:0]  dcache__probe_bits_address  ; 
   wire  dcache__s1_valid_masked  =  dcache__s1_valid  &~  dcache__io_cpu_s1_kill  ; 
   reg[33:0]  dcache__s1_vaddr  ; 
   reg[5:0]  dcache__s1_req_tag  ; 
   reg[4:0]  dcache__s1_req_cmd  ; 
   reg[1:0]  dcache__s1_req_size  ; 
   reg  dcache__s1_req_signed  ; 
   reg[1:0]  dcache__s1_req_dprv  ; 
   reg  dcache__s1_req_dv  ; 
   reg[1:0]  dcache__s1_tlb_req_size  ; 
   reg[4:0]  dcache__s1_tlb_req_cmd  ; 
   reg[1:0]  dcache__s1_tlb_req_prv  ; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_1  =  dcache__s1_req_cmd  ==5'h0; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_2  =  dcache__s1_req_cmd  ==5'h10; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_3  =  dcache__s1_req_cmd  ==5'h6; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_29  =  dcache__s1_req_cmd  ==5'h7; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_31  =  dcache__s1_req_cmd  ==5'h4; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_32  =  dcache__s1_req_cmd  ==5'h9; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_33  =  dcache__s1_req_cmd  ==5'hA; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_34  =  dcache__s1_req_cmd  ==5'hB; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_38  =  dcache__s1_req_cmd  ==5'h8; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_39  =  dcache__s1_req_cmd  ==5'hC; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_40  =  dcache__s1_req_cmd  ==5'hD; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_41  =  dcache__s1_req_cmd  ==5'hE; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_42  =  dcache__s1_req_cmd  ==5'hF; 
   wire  dcache__s1_read  =  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_1  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_2  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_3  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_29  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_31  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_32  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_33  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_34  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_38  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_39  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_40  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_41  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_42  ; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_26  =  dcache__s1_req_cmd  ==5'h1; 
   wire  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_51  =  dcache__s1_req_cmd  ==5'h11; 
   wire  dcache__s1_write  =  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_26  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_51  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_29  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_31  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_32  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_33  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_34  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_38  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_39  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_40  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_41  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_42  ; 
   reg  dcache__s1_flush_valid  ; 
   reg  dcache__cached_grant_wait  ; 
   reg  dcache__release_ack_wait  ; 
   reg[31:0]  dcache__release_ack_addr  ; 
   reg[3:0]  dcache__release_state  ; 
   wire  dcache___canAcceptCachedGrant_T  =  dcache__release_state  ==4'h1; 
   wire  dcache___inWriteback_T_1  =  dcache__release_state  ==4'h2; 
   wire  dcache__inWriteback  =  dcache___canAcceptCachedGrant_T  |  dcache___inWriteback_T_1  ; 
   wire  dcache___io_cpu_req_ready_T_4  =  dcache__release_state  ==4'h0&~  dcache__cached_grant_wait  &~  dcache__s1_nack  ; 
   reg  dcache__uncachedInFlight_0  ; 
   reg[33:0]  dcache__uncachedReqs_addr_0  ; 
   reg[5:0]  dcache__uncachedReqs_tag_0  ; 
   reg[1:0]  dcache__uncachedReqs_size_0  ; 
   reg  dcache__uncachedReqs_signed_0  ; 
   wire  dcache___pstore_drain_opportunistic_T  =  dcache__io_cpu_req_bits_cmd  ==5'h0; 
   wire  dcache___pstore_drain_opportunistic_T_1  =  dcache__io_cpu_req_bits_cmd  ==5'h10; 
   wire  dcache___pstore_drain_opportunistic_T_2  =  dcache__io_cpu_req_bits_cmd  ==5'h6; 
   wire  dcache___pstore_drain_opportunistic_T_28  =  dcache__io_cpu_req_bits_cmd  ==5'h7; 
   wire  dcache___pstore_drain_opportunistic_T_30  =  dcache__io_cpu_req_bits_cmd  ==5'h4; 
   wire  dcache___pstore_drain_opportunistic_T_31  =  dcache__io_cpu_req_bits_cmd  ==5'h9; 
   wire  dcache___pstore_drain_opportunistic_T_32  =  dcache__io_cpu_req_bits_cmd  ==5'hA; 
   wire  dcache___pstore_drain_opportunistic_T_33  =  dcache__io_cpu_req_bits_cmd  ==5'hB; 
   wire  dcache___pstore_drain_opportunistic_T_37  =  dcache__io_cpu_req_bits_cmd  ==5'h8; 
   wire  dcache___pstore_drain_opportunistic_T_38  =  dcache__io_cpu_req_bits_cmd  ==5'hC; 
   wire  dcache___pstore_drain_opportunistic_T_39  =  dcache__io_cpu_req_bits_cmd  ==5'hD; 
   wire  dcache___pstore_drain_opportunistic_T_40  =  dcache__io_cpu_req_bits_cmd  ==5'hE; 
   wire  dcache___pstore_drain_opportunistic_T_41  =  dcache__io_cpu_req_bits_cmd  ==5'hF; 
   wire  dcache___pstore_drain_opportunistic_T_25  =  dcache__io_cpu_req_bits_cmd  ==5'h1; 
   wire  dcache___pstore_drain_opportunistic_res_T_1  =  dcache__io_cpu_req_bits_cmd  ==5'h3; 
   wire  dcache___dataArb_io_in_3_valid_res_T_2  =  dcache___pstore_drain_opportunistic_T_25  |  dcache___pstore_drain_opportunistic_res_T_1  ; 
   wire  dcache___pstore_drain_opportunistic_T_50  =  dcache__io_cpu_req_bits_cmd  ==5'h11; 
  assign   dcache__dataArb_io_in_valid_3  =  dcache__io_cpu_req_valid  &~  dcache___dataArb_io_in_3_valid_res_T_2  ; 
  assign   dcache__dataArb_io_in_bits_addr_3  =  dcache__io_cpu_req_bits_addr  [11:0]; 
   wire  dcache___GEN_0  =  dcache__dataArb__grant_T_1  &(  dcache___pstore_drain_opportunistic_T  |  dcache___pstore_drain_opportunistic_T_1  |  dcache___pstore_drain_opportunistic_T_2  |  dcache___pstore_drain_opportunistic_T_28  |  dcache___pstore_drain_opportunistic_T_30  |  dcache___pstore_drain_opportunistic_T_31  |  dcache___pstore_drain_opportunistic_T_32  |  dcache___pstore_drain_opportunistic_T_33  |  dcache___pstore_drain_opportunistic_T_37  |  dcache___pstore_drain_opportunistic_T_38  |  dcache___pstore_drain_opportunistic_T_39  |  dcache___pstore_drain_opportunistic_T_40  |  dcache___pstore_drain_opportunistic_T_41  ); 
   reg  dcache__s1_did_read  ; 
  assign   dcache__metaArb_io_in_bits_idx_7  =  dcache__io_cpu_req_bits_addr  [11:6]; 
  assign   dcache__writeEnable  =  dcache__metaArb_io_out_valid  &  dcache__metaArb_io_out_bits_write  ; 
  assign   dcache__readEnable  =  dcache__metaArb_io_out_valid  &~  dcache__metaArb_io_out_bits_write  ; 
   wire[1:0]  dcache___s1_mask_xwr_T  ={  dcache__s1_vaddr  [0]|(|  dcache__s1_req_size  ),~(  dcache__s1_vaddr  [0])}; 
   wire[3:0]  dcache___s1_mask_xwr_T_1  ={(  dcache__s1_vaddr  [1] ?   dcache___s1_mask_xwr_T  :2'h0)|{2{  dcache__s1_req_size  [1]}},  dcache__s1_vaddr  [1] ? 2'h0:  dcache___s1_mask_xwr_T  }; 
   wire[7:0]  dcache__s1_mask_xwr  ={(  dcache__s1_vaddr  [2] ?   dcache___s1_mask_xwr_T_1  :4'h0)|{4{&  dcache__s1_req_size  }},  dcache__s1_vaddr  [2] ? 4'h0:  dcache___s1_mask_xwr_T_1  }; 
   reg  dcache__s2_valid  ; 
   wire  dcache__s2_valid_no_xcpt  =  dcache__s2_valid  &{  dcache__io_cpu_s2_xcpt_ma_ld_0  ,  dcache__io_cpu_s2_xcpt_ma_st_0  ,  dcache__io_cpu_s2_xcpt_pf_ld_0  ,  dcache__io_cpu_s2_xcpt_pf_st_0  ,  dcache__io_cpu_s2_xcpt_ae_ld_0  ,  dcache__io_cpu_s2_xcpt_ae_st_0  }==6'h0; 
   reg  dcache__s2_probe  ; 
   wire  dcache__releaseInFlight  =  dcache__s1_probe  |  dcache__s2_probe  |(|  dcache__release_state  ); 
   reg  dcache__s2_not_nacked_in_s1  ; 
   wire  dcache__s2_valid_masked  =  dcache__s2_valid_no_xcpt  &  dcache__s2_not_nacked_in_s1  ; 
   reg[5:0]  dcache__s2_req_tag  ; 
   reg[4:0]  dcache__s2_req_cmd  ; 
   reg[1:0]  dcache__s2_req_size  ; 
   reg  dcache__s2_req_signed  ; 
   reg[1:0]  dcache__s2_req_dprv  ; 
   reg  dcache__s2_req_dv  ; 
   reg  dcache__s2_tlb_xcpt_pf_ld  ; 
   reg  dcache__s2_tlb_xcpt_pf_st  ; 
   reg  dcache__s2_tlb_xcpt_ae_ld  ; 
   reg  dcache__s2_tlb_xcpt_ae_st  ; 
   reg  dcache__s2_tlb_xcpt_ma_ld  ; 
   reg  dcache__s2_tlb_xcpt_ma_st  ; 
   reg  dcache__s2_pma_cacheable  ; 
   reg[33:0]  dcache__s2_uncached_resp_addr  ; 
   reg[33:0]  dcache__s2_vaddr_r  ; 
   wire  dcache__s2_lr  =  dcache__s2_req_cmd  ==5'h6; 
   wire  dcache__s2_sc  =  dcache__s2_req_cmd  ==5'h7; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  =  dcache__s2_req_cmd  ==5'h4; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  =  dcache__s2_req_cmd  ==5'h9; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  =  dcache__s2_req_cmd  ==5'hA; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  =  dcache__s2_req_cmd  ==5'hB; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  =  dcache__s2_req_cmd  ==5'h8; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  =  dcache__s2_req_cmd  ==5'hC; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  =  dcache__s2_req_cmd  ==5'hD; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  =  dcache__s2_req_cmd  ==5'hE; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  =  dcache__s2_req_cmd  ==5'hF; 
   wire  dcache__s2_read  =  dcache__s2_req_cmd  ==5'h0|  dcache__s2_req_cmd  ==5'h10|  dcache__s2_lr  |  dcache__s2_sc  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  ; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_23  =  dcache__s2_req_cmd  ==5'h1; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  =  dcache__s2_req_cmd  ==5'h11; 
   wire  dcache__s2_write  =  dcache___metaArb_io_in_3_bits_data_c_cat_T_23  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |  dcache__s2_sc  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  ; 
   wire  dcache__s2_readwrite  =  dcache__s2_read  |  dcache__s2_write  ; 
   reg  dcache__s2_flush_valid  ; 
   reg[21:0]  dcache__s2_meta_corrected_r  ; 
   reg[63:0]  dcache__s2_data  ; 
   reg[1:0]  dcache__s2_probe_state_state  ; 
   reg[1:0]  dcache__s2_hit_state_state  ; 
   wire  dcache___metaArb_io_in_3_bits_data_c_cat_T_46  =  dcache__s2_req_cmd  ==5'h3; 
   wire[3:0]  dcache___GEN_1  ={  dcache___metaArb_io_in_3_bits_data_c_cat_T_23  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |  dcache__s2_sc  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  ,  dcache___metaArb_io_in_3_bits_data_c_cat_T_23  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |  dcache__s2_sc  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_46  |  dcache__s2_lr  ,  dcache__s2_hit_state_state  }; 
   wire  dcache__s2_hit  =  dcache___GEN_1  ==4'h3|  dcache___GEN_1  ==4'h2|  dcache___GEN_1  ==4'h1|  dcache___GEN_1  ==4'h7|  dcache___GEN_1  ==4'h6|(&  dcache___GEN_1  )|  dcache___GEN_1  ==4'hE; 
   reg[1:0]  dcache__casez_tmp  ; 
   wire[1:0]  dcache___GEN_2  ={1'h0,  dcache___GEN_1  ==4'hC}; 
  always @(*)
       begin 
         casez (  dcache___GEN_1  )
          4 'b0000: 
              dcache__casez_tmp   =2'h0;
          4 'b0001: 
              dcache__casez_tmp   =2'h1;
          4 'b0010: 
              dcache__casez_tmp   =2'h2;
          4 'b0011: 
              dcache__casez_tmp   =2'h3;
          4 'b0100: 
              dcache__casez_tmp   =2'h1;
          4 'b0101: 
              dcache__casez_tmp   =2'h2;
          4 'b0110: 
              dcache__casez_tmp   =2'h2;
          4 'b0111: 
              dcache__casez_tmp   =2'h3;
          4 'b1000: 
              dcache__casez_tmp   =  dcache___GEN_2  ;
          4 'b1001: 
              dcache__casez_tmp   =  dcache___GEN_2  ;
          4 'b1010: 
              dcache__casez_tmp   =  dcache___GEN_2  ;
          4 'b1011: 
              dcache__casez_tmp   =  dcache___GEN_2  ;
          4 'b1100: 
              dcache__casez_tmp   =  dcache___GEN_2  ;
          4 'b1101: 
              dcache__casez_tmp   =2'h2;
          4 'b1110: 
              dcache__casez_tmp   =2'h3;
          default : 
              dcache__casez_tmp   =2'h3;
         endcase 
       end
  
   wire  dcache__s2_valid_hit_maybe_flush_pre_data_ecc_and_waw  =  dcache__s2_valid_masked  &  dcache__s2_hit  ; 
   wire  dcache__s2_valid_hit_pre_data_ecc_and_waw  =  dcache__s2_valid_hit_maybe_flush_pre_data_ecc_and_waw  &  dcache__s2_readwrite  ; 
   wire  dcache__s2_valid_flush_line  =  dcache__s2_valid_hit_maybe_flush_pre_data_ecc_and_waw  &  dcache__s2_req_cmd  ==5'h5&  dcache__s2_req_size  [0]; 
   wire  dcache__s2_valid_miss  =  dcache__s2_valid_masked  &  dcache__s2_readwrite  &~  dcache__s2_hit  ; 
   wire  dcache__s2_valid_cached_miss  =  dcache__s2_valid_miss  &  dcache__s2_pma_cacheable  &~  dcache__uncachedInFlight_0  ; 
   wire  dcache__s2_want_victimize  =  dcache__s2_valid_cached_miss  |  dcache__s2_valid_flush_line  |  dcache__s2_flush_valid  ; 
   wire  dcache__s2_valid_uncached_pending  =  dcache__s2_valid_miss  &~  dcache__s2_pma_cacheable  &~  dcache__uncachedInFlight_0  ; 
   wire[1:0]  dcache__s2_victim_state_state  =(|  dcache__s2_hit_state_state  ) ?   dcache__s2_hit_state_state  :  dcache__s2_meta_corrected_r  [21:20]; 
   wire[3:0]  dcache___GEN_3  ={  dcache__probe_bits_param  ,  dcache__s2_probe_state_state  }; 
   wire  dcache___GEN_4  =  dcache___GEN_3  ==4'hB; 
   wire  dcache___GEN_5  =  dcache___GEN_3  ==4'h4; 
   wire  dcache___GEN_6  =  dcache___GEN_3  ==4'h5; 
   wire  dcache___GEN_7  =  dcache___GEN_3  ==4'h6; 
   wire  dcache___GEN_8  =  dcache___GEN_3  ==4'h7; 
   wire  dcache___GEN_9  =  dcache___GEN_3  ==4'h0; 
   wire  dcache___GEN_10  =  dcache___GEN_3  ==4'h1; 
   wire  dcache___GEN_11  =  dcache___GEN_3  ==4'h2; 
   wire  dcache___GEN_12  =  dcache___GEN_3  ==4'h3; 
   wire  dcache__s2_prb_ack_data  =  dcache___GEN_12  |~(  dcache___GEN_11  |  dcache___GEN_10  |  dcache___GEN_9  )&(  dcache___GEN_8  |~(  dcache___GEN_7  |  dcache___GEN_6  |  dcache___GEN_5  )&  dcache___GEN_4  ); 
   wire  dcache___GEN_13  =  dcache___GEN_12  |  dcache___GEN_11  ; 
   wire  dcache__s2_victim_dirty  =&  dcache__s2_victim_state_state  ; 
   wire  dcache__io_cpu_s2_nack_0  =  dcache__s2_valid_no_xcpt  &~(  dcache__s2_valid_uncached_pending  &  dcache__auto_out_a_ready  )&~(  dcache__s2_valid_masked  &  dcache__s2_req_cmd  ==5'h17)&~  dcache__s2_valid_hit_pre_data_ecc_and_waw  ; 
  assign   dcache__metaArb_io_in_valid_2  =  dcache__s2_valid_hit_pre_data_ecc_and_waw  &  dcache__s2_hit_state_state  !=  dcache__casez_tmp  ; 
   wire  dcache___GEN_14  =  dcache__io_cpu_s2_nack_0  |  dcache__metaArb_io_in_valid_2  ; 
  assign   dcache__metaArb_io_in_bits_idx_4  =  dcache__probe_bits_address  [11:6]; 
  assign   dcache__metaArb_io_in_bits_idx_3  =  dcache__s2_req_addr  [11:6]; 
  assign   dcache__metaArb_io_in_bits_data_2  ={  dcache__casez_tmp  ,  dcache__s2_req_addr  [31:12]}; 
   reg[6:0]  dcache__lrscCount  ; 
   reg[27:0]  dcache__lrscAddr  ; 
   wire  dcache__s2_sc_fail  =  dcache__s2_sc  &~((|(  dcache__lrscCount  [6:2]))&  dcache__lrscAddr  ==  dcache__s2_req_addr  [33:6]); 
   reg[4:0]  dcache__pstore1_cmd  ; 
   reg[33:0]  dcache__pstore1_addr  ; 
   reg[63:0]  dcache__pstore1_data  ; 
   reg[7:0]  dcache__pstore1_mask  ; 
   reg  dcache__pstore1_rmw  ; 
   wire  dcache___pstore1_held_T  =  dcache__s2_valid_hit_pre_data_ecc_and_waw  &  dcache__s2_write  ; 
   reg  dcache__pstore2_valid  ; 
   wire  dcache___pstore_drain_opportunistic_res_T_2  =  dcache___pstore_drain_opportunistic_T_25  |  dcache___pstore_drain_opportunistic_res_T_1  ; 
   reg  dcache__pstore_drain_on_miss_REG  ; 
   reg  dcache__pstore1_held  ; 
   wire  dcache__pstore1_valid_likely  =  dcache__s2_valid  &  dcache__s2_write  |  dcache__pstore1_held  ; 
   wire  dcache__pstore1_valid  =  dcache___pstore1_held_T  &~  dcache__s2_sc_fail  |  dcache__pstore1_held  ; 
   wire  dcache__pstore_drain_structural  =  dcache__pstore1_valid_likely  &  dcache__pstore2_valid  &(  dcache__s1_valid  &  dcache__s1_write  |  dcache__pstore1_rmw  ); 
   wire  dcache___dataArb_io_in_0_valid_T_4  =  dcache__s2_valid_hit_pre_data_ecc_and_waw  &  dcache__s2_write  ; 
   wire  dcache___dataArb_io_in_0_valid_T_9  =~(  dcache__io_cpu_req_valid  &~  dcache___pstore_drain_opportunistic_res_T_2  )|  dcache__releaseInFlight  |  dcache__pstore_drain_on_miss_REG  ; 
  assign   dcache__pstore_drain  =  dcache__pstore_drain_structural  |((  dcache___dataArb_io_in_0_valid_T_4  |  dcache__pstore1_held  )&~  dcache__pstore1_rmw  |  dcache__pstore2_valid  )&  dcache___dataArb_io_in_0_valid_T_9  ; 
   reg[33:0]  dcache__pstore2_addr  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r_1  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r_2  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r_3  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r_4  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r_5  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r_6  ; 
   reg[7:0]  dcache__pstore2_storegen_data_r_7  ; 
   reg[7:0]  dcache__pstore2_storegen_mask  ; 
  assign   dcache__dataArb_io_in_valid_0  =  dcache__pstore_drain_structural  |((  dcache___dataArb_io_in_0_valid_T_4  |  dcache__pstore1_held  )&~  dcache__pstore1_rmw  |  dcache__pstore2_valid  )&  dcache___dataArb_io_in_0_valid_T_9  ; 
  assign   dcache___dataArb_io_in_0_bits_wordMask_wordMask_T  =  dcache__pstore2_valid   ?   dcache__pstore2_addr  [11:0]:  dcache__pstore1_addr  [11:0]; 
  assign   dcache__dataArb_io_in_bits_wdata_0  =  dcache__pstore2_valid   ? {  dcache__pstore2_storegen_data_r_7  ,  dcache__pstore2_storegen_data_r_6  ,  dcache__pstore2_storegen_data_r_5  ,  dcache__pstore2_storegen_data_r_4  ,  dcache__pstore2_storegen_data_r_3  ,  dcache__pstore2_storegen_data_r_2  ,  dcache__pstore2_storegen_data_r_1  ,  dcache__pstore2_storegen_data_r  }:  dcache__pstore1_data  ; 
  assign   dcache__dataArb_io_in_bits_eccMask_0  =  dcache__pstore2_valid   ?   dcache__pstore2_storegen_mask  :  dcache__pstore1_mask  ; 
   wire  dcache___GEN_15  =  dcache__s1_valid  &  dcache__s1_read  &(  dcache__pstore1_valid_likely  &  dcache__pstore1_addr  [11:3]==  dcache__s1_vaddr  [11:3]&(  dcache__s1_write   ? (|(  dcache__pstore1_mask  &  dcache__s1_mask_xwr  )):(|(  dcache__pstore1_mask  &  dcache__s1_mask_xwr  )))|  dcache__pstore2_valid  &  dcache__pstore2_addr  [11:3]==  dcache__s1_vaddr  [11:3]&(  dcache__s1_write   ? (|(  dcache__pstore2_storegen_mask  &  dcache__s1_mask_xwr  )):(|(  dcache__pstore2_storegen_mask  &  dcache__s1_mask_xwr  )))); 
   wire  dcache__get_a_mask_size  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__get_a_mask_acc  =(&  dcache__s2_req_size  )|  dcache__get_a_mask_size  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__get_a_mask_acc_1  =(&  dcache__s2_req_size  )|  dcache__get_a_mask_size  &  dcache__s2_req_addr  [2]; 
   wire  dcache__get_a_mask_size_1  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__get_a_mask_eq_2  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__get_a_mask_acc_2  =  dcache__get_a_mask_acc  |  dcache__get_a_mask_size_1  &  dcache__get_a_mask_eq_2  ; 
   wire  dcache__get_a_mask_eq_3  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__get_a_mask_acc_3  =  dcache__get_a_mask_acc  |  dcache__get_a_mask_size_1  &  dcache__get_a_mask_eq_3  ; 
   wire  dcache__get_a_mask_eq_4  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__get_a_mask_acc_4  =  dcache__get_a_mask_acc_1  |  dcache__get_a_mask_size_1  &  dcache__get_a_mask_eq_4  ; 
   wire  dcache__get_a_mask_eq_5  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__get_a_mask_acc_5  =  dcache__get_a_mask_acc_1  |  dcache__get_a_mask_size_1  &  dcache__get_a_mask_eq_5  ; 
   wire  dcache__put_a_mask_size  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__put_a_mask_acc  =(&  dcache__s2_req_size  )|  dcache__put_a_mask_size  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__put_a_mask_acc_1  =(&  dcache__s2_req_size  )|  dcache__put_a_mask_size  &  dcache__s2_req_addr  [2]; 
   wire  dcache__put_a_mask_size_1  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__put_a_mask_eq_2  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__put_a_mask_acc_2  =  dcache__put_a_mask_acc  |  dcache__put_a_mask_size_1  &  dcache__put_a_mask_eq_2  ; 
   wire  dcache__put_a_mask_eq_3  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__put_a_mask_acc_3  =  dcache__put_a_mask_acc  |  dcache__put_a_mask_size_1  &  dcache__put_a_mask_eq_3  ; 
   wire  dcache__put_a_mask_eq_4  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__put_a_mask_acc_4  =  dcache__put_a_mask_acc_1  |  dcache__put_a_mask_size_1  &  dcache__put_a_mask_eq_4  ; 
   wire  dcache__put_a_mask_eq_5  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__put_a_mask_acc_5  =  dcache__put_a_mask_acc_1  |  dcache__put_a_mask_size_1  &  dcache__put_a_mask_eq_5  ; 
   wire  dcache__atomics_a_mask_size  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_1  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_1  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_2  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_2  =  dcache__atomics_a_mask_acc  |  dcache__atomics_a_mask_size_1  &  dcache__atomics_a_mask_eq_2  ; 
   wire  dcache__atomics_a_mask_eq_3  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_3  =  dcache__atomics_a_mask_acc  |  dcache__atomics_a_mask_size_1  &  dcache__atomics_a_mask_eq_3  ; 
   wire  dcache__atomics_a_mask_eq_4  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_4  =  dcache__atomics_a_mask_acc_1  |  dcache__atomics_a_mask_size_1  &  dcache__atomics_a_mask_eq_4  ; 
   wire  dcache__atomics_a_mask_eq_5  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_5  =  dcache__atomics_a_mask_acc_1  |  dcache__atomics_a_mask_size_1  &  dcache__atomics_a_mask_eq_5  ; 
   wire  dcache__atomics_a_mask_size_3  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_14  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_3  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_15  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_3  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_4  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_16  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_16  =  dcache__atomics_a_mask_acc_14  |  dcache__atomics_a_mask_size_4  &  dcache__atomics_a_mask_eq_16  ; 
   wire  dcache__atomics_a_mask_eq_17  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_17  =  dcache__atomics_a_mask_acc_14  |  dcache__atomics_a_mask_size_4  &  dcache__atomics_a_mask_eq_17  ; 
   wire  dcache__atomics_a_mask_eq_18  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_18  =  dcache__atomics_a_mask_acc_15  |  dcache__atomics_a_mask_size_4  &  dcache__atomics_a_mask_eq_18  ; 
   wire  dcache__atomics_a_mask_eq_19  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_19  =  dcache__atomics_a_mask_acc_15  |  dcache__atomics_a_mask_size_4  &  dcache__atomics_a_mask_eq_19  ; 
   wire  dcache__atomics_a_mask_size_6  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_28  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_6  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_29  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_6  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_7  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_30  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_30  =  dcache__atomics_a_mask_acc_28  |  dcache__atomics_a_mask_size_7  &  dcache__atomics_a_mask_eq_30  ; 
   wire  dcache__atomics_a_mask_eq_31  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_31  =  dcache__atomics_a_mask_acc_28  |  dcache__atomics_a_mask_size_7  &  dcache__atomics_a_mask_eq_31  ; 
   wire  dcache__atomics_a_mask_eq_32  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_32  =  dcache__atomics_a_mask_acc_29  |  dcache__atomics_a_mask_size_7  &  dcache__atomics_a_mask_eq_32  ; 
   wire  dcache__atomics_a_mask_eq_33  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_33  =  dcache__atomics_a_mask_acc_29  |  dcache__atomics_a_mask_size_7  &  dcache__atomics_a_mask_eq_33  ; 
   wire  dcache__atomics_a_mask_size_9  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_42  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_9  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_43  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_9  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_10  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_44  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_44  =  dcache__atomics_a_mask_acc_42  |  dcache__atomics_a_mask_size_10  &  dcache__atomics_a_mask_eq_44  ; 
   wire  dcache__atomics_a_mask_eq_45  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_45  =  dcache__atomics_a_mask_acc_42  |  dcache__atomics_a_mask_size_10  &  dcache__atomics_a_mask_eq_45  ; 
   wire  dcache__atomics_a_mask_eq_46  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_46  =  dcache__atomics_a_mask_acc_43  |  dcache__atomics_a_mask_size_10  &  dcache__atomics_a_mask_eq_46  ; 
   wire  dcache__atomics_a_mask_eq_47  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_47  =  dcache__atomics_a_mask_acc_43  |  dcache__atomics_a_mask_size_10  &  dcache__atomics_a_mask_eq_47  ; 
   wire  dcache__atomics_a_mask_size_12  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_56  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_12  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_57  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_12  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_13  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_58  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_58  =  dcache__atomics_a_mask_acc_56  |  dcache__atomics_a_mask_size_13  &  dcache__atomics_a_mask_eq_58  ; 
   wire  dcache__atomics_a_mask_eq_59  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_59  =  dcache__atomics_a_mask_acc_56  |  dcache__atomics_a_mask_size_13  &  dcache__atomics_a_mask_eq_59  ; 
   wire  dcache__atomics_a_mask_eq_60  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_60  =  dcache__atomics_a_mask_acc_57  |  dcache__atomics_a_mask_size_13  &  dcache__atomics_a_mask_eq_60  ; 
   wire  dcache__atomics_a_mask_eq_61  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_61  =  dcache__atomics_a_mask_acc_57  |  dcache__atomics_a_mask_size_13  &  dcache__atomics_a_mask_eq_61  ; 
   wire  dcache__atomics_a_mask_size_15  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_70  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_15  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_71  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_15  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_16  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_72  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_72  =  dcache__atomics_a_mask_acc_70  |  dcache__atomics_a_mask_size_16  &  dcache__atomics_a_mask_eq_72  ; 
   wire  dcache__atomics_a_mask_eq_73  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_73  =  dcache__atomics_a_mask_acc_70  |  dcache__atomics_a_mask_size_16  &  dcache__atomics_a_mask_eq_73  ; 
   wire  dcache__atomics_a_mask_eq_74  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_74  =  dcache__atomics_a_mask_acc_71  |  dcache__atomics_a_mask_size_16  &  dcache__atomics_a_mask_eq_74  ; 
   wire  dcache__atomics_a_mask_eq_75  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_75  =  dcache__atomics_a_mask_acc_71  |  dcache__atomics_a_mask_size_16  &  dcache__atomics_a_mask_eq_75  ; 
   wire  dcache__atomics_a_mask_size_18  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_84  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_18  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_85  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_18  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_19  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_86  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_86  =  dcache__atomics_a_mask_acc_84  |  dcache__atomics_a_mask_size_19  &  dcache__atomics_a_mask_eq_86  ; 
   wire  dcache__atomics_a_mask_eq_87  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_87  =  dcache__atomics_a_mask_acc_84  |  dcache__atomics_a_mask_size_19  &  dcache__atomics_a_mask_eq_87  ; 
   wire  dcache__atomics_a_mask_eq_88  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_88  =  dcache__atomics_a_mask_acc_85  |  dcache__atomics_a_mask_size_19  &  dcache__atomics_a_mask_eq_88  ; 
   wire  dcache__atomics_a_mask_eq_89  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_89  =  dcache__atomics_a_mask_acc_85  |  dcache__atomics_a_mask_size_19  &  dcache__atomics_a_mask_eq_89  ; 
   wire  dcache__atomics_a_mask_size_21  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_98  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_21  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_99  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_21  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_22  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_100  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_100  =  dcache__atomics_a_mask_acc_98  |  dcache__atomics_a_mask_size_22  &  dcache__atomics_a_mask_eq_100  ; 
   wire  dcache__atomics_a_mask_eq_101  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_101  =  dcache__atomics_a_mask_acc_98  |  dcache__atomics_a_mask_size_22  &  dcache__atomics_a_mask_eq_101  ; 
   wire  dcache__atomics_a_mask_eq_102  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_102  =  dcache__atomics_a_mask_acc_99  |  dcache__atomics_a_mask_size_22  &  dcache__atomics_a_mask_eq_102  ; 
   wire  dcache__atomics_a_mask_eq_103  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_103  =  dcache__atomics_a_mask_acc_99  |  dcache__atomics_a_mask_size_22  &  dcache__atomics_a_mask_eq_103  ; 
   wire  dcache__atomics_a_mask_size_24  =  dcache__s2_req_size  ==2'h2; 
   wire  dcache__atomics_a_mask_acc_112  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_24  &~(  dcache__s2_req_addr  [2]); 
   wire  dcache__atomics_a_mask_acc_113  =(&  dcache__s2_req_size  )|  dcache__atomics_a_mask_size_24  &  dcache__s2_req_addr  [2]; 
   wire  dcache__atomics_a_mask_size_25  =  dcache__s2_req_size  ==2'h1; 
   wire  dcache__atomics_a_mask_eq_114  =~(  dcache__s2_req_addr  [2])&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_114  =  dcache__atomics_a_mask_acc_112  |  dcache__atomics_a_mask_size_25  &  dcache__atomics_a_mask_eq_114  ; 
   wire  dcache__atomics_a_mask_eq_115  =~(  dcache__s2_req_addr  [2])&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_115  =  dcache__atomics_a_mask_acc_112  |  dcache__atomics_a_mask_size_25  &  dcache__atomics_a_mask_eq_115  ; 
   wire  dcache__atomics_a_mask_eq_116  =  dcache__s2_req_addr  [2]&~(  dcache__s2_req_addr  [1]); 
   wire  dcache__atomics_a_mask_acc_116  =  dcache__atomics_a_mask_acc_113  |  dcache__atomics_a_mask_size_25  &  dcache__atomics_a_mask_eq_116  ; 
   wire  dcache__atomics_a_mask_eq_117  =  dcache__s2_req_addr  [2]&  dcache__s2_req_addr  [1]; 
   wire  dcache__atomics_a_mask_acc_117  =  dcache__atomics_a_mask_acc_113  |  dcache__atomics_a_mask_size_25  &  dcache__atomics_a_mask_eq_117  ; 
   wire[7:0]  dcache__atomics_mask  =  dcache___metaArb_io_in_3_bits_data_c_cat_T_39   ? {  dcache__atomics_a_mask_acc_117  |  dcache__atomics_a_mask_eq_117  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_117  |  dcache__atomics_a_mask_eq_117  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_116  |  dcache__atomics_a_mask_eq_116  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_116  |  dcache__atomics_a_mask_eq_116  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_115  |  dcache__atomics_a_mask_eq_115  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_115  |  dcache__atomics_a_mask_eq_115  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_114  |  dcache__atomics_a_mask_eq_114  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_114  |  dcache__atomics_a_mask_eq_114  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_38   ? {  dcache__atomics_a_mask_acc_103  |  dcache__atomics_a_mask_eq_103  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_103  |  dcache__atomics_a_mask_eq_103  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_102  |  dcache__atomics_a_mask_eq_102  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_102  |  dcache__atomics_a_mask_eq_102  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_101  |  dcache__atomics_a_mask_eq_101  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_101  |  dcache__atomics_a_mask_eq_101  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_100  |  dcache__atomics_a_mask_eq_100  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_100  |  dcache__atomics_a_mask_eq_100  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_37   ? {  dcache__atomics_a_mask_acc_89  |  dcache__atomics_a_mask_eq_89  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_89  |  dcache__atomics_a_mask_eq_89  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_88  |  dcache__atomics_a_mask_eq_88  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_88  |  dcache__atomics_a_mask_eq_88  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_87  |  dcache__atomics_a_mask_eq_87  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_87  |  dcache__atomics_a_mask_eq_87  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_86  |  dcache__atomics_a_mask_eq_86  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_86  |  dcache__atomics_a_mask_eq_86  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_36   ? {  dcache__atomics_a_mask_acc_75  |  dcache__atomics_a_mask_eq_75  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_75  |  dcache__atomics_a_mask_eq_75  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_74  |  dcache__atomics_a_mask_eq_74  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_74  |  dcache__atomics_a_mask_eq_74  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_73  |  dcache__atomics_a_mask_eq_73  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_73  |  dcache__atomics_a_mask_eq_73  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_72  |  dcache__atomics_a_mask_eq_72  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_72  |  dcache__atomics_a_mask_eq_72  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_35   ? {  dcache__atomics_a_mask_acc_61  |  dcache__atomics_a_mask_eq_61  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_61  |  dcache__atomics_a_mask_eq_61  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_60  |  dcache__atomics_a_mask_eq_60  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_60  |  dcache__atomics_a_mask_eq_60  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_59  |  dcache__atomics_a_mask_eq_59  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_59  |  dcache__atomics_a_mask_eq_59  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_58  |  dcache__atomics_a_mask_eq_58  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_58  |  dcache__atomics_a_mask_eq_58  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_31   ? {  dcache__atomics_a_mask_acc_47  |  dcache__atomics_a_mask_eq_47  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_47  |  dcache__atomics_a_mask_eq_47  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_46  |  dcache__atomics_a_mask_eq_46  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_46  |  dcache__atomics_a_mask_eq_46  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_45  |  dcache__atomics_a_mask_eq_45  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_45  |  dcache__atomics_a_mask_eq_45  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_44  |  dcache__atomics_a_mask_eq_44  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_44  |  dcache__atomics_a_mask_eq_44  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_30   ? {  dcache__atomics_a_mask_acc_33  |  dcache__atomics_a_mask_eq_33  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_33  |  dcache__atomics_a_mask_eq_33  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_32  |  dcache__atomics_a_mask_eq_32  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_32  |  dcache__atomics_a_mask_eq_32  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_31  |  dcache__atomics_a_mask_eq_31  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_31  |  dcache__atomics_a_mask_eq_31  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_30  |  dcache__atomics_a_mask_eq_30  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_30  |  dcache__atomics_a_mask_eq_30  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_29   ? {  dcache__atomics_a_mask_acc_19  |  dcache__atomics_a_mask_eq_19  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_19  |  dcache__atomics_a_mask_eq_19  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_18  |  dcache__atomics_a_mask_eq_18  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_18  |  dcache__atomics_a_mask_eq_18  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_17  |  dcache__atomics_a_mask_eq_17  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_17  |  dcache__atomics_a_mask_eq_17  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_16  |  dcache__atomics_a_mask_eq_16  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_16  |  dcache__atomics_a_mask_eq_16  &~(  dcache__s2_req_addr  [0])}:  dcache___metaArb_io_in_3_bits_data_c_cat_T_28   ? {  dcache__atomics_a_mask_acc_5  |  dcache__atomics_a_mask_eq_5  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_5  |  dcache__atomics_a_mask_eq_5  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_4  |  dcache__atomics_a_mask_eq_4  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_4  |  dcache__atomics_a_mask_eq_4  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_3  |  dcache__atomics_a_mask_eq_3  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_3  |  dcache__atomics_a_mask_eq_3  &~(  dcache__s2_req_addr  [0]),  dcache__atomics_a_mask_acc_2  |  dcache__atomics_a_mask_eq_2  &  dcache__s2_req_addr  [0],  dcache__atomics_a_mask_acc_2  |  dcache__atomics_a_mask_eq_2  &~(  dcache__s2_req_addr  [0])}:8'h0; 
   wire  dcache__tl_out_a_valid  =  dcache__s2_valid_uncached_pending  |  dcache__s2_valid_cached_miss  &~(  dcache__release_ack_wait  &(  dcache__s2_req_addr  [20:6]^  dcache__release_ack_addr  [20:6])==15'h0)&~  dcache__s2_victim_dirty  ; 
   wire  dcache___GEN_16  =~  dcache__s2_write  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |~  dcache__s2_read  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  ; 
   wire  dcache___io_errors_bus_valid_T  =  dcache__nodeOut_d_ready  &  dcache__auto_out_d_valid  ; 
   wire[26:0]  dcache___beats1_decode_T_1  =27'hFFF<<  dcache__auto_out_d_bits_size  ; 
   wire[8:0]  dcache__beats1  =  dcache__auto_out_d_bits_opcode  [0] ? ~(  dcache___beats1_decode_T_1  [11:3]):9'h0; 
   reg[8:0]  dcache__counter  ; 
   wire[8:0]  dcache___counter1_T  =  dcache__counter  -9'h1; 
   wire  dcache__d_last  =  dcache__counter  ==9'h1|  dcache__beats1  ==9'h0; 
   wire[8:0]  dcache__count  =  dcache__beats1  &~  dcache___counter1_T  ; 
   wire  dcache__grantIsUncachedData  =  dcache__auto_out_d_bits_opcode  ==3'h1; 
   wire  dcache__grantIsUncached  =  dcache__grantIsUncachedData  |  dcache__auto_out_d_bits_opcode  ==3'h0|  dcache__auto_out_d_bits_opcode  ==3'h2; 
   wire  dcache__grantIsRefill  =  dcache__auto_out_d_bits_opcode  ==3'h5; 
   wire  dcache__grantIsCached  =  dcache__auto_out_d_bits_opcode  ==3'h4|  dcache__grantIsRefill  ; 
   wire  dcache__grantIsVoluntary  =  dcache__auto_out_d_bits_opcode  ==3'h6; 
   reg  dcache__grantInProgress  ; 
   reg[2:0]  dcache__blockProbeAfterGrantCount  ; 
   wire  dcache___metaArb_io_in_4_valid_T  =  dcache__release_state  ==4'h6; 
   wire  dcache___nodeOut_c_valid_T_1  =  dcache__release_state  ==4'h9; 
   wire  dcache___canAcceptCachedGrant_T_4  =  dcache___canAcceptCachedGrant_T  |  dcache___metaArb_io_in_4_valid_T  |  dcache___nodeOut_c_valid_T_1  ; 
   wire  dcache___GEN_17  =  dcache___io_errors_bus_valid_T  &  dcache__grantIsCached  ; 
   wire  dcache___GEN_18  =  dcache__auto_out_d_bits_source  &  dcache__d_last  ; 
   wire  dcache___GEN_19  =~  dcache___io_errors_bus_valid_T  |  dcache__grantIsCached  |~(  dcache__grantIsUncached  &  dcache__grantIsUncachedData  ); 
   wire  dcache___GEN_20  =  dcache__grantIsRefill  &  dcache__dataArb_io_in_valid_0  ; 
   wire  dcache__nodeOut_e_valid  =~  dcache___GEN_20  &  dcache__auto_out_d_valid  &~(|  dcache__counter  )&  dcache__grantIsCached  &~  dcache___canAcceptCachedGrant_T_4  ; 
  assign   dcache__dataArb_io_in_bits_addr_1  ={  dcache__s2_req_addr  [11:6]|  dcache__count  [8:3],  dcache__count  [2:0],3'h0}; 
  assign   dcache__metaArb_io_in_valid_3  =  dcache__grantIsCached  &  dcache__d_last  &  dcache___io_errors_bus_valid_T  &~  dcache__auto_out_d_bits_denied  ; 
   wire[3:0]  dcache___metaArb_io_in_3_bits_data_T_1  ={  dcache___metaArb_io_in_3_bits_data_c_cat_T_23  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |  dcache__s2_sc  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  ,  dcache___metaArb_io_in_3_bits_data_c_cat_T_23  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |  dcache__s2_sc  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_46  |  dcache__s2_lr  ,  dcache__auto_out_d_bits_param  }; 
  assign   dcache__metaArb_io_in_bits_data_3  ={  dcache___metaArb_io_in_3_bits_data_T_1  ==4'hC ? 2'h3:  dcache___metaArb_io_in_3_bits_data_T_1  ==4'h4|  dcache___metaArb_io_in_3_bits_data_T_1  ==4'h0 ? 2'h2:{1'h0,  dcache___metaArb_io_in_3_bits_data_T_1  ==4'h1},  dcache__s2_req_addr  [31:12]}; 
   reg  dcache__blockUncachedGrant  ; 
   wire  dcache___GEN_21  =  dcache__grantIsUncachedData  &(  dcache__blockUncachedGrant  |  dcache__s1_valid  ); 
  assign   dcache__nodeOut_d_ready  =~(  dcache___GEN_21  |  dcache___GEN_20  )&(~  dcache__grantIsCached  |((|  dcache__counter  )|  dcache__auto_out_e_ready  )&~  dcache___canAcceptCachedGrant_T_4  ); 
   wire  dcache__io_cpu_req_ready_0  =  dcache___GEN_21   ? ~(  dcache__auto_out_d_valid  |  dcache__metaArb__grant_T_5  |  dcache___GEN_0  )&  dcache___io_cpu_req_ready_T_4  :~(  dcache__metaArb__grant_T_5  |  dcache___GEN_0  )&  dcache___io_cpu_req_ready_T_4  ; 
   wire  dcache___GEN_22  =  dcache___GEN_21  &  dcache__auto_out_d_valid  ; 
  assign   dcache__dataArb_io_in_valid_1  =  dcache___GEN_22  |  dcache__auto_out_d_valid  &  dcache__grantIsRefill  &~  dcache___canAcceptCachedGrant_T_4  ; 
  assign   dcache__dataArb_io_in_bits_write_1  =~  dcache___GEN_21  |~  dcache__auto_out_d_valid  ; 
   wire  dcache__block_probe_for_core_progress  =(|  dcache__blockProbeAfterGrantCount  )|(|(  dcache__lrscCount  [6:2])); 
   wire  dcache__nodeOut_b_ready  =~  dcache__metaArb__grant_T_3  &~(  dcache__block_probe_for_core_progress  |  dcache__releaseInFlight  |  dcache__release_ack_wait  &(  dcache__auto_out_b_bits_address  [20:6]^  dcache__release_ack_addr  [20:6])==15'h0|  dcache__grantInProgress  |  dcache__s1_valid  |  dcache__s2_valid  ); 
   wire  dcache___io_cpu_perf_release_T  =  dcache__auto_out_c_ready  &  dcache__nodeOut_c_valid  ; 
   wire[26:0]  dcache___GEN_23  ={23'h0,  dcache__nodeOut_c_bits_size  }; 
   wire[26:0]  dcache___beats1_decode_T_5  =27'hFFF<<  dcache___GEN_23  ; 
   wire[8:0]  dcache__beats1_1  =  dcache__nodeOut_c_bits_opcode  [0] ? ~(  dcache___beats1_decode_T_5  [11:3]):9'h0; 
   reg[8:0]  dcache__counter_1  ; 
   wire[8:0]  dcache___counter1_T_1  =  dcache__counter_1  -9'h1; 
   wire  dcache__c_first  =  dcache__counter_1  ==9'h0; 
   wire  dcache__releaseDone  =(  dcache__counter_1  ==9'h1|  dcache__beats1_1  ==9'h0)&  dcache___io_cpu_perf_release_T  ; 
   reg  dcache__s1_release_data_valid  ; 
   reg  dcache__s2_release_data_valid  ; 
   wire  dcache__releaseRejected  =  dcache__s2_release_data_valid  &~  dcache___io_cpu_perf_release_T  ; 
   wire[9:0]  dcache___releaseDataBeat_T_5  ={1'h0,  dcache__beats1_1  &~  dcache___counter1_T_1  }+{8'h0,  dcache__releaseRejected   ? 2'h0:{1'h0,  dcache__s1_release_data_valid  }+{1'h0,  dcache__s2_release_data_valid  }}; 
  assign   dcache__s1_nack  =  dcache__s2_probe   ?   dcache__s2_prb_ack_data  |(|  dcache__s2_probe_state_state  )|~  dcache__releaseDone  |  dcache___GEN_15  |  dcache___GEN_14  :  dcache___GEN_15  |  dcache___GEN_14  ; 
   wire  dcache___GEN_24  =  dcache__release_state  ==4'h4; 
  assign   dcache__metaArb_io_in_valid_6  =  dcache___GEN_24  |  dcache__auto_out_b_valid  &(~  dcache__block_probe_for_core_progress  |(|  dcache__lrscCount  )&~(|(  dcache__lrscCount  [6:2]))); 
  assign   dcache__metaArb_io_in_bits_idx_6  =  dcache___GEN_24   ?   dcache__metaArb_io_in_bits_idx_4  :  dcache__auto_out_b_bits_address  [11:6]; 
   wire  dcache___GEN_25  =  dcache__release_state  ==4'h5; 
   wire  dcache___GEN_26  =  dcache__release_state  ==4'h3; 
  assign   dcache__nodeOut_c_valid  =  dcache___GEN_26  |  dcache___GEN_25  |  dcache__s2_probe  &~  dcache__s2_prb_ack_data  |  dcache__s2_release_data_valid  &~(  dcache__c_first  &  dcache__release_ack_wait  ); 
   wire  dcache___GEN_27  =  dcache___canAcceptCachedGrant_T  |  dcache___metaArb_io_in_4_valid_T  |  dcache___nodeOut_c_valid_T_1  ; 
  assign   dcache__nodeOut_c_bits_opcode  =  dcache___GEN_27   ? {2'h3,~  dcache___nodeOut_c_valid_T_1  }:{2'h2,  dcache___inWriteback_T_1  }; 
  assign   dcache__nodeOut_c_bits_size  =  dcache___GEN_27   ? 4'h6:  dcache__probe_bits_size  ; 
  assign   dcache__dataArb_io_in_valid_2  =  dcache__inWriteback  &  dcache___releaseDataBeat_T_5  <10'h8; 
  assign   dcache__dataArb_io_in_bits_addr_2  ={  dcache__metaArb_io_in_bits_idx_4  ,  dcache___releaseDataBeat_T_5  [2:0],3'h0}; 
  assign   dcache__metaArb_io_in_valid_4  =  dcache___metaArb_io_in_4_valid_T  |  dcache__release_state  ==4'h7; 
  assign   dcache__metaArb_io_in_bits_data_7  ={  dcache___GEN_27   ? 2'h0:  dcache___GEN_13   ? 2'h2:  dcache___GEN_10   ? 2'h1:  dcache___GEN_9   ? 2'h0:{1'h0,  dcache___GEN_8  |  dcache___GEN_7  |  dcache___GEN_6  },  dcache__probe_bits_address  [31:12]}; 
   reg  dcache__io_cpu_s2_xcpt_REG  ; 
  assign   dcache__io_cpu_s2_xcpt_pf_ld_0  =  dcache__io_cpu_s2_xcpt_REG  &  dcache__s2_tlb_xcpt_pf_ld  ; 
  assign   dcache__io_cpu_s2_xcpt_pf_st_0  =  dcache__io_cpu_s2_xcpt_REG  &  dcache__s2_tlb_xcpt_pf_st  ; 
  assign   dcache__io_cpu_s2_xcpt_ae_ld_0  =  dcache__io_cpu_s2_xcpt_REG  &  dcache__s2_tlb_xcpt_ae_ld  ; 
  assign   dcache__io_cpu_s2_xcpt_ae_st_0  =  dcache__io_cpu_s2_xcpt_REG  &  dcache__s2_tlb_xcpt_ae_st  ; 
  assign   dcache__io_cpu_s2_xcpt_ma_ld_0  =  dcache__io_cpu_s2_xcpt_REG  &  dcache__s2_tlb_xcpt_ma_ld  ; 
  assign   dcache__io_cpu_s2_xcpt_ma_st_0  =  dcache__io_cpu_s2_xcpt_REG  &  dcache__s2_tlb_xcpt_ma_st  ; 
   reg  dcache__doUncachedResp  ; 
   wire  dcache__io_cpu_replay_next_0  =  dcache___io_errors_bus_valid_T  &  dcache__grantIsUncachedData  ; 
   wire  dcache___GEN_28  =  dcache___io_errors_bus_valid_T  &~  dcache__grantIsCached  ; 
  always @( posedge   dcache__clock  )
       begin 
         if (~  dcache__reset  &~(~(  dcache___pstore_drain_opportunistic_T  |  dcache___pstore_drain_opportunistic_T_1  |  dcache___pstore_drain_opportunistic_T_2  |  dcache___pstore_drain_opportunistic_T_28  |  dcache___pstore_drain_opportunistic_T_30  |  dcache___pstore_drain_opportunistic_T_31  |  dcache___pstore_drain_opportunistic_T_32  |  dcache___pstore_drain_opportunistic_T_33  |  dcache___pstore_drain_opportunistic_T_37  |  dcache___pstore_drain_opportunistic_T_38  |  dcache___pstore_drain_opportunistic_T_39  |  dcache___pstore_drain_opportunistic_T_40  |  dcache___pstore_drain_opportunistic_T_41  |(  dcache___pstore_drain_opportunistic_T_25  |  dcache___pstore_drain_opportunistic_T_50  |  dcache___pstore_drain_opportunistic_T_28  |  dcache___pstore_drain_opportunistic_T_30  |  dcache___pstore_drain_opportunistic_T_31  |  dcache___pstore_drain_opportunistic_T_32  |  dcache___pstore_drain_opportunistic_T_33  |  dcache___pstore_drain_opportunistic_T_37  |  dcache___pstore_drain_opportunistic_T_38  |  dcache___pstore_drain_opportunistic_T_39  |  dcache___pstore_drain_opportunistic_T_40  |  dcache___pstore_drain_opportunistic_T_41  )&  dcache___pstore_drain_opportunistic_T_50  )|~  dcache___dataArb_io_in_3_valid_res_T_2  ))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
              if (1)$display("");
            end 
         if (~  dcache__reset  &~(~(  dcache__s1_valid_masked  &  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_51  )|(&(  dcache__s1_mask_xwr  |~  dcache__io_cpu_s1_data_mask  ))))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:306 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n");
              if (1)$display("");
            end 
         if (~  dcache__reset  &~(~(  dcache___pstore_drain_opportunistic_T  |  dcache___pstore_drain_opportunistic_T_1  |  dcache___pstore_drain_opportunistic_T_2  |  dcache___pstore_drain_opportunistic_T_28  |  dcache___pstore_drain_opportunistic_T_30  |  dcache___pstore_drain_opportunistic_T_31  |  dcache___pstore_drain_opportunistic_T_32  |  dcache___pstore_drain_opportunistic_T_33  |  dcache___pstore_drain_opportunistic_T_37  |  dcache___pstore_drain_opportunistic_T_38  |  dcache___pstore_drain_opportunistic_T_39  |  dcache___pstore_drain_opportunistic_T_40  |  dcache___pstore_drain_opportunistic_T_41  |(  dcache___pstore_drain_opportunistic_T_25  |  dcache___pstore_drain_opportunistic_T_50  |  dcache___pstore_drain_opportunistic_T_28  |  dcache___pstore_drain_opportunistic_T_30  |  dcache___pstore_drain_opportunistic_T_31  |  dcache___pstore_drain_opportunistic_T_32  |  dcache___pstore_drain_opportunistic_T_33  |  dcache___pstore_drain_opportunistic_T_37  |  dcache___pstore_drain_opportunistic_T_38  |  dcache___pstore_drain_opportunistic_T_39  |  dcache___pstore_drain_opportunistic_T_40  |  dcache___pstore_drain_opportunistic_T_41  )&  dcache___pstore_drain_opportunistic_T_50  )|~  dcache___pstore_drain_opportunistic_res_T_2  ))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
              if (1)$display("");
            end 
         if (~  dcache__reset  &~(  dcache__pstore1_rmw  |(  dcache___dataArb_io_in_0_valid_T_4  |  dcache__pstore1_held  )==  dcache__pstore1_valid  ))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:487 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n");
              if (1)$display("");
            end 
         if (  dcache___GEN_17  &~  dcache__reset  &~  dcache__cached_grant_wait  )
            begin 
              if (1)$display("Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:654 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n");
              if (1)$display("");
            end 
         if (  dcache___GEN_28  &  dcache__grantIsUncached  &  dcache___GEN_18  &~  dcache__reset  &~  dcache__uncachedInFlight_0  )
            begin 
              if (1)$display("Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:664 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n");
              if (1)$display("");
            end 
         if (  dcache___GEN_28  &~  dcache__grantIsUncached  &  dcache__grantIsVoluntary  &~  dcache__reset  &~  dcache__release_ack_wait  )
            begin 
              if (1)$display("Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:685 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n");
              if (1)$display("");
            end 
         if (~  dcache__reset  &(  dcache__auto_out_e_ready  &  dcache__nodeOut_e_valid  )!=(  dcache___io_errors_bus_valid_T  &~(|  dcache__counter  )&  dcache__grantIsCached  ))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:693 assert(tl_out.e.fire === (tl_out.d.fire && d_first && grantIsCached))\n");
              if (1)$display("");
            end 
         if (  dcache__s2_want_victimize  &~  dcache__reset  &~(  dcache__s2_valid_flush_line  |  dcache__s2_flush_valid  |  dcache__io_cpu_s2_nack_0  ))
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:794 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n");
              if (1)$display("");
            end 
         if (  dcache__doUncachedResp  &~  dcache__reset  &  dcache__s2_valid_hit_pre_data_ecc_and_waw  )
            begin 
              if (1)$display("Assertion failed\n    at DCache.scala:928 assert(!s2_valid_hit)\n");
              if (1)$display("");
            end 
       end
  
   wire[31:0]  dcache__io_cpu_resp_bits_data_zeroed  =  dcache__s2_req_addr  [2] ?   dcache__s2_data  [63:32]:  dcache__s2_data  [31:0]; 
   wire  dcache___io_cpu_resp_bits_data_word_bypass_T_1  =  dcache__s2_req_size  ==2'h2; 
   wire[15:0]  dcache__io_cpu_resp_bits_data_zeroed_1  =  dcache__s2_req_addr  [1] ?   dcache__io_cpu_resp_bits_data_zeroed  [31:16]:  dcache__io_cpu_resp_bits_data_zeroed  [15:0]; 
   wire[7:0]  dcache__io_cpu_resp_bits_data_zeroed_2  =  dcache__s2_sc   ? 8'h0:  dcache__s2_req_addr  [0] ?   dcache__io_cpu_resp_bits_data_zeroed_1  [15:8]:  dcache__io_cpu_resp_bits_data_zeroed_1  [7:0]; 
   wire[31:0]  dcache__io_cpu_resp_bits_data_word_bypass_zeroed  =  dcache__s2_req_addr  [2] ?   dcache__s2_data  [63:32]:  dcache__s2_data  [31:0]; 
   reg  dcache__REG  ; 
   wire[26:0]  dcache___io_cpu_perf_release_beats1_decode_T_1  =27'hFFF<<  dcache___GEN_23  ; 
   wire[8:0]  dcache__io_cpu_perf_release_beats1  =  dcache__nodeOut_c_bits_opcode  [0] ? ~(  dcache___io_cpu_perf_release_beats1_decode_T_1  [11:3]):9'h0; 
   reg[8:0]  dcache__io_cpu_perf_release_counter  ; 
   wire[3:0]  dcache___release_state_T_14  =  dcache__s2_victim_dirty  &~(  dcache__s2_valid_flush_line  &  dcache__s2_req_size  [1]) ? 4'h1:4'h6; 
   wire[3:0]  dcache___release_state_T_15  ={1'h0,  dcache__releaseDone  ,2'h3}; 
   wire[3:0]  dcache___GEN_29  =  dcache__s2_prb_ack_data   ? 4'h2:(|  dcache__s2_probe_state_state  ) ? 4'h3:4'h5; 
   wire[3:0]  dcache___GEN_30  =  dcache__s2_want_victimize   ?   dcache___release_state_T_14  :  dcache__release_state  ; 
   wire[3:0]  dcache___GEN_31  =  dcache__s2_probe   ?   dcache___GEN_29  :  dcache___GEN_30  ; 
   wire  dcache___GEN_32  =  dcache___io_errors_bus_valid_T  &  dcache__grantIsCached  &  dcache__d_last  ; 
   wire  dcache___GEN_33  =  dcache___GEN_24  &~  dcache__metaArb__grant_T_3  ; 
   wire[6:0]  dcache__flushCounterNext  ={1'h0,  dcache__flushCounter  }+7'h1; 
   wire  dcache___GEN_34  =  dcache___GEN_25  &  dcache__releaseDone  |  dcache___GEN_33  ; 
   wire[33:0]  dcache__s0_req_addr  ={  dcache__resetting   ? {  dcache__io_cpu_req_bits_addr  [33:12],  dcache__flushCounter  }:  dcache___GEN   ? {  dcache__io_cpu_req_bits_addr  [33:12],  dcache__s2_req_addr  [11:6]}:  dcache__metaArb_io_in_valid_4   ? {  dcache__io_cpu_req_bits_addr  [33:12],  dcache__probe_bits_address  [11:6]}:  dcache__metaArb_io_in_valid_6   ? {  dcache__io_cpu_req_bits_addr  [33:32],  dcache___GEN_24   ?   dcache__probe_bits_address  [31:6]:  dcache__auto_out_b_bits_address  [31:6]}:  dcache__io_cpu_req_bits_addr  [33:6],  dcache__io_cpu_req_bits_addr  [5:0]}; 
   wire[9:0]  dcache___GEN_35  =  dcache__s1_tlb_req_vaddr  [25:16]^10'h200; 
   wire[3:0]  dcache___GEN_36  =  dcache__s1_tlb_req_vaddr  [31:28]^4'h8; 
   wire  dcache__tlb_legal_address  ={  dcache__s1_tlb_req_vaddr  [33:14],~(  dcache__s1_tlb_req_vaddr  [13:12])}==22'h0|{  dcache__s1_tlb_req_vaddr  [33:28],~(  dcache__s1_tlb_req_vaddr  [27:26])}==8'h0|{  dcache__s1_tlb_req_vaddr  [33:26],  dcache___GEN_35  }==18'h0|~(|(  dcache__s1_tlb_req_vaddr  [33:12]))|{  dcache__s1_tlb_req_vaddr  [33:17],~(  dcache__s1_tlb_req_vaddr  [16])}==18'h0|{  dcache__s1_tlb_req_vaddr  [33:32],  dcache___GEN_36  }==6'h0|{  dcache__s1_tlb_req_vaddr  [33:31],~(  dcache__s1_tlb_req_vaddr  [30:29])}==5'h0; 
   wire  dcache__tlb_cacheable  =  dcache__tlb_legal_address  &~(  dcache___GEN_36  [3]); 
   wire  dcache__tlb_deny_access_to_debug  =~  dcache__io_ptw_status_debug  &~(|(  dcache__s1_tlb_req_vaddr  [33:12])); 
   wire[3:0]  dcache___GEN_37  ={  dcache__s1_tlb_req_vaddr  [31:30],  dcache__s1_tlb_req_vaddr  [27],  dcache__s1_tlb_req_vaddr  [16]}; 
   wire[2:0]  dcache___GEN_38  ={  dcache__s1_tlb_req_vaddr  [31:30],~(  dcache__s1_tlb_req_vaddr  [27])}; 
   wire[1:0]  dcache___GEN_39  ={  dcache__s1_tlb_req_vaddr  [31],~(  dcache__s1_tlb_req_vaddr  [30])}; 
   wire[3:0]  dcache___GEN_40  =  dcache__s1_tlb_req_vaddr  [3:0]&(4'h1<<  dcache__s1_tlb_req_size  )-4'h1; 
   wire  dcache__tlb__cmd_lrsc_T  =  dcache__s1_tlb_req_cmd  ==5'h6; 
   wire  dcache__tlb__cmd_lrsc_T_1  =  dcache__s1_tlb_req_cmd  ==5'h7; 
   wire  dcache__tlb__cmd_read_T_7  =  dcache__s1_tlb_req_cmd  ==5'h4; 
   wire  dcache__tlb__cmd_read_T_8  =  dcache__s1_tlb_req_cmd  ==5'h9; 
   wire  dcache__tlb__cmd_read_T_9  =  dcache__s1_tlb_req_cmd  ==5'hA; 
   wire  dcache__tlb__cmd_read_T_10  =  dcache__s1_tlb_req_cmd  ==5'hB; 
   wire  dcache__tlb__cmd_read_T_14  =  dcache__s1_tlb_req_cmd  ==5'h8; 
   wire  dcache__tlb__cmd_read_T_15  =  dcache__s1_tlb_req_cmd  ==5'hC; 
   wire  dcache__tlb__cmd_read_T_16  =  dcache__s1_tlb_req_cmd  ==5'hD; 
   wire  dcache__tlb__cmd_read_T_17  =  dcache__s1_tlb_req_cmd  ==5'hE; 
   wire  dcache__tlb__cmd_read_T_18  =  dcache__s1_tlb_req_cmd  ==5'hF; 
   wire  dcache__tlb_cmd_put_partial  =  dcache__s1_tlb_req_cmd  ==5'h11; 
   wire  dcache__tlb_cmd_read  =  dcache__s1_tlb_req_cmd  ==5'h0|  dcache__s1_tlb_req_cmd  ==5'h10|  dcache__tlb__cmd_lrsc_T  |  dcache__tlb__cmd_lrsc_T_1  |  dcache__tlb__cmd_read_T_7  |  dcache__tlb__cmd_read_T_8  |  dcache__tlb__cmd_read_T_9  |  dcache__tlb__cmd_read_T_10  |  dcache__tlb__cmd_read_T_14  |  dcache__tlb__cmd_read_T_15  |  dcache__tlb__cmd_read_T_16  |  dcache__tlb__cmd_read_T_17  |  dcache__tlb__cmd_read_T_18  ; 
   wire  dcache__tlb_cmd_write  =  dcache__s1_tlb_req_cmd  ==5'h1|  dcache__tlb_cmd_put_partial  |  dcache__tlb__cmd_lrsc_T_1  |  dcache__tlb__cmd_read_T_7  |  dcache__tlb__cmd_read_T_8  |  dcache__tlb__cmd_read_T_9  |  dcache__tlb__cmd_read_T_10  |  dcache__tlb__cmd_read_T_14  |  dcache__tlb__cmd_read_T_15  |  dcache__tlb__cmd_read_T_16  |  dcache__tlb__cmd_read_T_17  |  dcache__tlb__cmd_read_T_18  ; 
   wire  dcache__tlb_ae_array  =(|  dcache___GEN_40  )&  dcache__tlb_legal_address  &({  dcache__s1_tlb_req_vaddr  [31:30],  dcache__s1_tlb_req_vaddr  [27],  dcache__s1_tlb_req_vaddr  [25],  dcache__s1_tlb_req_vaddr  [16],  dcache__s1_tlb_req_vaddr  [13]}==6'h0|{  dcache__s1_tlb_req_vaddr  [31:30],  dcache__s1_tlb_req_vaddr  [27],  dcache___GEN_35  [9],  dcache__s1_tlb_req_vaddr  [16]}==5'h0|~(|  dcache___GEN_38  )|~(|  dcache___GEN_39  ))|(  dcache__tlb__cmd_lrsc_T  |  dcache__tlb__cmd_lrsc_T_1  )&~  dcache__tlb_cacheable  ; 
   wire[1:0]  dcache___s2_data_T_1  =  dcache__io_cpu_replay_next_0  |  dcache__inWriteback  |  dcache__s1_did_read   ? (  dcache___GEN_19   ? 2'h1:2'h2):2'h0; 
   wire  dcache___probe_bits_T  =  dcache__nodeOut_b_ready  &  dcache__auto_out_b_valid  ; 
   wire  dcache__s1_valid_not_nacked  =  dcache__s1_valid  &~  dcache__s1_nack  ; 
   wire  dcache___s1_meta_hit_state_T_2  =  dcache___tag_array_0_ext_RW0_rdata  [19:0]==  dcache__s1_tlb_req_vaddr  [31:12]&~  dcache__s1_flush_valid  ; 
   wire  dcache___s2_victim_way_T  =  dcache__s1_valid_not_nacked  |  dcache__s1_flush_valid  ; 
   wire  dcache___GEN_41  =  dcache__s2_valid_hit_pre_data_ecc_and_waw  &  dcache__s2_lr  &~  dcache__cached_grant_wait  |  dcache__s2_valid_cached_miss  ; 
   wire  dcache__advance_pstore1  =  dcache__pstore1_valid  &  dcache__pstore2_valid  ==  dcache__pstore_drain  ; 
   wire  dcache___io_cpu_perf_acquire_T  =  dcache__auto_out_a_ready  &  dcache__tl_out_a_valid  ; 
   wire  dcache___GEN_42  =  dcache___io_cpu_perf_acquire_T  &~  dcache__s2_pma_cacheable  ; 
   wire  dcache___GEN_43  =  dcache___GEN_27  &  dcache___io_cpu_perf_release_T  &  dcache__c_first  ; 
  always @( posedge   dcache__clock  )
       begin 
         if (  dcache__reset  )
            begin  
               dcache__s1_valid   <=1'h0; 
               dcache__s1_probe   <=1'h0; 
               dcache__cached_grant_wait   <=1'h0; 
               dcache__resetting   <=1'h0; 
               dcache__flushCounter   <=6'h0; 
               dcache__release_ack_wait   <=1'h0; 
               dcache__release_state   <=4'h0; 
               dcache__uncachedInFlight_0   <=1'h0; 
               dcache__s2_valid   <=1'h0; 
               dcache__s2_probe   <=1'h0; 
               dcache__lrscCount   <=7'h0; 
               dcache__pstore2_valid   <=1'h0; 
               dcache__pstore1_held   <=1'h0; 
               dcache__counter   <=9'h0; 
               dcache__grantInProgress   <=1'h0; 
               dcache__blockProbeAfterGrantCount   <=3'h0; 
               dcache__counter_1   <=9'h0; 
               dcache__io_cpu_perf_release_counter   <=9'h0;
            end 
          else 
            begin  
               dcache__s1_valid   <=  dcache__io_cpu_req_ready_0  &  dcache__io_cpu_req_valid  ; 
               dcache__s1_probe   <=  dcache___GEN_33  |  dcache___probe_bits_T  ; 
               dcache__cached_grant_wait   <=~  dcache___GEN_32  &(  dcache___io_cpu_perf_acquire_T  &  dcache__s2_pma_cacheable  |  dcache__cached_grant_wait  ); 
               dcache__resetting   <=~(  dcache__resetting  &  dcache__flushCounterNext  [6])&(  dcache__REG  |  dcache__resetting  );
              if (  dcache__resetting  ) 
                  dcache__flushCounter   <=  dcache__flushCounterNext  [5:0]; 
               dcache__release_ack_wait   <=  dcache___GEN_43  |(~  dcache___io_errors_bus_valid_T  |  dcache__grantIsCached  |  dcache__grantIsUncached  |~  dcache__grantIsVoluntary  )&  dcache__release_ack_wait  ;
              if (~  dcache__metaArb__grant_T_2  &  dcache__metaArb_io_in_valid_4  ) 
                  dcache__release_state   <=4'h0;
               else 
                 if (  dcache___GEN_27  )
                    begin 
                      if (  dcache__releaseDone  ) 
                          dcache__release_state   <=4'h6;
                       else 
                         if (  dcache___GEN_26  ) 
                             dcache__release_state   <=  dcache___inWriteback_T_1   ? (  dcache___GEN_34   ? 4'h0:  dcache___GEN_31  ):  dcache___GEN_25   ? (  dcache__releaseDone  |  dcache___GEN_33   ? 4'h0:  dcache___GEN_31  ):  dcache___GEN_33   ? 4'h0:  dcache__s2_probe   ? (  dcache__s2_prb_ack_data   ? 4'h2:(|  dcache__s2_probe_state_state  ) ? 4'h3:  dcache__releaseDone   ? 4'h0:4'h5):  dcache___GEN_30  ;
                          else 
                            if (  dcache___GEN_34  ) 
                                dcache__release_state   <=4'h0;
                             else 
                               if (  dcache__s2_probe  )
                                  begin 
                                    if (  dcache__s2_prb_ack_data  ) 
                                        dcache__release_state   <=4'h2;
                                     else 
                                       if (|  dcache__s2_probe_state_state  ) 
                                           dcache__release_state   <=  dcache___release_state_T_15  ;
                                        else 
                                          if (  dcache__releaseDone  ) 
                                              dcache__release_state   <=4'h0;
                                           else  
                                              dcache__release_state   <=4'h5;
                                  end 
                                else 
                                  if (  dcache__s2_want_victimize  ) 
                                      dcache__release_state   <=  dcache___release_state_T_14  ;
                    end 
                  else 
                    if (  dcache___inWriteback_T_1  )
                       begin 
                         if (  dcache__releaseDone  ) 
                             dcache__release_state   <=4'h7;
                          else 
                            if (  dcache___GEN_34  ) 
                                dcache__release_state   <=4'h0;
                             else 
                               if (  dcache__s2_probe  ) 
                                   dcache__release_state   <=  dcache___GEN_29  ;
                                else 
                                  if (  dcache__s2_want_victimize  ) 
                                      dcache__release_state   <=  dcache___release_state_T_14  ;
                       end 
                     else 
                       if (  dcache___GEN_26  )
                          begin 
                            if (  dcache__releaseDone  ) 
                                dcache__release_state   <=4'h7;
                             else 
                               if (  dcache___GEN_34  ) 
                                   dcache__release_state   <=4'h0;
                                else 
                                  if (  dcache__s2_probe  ) 
                                      dcache__release_state   <=  dcache___GEN_29  ;
                                   else 
                                     if (  dcache__s2_want_victimize  ) 
                                         dcache__release_state   <=  dcache___release_state_T_14  ;
                          end 
                        else 
                          if (  dcache___GEN_34  ) 
                              dcache__release_state   <=4'h0;
                           else 
                             if (  dcache__s2_probe  )
                                begin 
                                  if (  dcache__s2_prb_ack_data  ) 
                                      dcache__release_state   <=4'h2;
                                   else 
                                     if (|  dcache__s2_probe_state_state  ) 
                                         dcache__release_state   <=  dcache___release_state_T_15  ;
                                      else 
                                        if (  dcache__releaseDone  ) 
                                            dcache__release_state   <=4'h0;
                                         else  
                                            dcache__release_state   <=4'h5;
                                end 
                              else 
                                if (  dcache__s2_want_victimize  ) 
                                    dcache__release_state   <=  dcache___release_state_T_14  ; 
               dcache__uncachedInFlight_0   <=(~  dcache___io_errors_bus_valid_T  |  dcache__grantIsCached  |~(  dcache__grantIsUncached  &  dcache___GEN_18  ))&(  dcache___GEN_42  |  dcache__uncachedInFlight_0  ); 
               dcache__s2_valid   <=  dcache__s1_valid_masked  &~(  dcache__s1_req_cmd  ==5'h14|  dcache__s1_req_cmd  ==5'h15|  dcache__s1_req_cmd  ==5'h16); 
               dcache__s2_probe   <=  dcache__s1_probe  ;
              if (  dcache__s1_probe  ) 
                  dcache__lrscCount   <=7'h0;
               else 
                 if (  dcache__s2_valid_masked  &(|(  dcache__lrscCount  [6:2]))) 
                     dcache__lrscCount   <=7'h3;
                  else 
                    if (|  dcache__lrscCount  ) 
                        dcache__lrscCount   <=  dcache__lrscCount  -7'h1;
                     else 
                       if (  dcache___GEN_41  ) 
                           dcache__lrscCount   <=  dcache__s2_hit   ? 7'h4F:7'h0; 
               dcache__pstore2_valid   <=  dcache__pstore2_valid  &~  dcache__pstore_drain  |  dcache__advance_pstore1  ; 
               dcache__pstore1_held   <=(  dcache___pstore1_held_T  &~  dcache__s2_sc_fail  |  dcache__pstore1_held  )&  dcache__pstore2_valid  &~  dcache__pstore_drain  ;
              if (  dcache___io_errors_bus_valid_T  )
                 begin 
                   if (|  dcache__counter  ) 
                       dcache__counter   <=  dcache___counter1_T  ;
                    else  
                       dcache__counter   <=  dcache__beats1  ;
                 end 
              if (  dcache___GEN_17  ) 
                  dcache__grantInProgress   <=~  dcache__d_last  ;
              if (  dcache___GEN_32  ) 
                  dcache__blockProbeAfterGrantCount   <=3'h7;
               else 
                 if (|  dcache__blockProbeAfterGrantCount  ) 
                     dcache__blockProbeAfterGrantCount   <=  dcache__blockProbeAfterGrantCount  -3'h1;
              if (  dcache___io_cpu_perf_release_T  )
                 begin 
                   if (  dcache__c_first  ) 
                       dcache__counter_1   <=  dcache__beats1_1  ;
                    else  
                       dcache__counter_1   <=  dcache___counter1_T_1  ;
                   if (  dcache__io_cpu_perf_release_counter  ==9'h0) 
                       dcache__io_cpu_perf_release_counter   <=  dcache__io_cpu_perf_release_beats1  ;
                    else  
                       dcache__io_cpu_perf_release_counter   <=  dcache__io_cpu_perf_release_counter  -9'h1;
                 end 
            end 
         if (  dcache__s2_want_victimize  )
            begin  
               dcache__probe_bits_param   <=2'h0; 
               dcache__probe_bits_size   <=4'h0; 
               dcache__probe_bits_address   <={  dcache__s2_valid_flush_line   ?   dcache__s2_req_addr  [31:12]:  dcache__s2_meta_corrected_r  [19:0],  dcache__s2_req_addr  [11:6],6'h0};
            end 
          else 
            if (  dcache___probe_bits_T  )
               begin  
                  dcache__probe_bits_param   <=  dcache__auto_out_b_bits_param  ; 
                  dcache__probe_bits_size   <=  dcache__auto_out_b_bits_size  ; 
                  dcache__probe_bits_address   <=  dcache__auto_out_b_bits_address  ;
               end  
          dcache__probe_bits_source   <=~  dcache__s2_want_victimize  &(  dcache___probe_bits_T   ?   dcache__auto_out_b_bits_source  :  dcache__probe_bits_source  );
         if (  dcache__metaArb_io_out_valid  &~  dcache__metaArb_io_out_bits_write  )
            begin  
               dcache__s1_vaddr   <=  dcache__s0_req_addr  ; 
               dcache__s1_req_tag   <=  dcache__io_cpu_req_bits_tag  ; 
               dcache__s1_req_cmd   <=  dcache__io_cpu_req_bits_cmd  ; 
               dcache__s1_req_size   <=  dcache__io_cpu_req_bits_size  ; 
               dcache__s1_req_signed   <=  dcache__io_cpu_req_bits_signed  ; 
               dcache__s1_req_dprv   <=2'h3; 
               dcache__s1_req_dv   <=  dcache__io_cpu_req_bits_dv  ; 
               dcache__s1_tlb_req_vaddr   <=  dcache__s0_req_addr  ; 
               dcache__s1_tlb_req_size   <=  dcache__io_cpu_req_bits_size  ; 
               dcache__s1_tlb_req_cmd   <=  dcache__io_cpu_req_bits_cmd  ; 
               dcache__s1_tlb_req_prv   <=2'h3; 
               dcache__s1_did_read   <=~  dcache__dataArb__grant_T_1  &  dcache__io_cpu_req_valid  &(  dcache___pstore_drain_opportunistic_T  |  dcache___pstore_drain_opportunistic_T_1  |  dcache___pstore_drain_opportunistic_T_2  |  dcache___pstore_drain_opportunistic_T_28  |  dcache___pstore_drain_opportunistic_T_30  |  dcache___pstore_drain_opportunistic_T_31  |  dcache___pstore_drain_opportunistic_T_32  |  dcache___pstore_drain_opportunistic_T_33  |  dcache___pstore_drain_opportunistic_T_37  |  dcache___pstore_drain_opportunistic_T_38  |  dcache___pstore_drain_opportunistic_T_39  |  dcache___pstore_drain_opportunistic_T_40  |  dcache___pstore_drain_opportunistic_T_41  |(  dcache___pstore_drain_opportunistic_T_25  |  dcache___pstore_drain_opportunistic_T_50  |  dcache___pstore_drain_opportunistic_T_28  |  dcache___pstore_drain_opportunistic_T_30  |  dcache___pstore_drain_opportunistic_T_31  |  dcache___pstore_drain_opportunistic_T_32  |  dcache___pstore_drain_opportunistic_T_33  |  dcache___pstore_drain_opportunistic_T_37  |  dcache___pstore_drain_opportunistic_T_38  |  dcache___pstore_drain_opportunistic_T_39  |  dcache___pstore_drain_opportunistic_T_40  |  dcache___pstore_drain_opportunistic_T_41  )&  dcache___pstore_drain_opportunistic_T_50  );
            end  
          dcache__s1_flush_valid   <=1'h0;
         if (  dcache___GEN_43  ) 
             dcache__release_ack_addr   <=  dcache__probe_bits_address  ;
         if (  dcache___GEN_42  )
            begin  
               dcache__uncachedReqs_addr_0   <=  dcache__s2_req_addr  ; 
               dcache__uncachedReqs_tag_0   <=  dcache__s2_req_tag  ; 
               dcache__uncachedReqs_size_0   <=  dcache__s2_req_size  ; 
               dcache__uncachedReqs_signed_0   <=  dcache__s2_req_signed  ;
            end  
          dcache__s2_not_nacked_in_s1   <=~  dcache__s1_nack  ;
         if (  dcache___GEN_19  )
            begin 
              if (  dcache___s2_victim_way_T  )
                 begin  
                    dcache__s2_req_addr   <={2'h0,  dcache__s1_tlb_req_vaddr  [31:12],  dcache__s1_vaddr  [11:0]}; 
                    dcache__s2_req_tag   <=  dcache__s1_req_tag  ; 
                    dcache__s2_req_cmd   <=  dcache__s1_req_cmd  ; 
                    dcache__s2_req_size   <=  dcache__s1_req_size  ; 
                    dcache__s2_req_signed   <=  dcache__s1_req_signed  ;
                 end 
            end 
          else 
            begin  
               dcache__s2_req_addr   <={2'h0,  dcache__s1_tlb_req_vaddr  [31:12],  dcache__s1_vaddr  [11:3],  dcache__uncachedReqs_addr_0  [2:0]}; 
               dcache__s2_req_tag   <=  dcache__uncachedReqs_tag_0  ; 
               dcache__s2_req_cmd   <=5'h0; 
               dcache__s2_req_size   <=  dcache__uncachedReqs_size_0  ; 
               dcache__s2_req_signed   <=  dcache__uncachedReqs_signed_0  ;
            end 
         if (  dcache___s2_victim_way_T  )
            begin  
               dcache__s2_req_dprv   <=  dcache__s1_req_dprv  ; 
               dcache__s2_req_dv   <=  dcache__s1_req_dv  ; 
               dcache__s2_tlb_xcpt_ae_ld   <=  dcache__tlb_cmd_read  &(  dcache__tlb_ae_array  |~(  dcache__tlb_legal_address  &~  dcache__tlb_deny_access_to_debug  &  dcache___tlb_pmp_io_r  )); 
               dcache__s2_tlb_xcpt_ae_st   <=(  dcache__tlb_cmd_write  |  dcache__s1_tlb_req_cmd  ==5'h5|  dcache__s1_tlb_req_cmd  ==5'h17)&(  dcache__tlb_ae_array  |~(  dcache__tlb_legal_address  &(~(|  dcache___GEN_37  )|~(|  dcache___GEN_38  )|~(|  dcache___GEN_39  )|~(|(  dcache___GEN_36  [3:2])))&~  dcache__tlb_deny_access_to_debug  &  dcache___tlb_pmp_io_w  ))|  dcache__tlb_cmd_put_partial  &~(  dcache__tlb_legal_address  &(~(|  dcache___GEN_37  )|~(|  dcache___GEN_38  )|~(|  dcache___GEN_39  )|~(|(  dcache___GEN_36  [3:2])))|  dcache__tlb_cacheable  )|(  dcache__tlb__cmd_read_T_7  |  dcache__tlb__cmd_read_T_8  |  dcache__tlb__cmd_read_T_9  |  dcache__tlb__cmd_read_T_10  )&~(  dcache__tlb_legal_address  &(~(|  dcache___GEN_37  )|~(|  dcache___GEN_38  ))|  dcache__tlb_cacheable  )|(  dcache__tlb__cmd_read_T_14  |  dcache__tlb__cmd_read_T_15  |  dcache__tlb__cmd_read_T_16  |  dcache__tlb__cmd_read_T_17  |  dcache__tlb__cmd_read_T_18  )&~(  dcache__tlb_legal_address  &(~(|  dcache___GEN_37  )|~(|  dcache___GEN_38  ))|  dcache__tlb_cacheable  ); 
               dcache__s2_tlb_xcpt_ma_ld   <=(|  dcache___GEN_40  )&  dcache__tlb_cmd_read  ; 
               dcache__s2_tlb_xcpt_ma_st   <=(|  dcache___GEN_40  )&  dcache__tlb_cmd_write  ; 
               dcache__s2_pma_cacheable   <=  dcache__tlb_cacheable  ; 
               dcache__s2_vaddr_r   <=  dcache__s1_vaddr  ;
              if (  dcache___s1_meta_hit_state_T_2  ) 
                  dcache__s2_hit_state_state   <=  dcache___tag_array_0_ext_RW0_rdata  [21:20];
               else  
                  dcache__s2_hit_state_state   <=2'h0;
            end  
          dcache__s2_tlb_xcpt_pf_ld   <=~  dcache___s2_victim_way_T  &  dcache__s2_tlb_xcpt_pf_ld  ; 
          dcache__s2_tlb_xcpt_pf_st   <=~  dcache___s2_victim_way_T  &  dcache__s2_tlb_xcpt_pf_st  ;
         if (  dcache___GEN_19  )
            begin 
            end 
          else  
             dcache__s2_uncached_resp_addr   <=  dcache__uncachedReqs_addr_0  ; 
          dcache__s2_flush_valid   <=  dcache__s1_flush_valid  ;
         if (  dcache___s2_victim_way_T  |  dcache__s1_probe  ) 
             dcache__s2_meta_corrected_r   <=  dcache___tag_array_0_ext_RW0_rdata  ;
         if (  dcache__s1_valid  |  dcache__inWriteback  |  dcache__io_cpu_replay_next_0  ) 
             dcache__s2_data   <=(  dcache___s2_data_T_1  [0] ?   dcache___data_io_resp_0  :64'h0)|(  dcache___s2_data_T_1  [1] ?   dcache__auto_out_d_bits_data  :64'h0);
         if (  dcache__s1_probe  )
            begin 
              if (  dcache___s1_meta_hit_state_T_2  ) 
                  dcache__s2_probe_state_state   <=  dcache___tag_array_0_ext_RW0_rdata  [21:20];
               else  
                  dcache__s2_probe_state_state   <=2'h0;
            end 
         if (  dcache___GEN_41  ) 
             dcache__lrscAddr   <=  dcache__s2_req_addr  [33:6];
         if (  dcache__s1_valid_not_nacked  &  dcache__s1_write  )
            begin  
               dcache__pstore1_cmd   <=  dcache__s1_req_cmd  ; 
               dcache__pstore1_addr   <=  dcache__s1_vaddr  ; 
               dcache__pstore1_data   <=  dcache__io_cpu_s1_data_data  ; 
               dcache__pstore1_mask   <=  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_51   ?   dcache__io_cpu_s1_data_mask  :  dcache__s1_mask_xwr  ; 
               dcache__pstore1_rmw   <=  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_1  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_2  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_3  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_29  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_31  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_32  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_33  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_34  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_38  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_39  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_40  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_41  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_42  |(  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_26  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_51  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_29  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_31  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_32  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_33  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_34  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_38  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_39  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_40  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_41  |  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_42  )&  dcache___io_cpu_perf_canAcceptLoadThenLoad_T_51  ;
            end  
          dcache__pstore_drain_on_miss_REG   <=  dcache__io_cpu_s2_nack_0  ;
         if (  dcache__advance_pstore1  )
            begin  
               dcache__pstore2_addr   <=  dcache__pstore1_addr  ; 
               dcache__pstore2_storegen_data_r   <=  dcache___amoalus_0_io_out  [7:0]; 
               dcache__pstore2_storegen_data_r_1   <=  dcache___amoalus_0_io_out  [15:8]; 
               dcache__pstore2_storegen_data_r_2   <=  dcache___amoalus_0_io_out  [23:16]; 
               dcache__pstore2_storegen_data_r_3   <=  dcache___amoalus_0_io_out  [31:24]; 
               dcache__pstore2_storegen_data_r_4   <=  dcache___amoalus_0_io_out  [39:32]; 
               dcache__pstore2_storegen_data_r_5   <=  dcache___amoalus_0_io_out  [47:40]; 
               dcache__pstore2_storegen_data_r_6   <=  dcache___amoalus_0_io_out  [55:48]; 
               dcache__pstore2_storegen_data_r_7   <=  dcache___amoalus_0_io_out  [63:56]; 
               dcache__pstore2_storegen_mask   <=  dcache__pstore1_mask  ;
            end 
         if (  dcache___GEN_22  ) 
             dcache__blockUncachedGrant   <=  dcache__dataArb_io_in_valid_0  ;
          else  
             dcache__blockUncachedGrant   <=  dcache__dataArb_io_out_valid  ; 
          dcache__s1_release_data_valid   <=~  dcache__dataArb__grant_T  &  dcache__dataArb_io_in_valid_2  ; 
          dcache__s2_release_data_valid   <=  dcache__s1_release_data_valid  &~  dcache__releaseRejected  ; 
          dcache__io_cpu_s2_xcpt_REG   <=  dcache__s1_valid  &~  dcache__io_cpu_s1_kill  &(  dcache__s1_read  |  dcache__s1_write  |  dcache__s1_req_cmd  ==5'h5&  dcache__s1_req_size  [0]|  dcache__s1_req_cmd  ==5'h17)&~  dcache__s1_nack  ; 
          dcache__doUncachedResp   <=  dcache__io_cpu_replay_next_0  ; 
          dcache__REG   <=  dcache__reset  ;
       end
   
  
wire [1:0] dcache__tlb_pmp__io_prv;
wire  dcache__tlb_pmp__io_pmp_cfg_l_0;
wire  dcache__tlb_pmp__io_pmp_cfg_l_1;
wire  dcache__tlb_pmp__io_pmp_cfg_l_2;
wire  dcache__tlb_pmp__io_pmp_cfg_l_3;
wire  dcache__tlb_pmp__io_pmp_cfg_l_4;
wire  dcache__tlb_pmp__io_pmp_cfg_l_5;
wire  dcache__tlb_pmp__io_pmp_cfg_l_6;
wire  dcache__tlb_pmp__io_pmp_cfg_l_7;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_0;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_1;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_2;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_3;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_4;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_5;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_6;
wire [1:0] dcache__tlb_pmp__io_pmp_cfg_a_7;
wire  dcache__tlb_pmp__io_pmp_cfg_w_0;
wire  dcache__tlb_pmp__io_pmp_cfg_w_1;
wire  dcache__tlb_pmp__io_pmp_cfg_w_2;
wire  dcache__tlb_pmp__io_pmp_cfg_w_3;
wire  dcache__tlb_pmp__io_pmp_cfg_w_4;
wire  dcache__tlb_pmp__io_pmp_cfg_w_5;
wire  dcache__tlb_pmp__io_pmp_cfg_w_6;
wire  dcache__tlb_pmp__io_pmp_cfg_w_7;
wire  dcache__tlb_pmp__io_pmp_cfg_r_0;
wire  dcache__tlb_pmp__io_pmp_cfg_r_1;
wire  dcache__tlb_pmp__io_pmp_cfg_r_2;
wire  dcache__tlb_pmp__io_pmp_cfg_r_3;
wire  dcache__tlb_pmp__io_pmp_cfg_r_4;
wire  dcache__tlb_pmp__io_pmp_cfg_r_5;
wire  dcache__tlb_pmp__io_pmp_cfg_r_6;
wire  dcache__tlb_pmp__io_pmp_cfg_r_7;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_0;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_1;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_2;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_3;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_4;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_5;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_6;
wire [29:0] dcache__tlb_pmp__io_pmp_addr_7;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_0;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_1;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_2;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_3;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_4;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_5;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_6;
wire [31:0] dcache__tlb_pmp__io_pmp_mask_7;
wire [31:0] dcache__tlb_pmp__io_addr;
wire [1:0] dcache__tlb_pmp__io_size;
wire  dcache__tlb_pmp__io_r;
wire  dcache__tlb_pmp__io_w;
 
   wire[5:0]  dcache__tlb_pmp___GEN  ={4'h0,  dcache__tlb_pmp__io_size  }; 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_1  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[5:0]  dcache__tlb_pmp___res_hit_T_4  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit  =  dcache__tlb_pmp__io_pmp_cfg_a_7  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_7  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_7  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_7  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_7  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_1  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_7  [0]&~(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_6  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_6  [29:1])==29'h0&(  dcache__tlb_pmp__io_addr  [2:0]|~(  dcache__tlb_pmp___res_hit_T_4  [2:0]))<{  dcache__tlb_pmp__io_pmp_addr_6  [0],2'h0})&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_7  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_7  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_7  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_7  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_1  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_1  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned  =  dcache__tlb_pmp__io_pmp_cfg_a_7  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask  &~(  dcache__tlb_pmp__io_pmp_mask_7  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_6  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_6  [0]&~(  dcache__tlb_pmp__io_addr  [2])|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_7  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_7  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask  [2])); 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_5  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[5:0]  dcache__tlb_pmp___res_hit_T_18  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit_1  =  dcache__tlb_pmp__io_pmp_cfg_a_6  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_6  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_6  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_6  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_6  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_5  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_6  [0]&~(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_5  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_5  [29:1])==29'h0&(  dcache__tlb_pmp__io_addr  [2:0]|~(  dcache__tlb_pmp___res_hit_T_18  [2:0]))<{  dcache__tlb_pmp__io_pmp_addr_5  [0],2'h0})&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_6  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_6  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_6  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore_1  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_6  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_4  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask_1  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_4  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned_1  =  dcache__tlb_pmp__io_pmp_cfg_a_6  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask_1  &~(  dcache__tlb_pmp__io_pmp_mask_6  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_5  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_5  [0]&~(  dcache__tlb_pmp__io_addr  [2])|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_6  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_6  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask_1  [2])); 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_9  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[5:0]  dcache__tlb_pmp___res_hit_T_32  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit_2  =  dcache__tlb_pmp__io_pmp_cfg_a_5  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_5  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_5  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_5  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_5  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_9  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_5  [0]&~(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_4  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_4  [29:1])==29'h0&(  dcache__tlb_pmp__io_addr  [2:0]|~(  dcache__tlb_pmp___res_hit_T_32  [2:0]))<{  dcache__tlb_pmp__io_pmp_addr_4  [0],2'h0})&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_5  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_5  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_5  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore_2  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_5  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_7  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask_2  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_7  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned_2  =  dcache__tlb_pmp__io_pmp_cfg_a_5  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask_2  &~(  dcache__tlb_pmp__io_pmp_mask_5  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_4  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_4  [0]&~(  dcache__tlb_pmp__io_addr  [2])|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_5  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_5  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask_2  [2])); 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_13  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[5:0]  dcache__tlb_pmp___res_hit_T_46  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit_3  =  dcache__tlb_pmp__io_pmp_cfg_a_4  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_4  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_4  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_4  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_4  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_13  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_4  [0]&~(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_3  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_3  [29:1])==29'h0&(  dcache__tlb_pmp__io_addr  [2:0]|~(  dcache__tlb_pmp___res_hit_T_46  [2:0]))<{  dcache__tlb_pmp__io_pmp_addr_3  [0],2'h0})&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_4  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_4  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_4  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore_3  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_4  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_10  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask_3  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_10  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned_3  =  dcache__tlb_pmp__io_pmp_cfg_a_4  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask_3  &~(  dcache__tlb_pmp__io_pmp_mask_4  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_3  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_3  [0]&~(  dcache__tlb_pmp__io_addr  [2])|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_4  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_4  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask_3  [2])); 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_17  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[5:0]  dcache__tlb_pmp___res_hit_T_60  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit_4  =  dcache__tlb_pmp__io_pmp_cfg_a_3  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_3  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_3  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_3  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_3  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_17  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_3  [0]&~(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_2  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_2  [29:1])==29'h0&(  dcache__tlb_pmp__io_addr  [2:0]|~(  dcache__tlb_pmp___res_hit_T_60  [2:0]))<{  dcache__tlb_pmp__io_pmp_addr_2  [0],2'h0})&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_3  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_3  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_3  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore_4  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_3  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_13  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask_4  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_13  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned_4  =  dcache__tlb_pmp__io_pmp_cfg_a_3  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask_4  &~(  dcache__tlb_pmp__io_pmp_mask_3  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_2  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_2  [0]&~(  dcache__tlb_pmp__io_addr  [2])|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_3  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_3  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask_4  [2])); 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_21  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[5:0]  dcache__tlb_pmp___res_hit_T_74  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit_5  =  dcache__tlb_pmp__io_pmp_cfg_a_2  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_2  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_2  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_2  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_2  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_21  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_2  [0]&~(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_1  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_1  [29:1])==29'h0&(  dcache__tlb_pmp__io_addr  [2:0]|~(  dcache__tlb_pmp___res_hit_T_74  [2:0]))<{  dcache__tlb_pmp__io_pmp_addr_1  [0],2'h0})&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_2  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_2  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_2  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore_5  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_2  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_16  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask_5  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_16  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned_5  =  dcache__tlb_pmp__io_pmp_cfg_a_2  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask_5  &~(  dcache__tlb_pmp__io_pmp_mask_2  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_1  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_1  [0]&~(  dcache__tlb_pmp__io_addr  [2])|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_2  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_2  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask_5  [2])); 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_25  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[5:0]  dcache__tlb_pmp___res_hit_T_88  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit_6  =  dcache__tlb_pmp__io_pmp_cfg_a_1  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_1  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_1  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_1  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_1  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_25  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_1  [0]&~(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_0  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_0  [29:1])==29'h0&(  dcache__tlb_pmp__io_addr  [2:0]|~(  dcache__tlb_pmp___res_hit_T_88  [2:0]))<{  dcache__tlb_pmp__io_pmp_addr_0  [0],2'h0})&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_1  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_1  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_1  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore_6  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_1  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_19  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask_6  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_19  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned_6  =  dcache__tlb_pmp__io_pmp_cfg_a_1  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask_6  &~(  dcache__tlb_pmp__io_pmp_mask_1  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_0  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_0  [0]&~(  dcache__tlb_pmp__io_addr  [2])|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_1  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_1  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask_6  [2])); 
   wire[5:0]  dcache__tlb_pmp___res_hit_lsbMask_T_29  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire  dcache__tlb_pmp__res_hit_7  =  dcache__tlb_pmp__io_pmp_cfg_a_0  [1] ? ((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_0  [29:1])&~(  dcache__tlb_pmp__io_pmp_mask_0  [31:3]))==29'h0&((  dcache__tlb_pmp__io_addr  [2:0]^{  dcache__tlb_pmp__io_pmp_addr_0  [0],2'h0})&~(  dcache__tlb_pmp__io_pmp_mask_0  [2:0]|~(  dcache__tlb_pmp___res_hit_lsbMask_T_29  [2:0])))==3'h0:  dcache__tlb_pmp__io_pmp_cfg_a_0  [0]&(  dcache__tlb_pmp__io_addr  [31:3]<  dcache__tlb_pmp__io_pmp_addr_0  [29:1]|(  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_0  [29:1])==29'h0&  dcache__tlb_pmp__io_addr  [2:0]<{  dcache__tlb_pmp__io_pmp_addr_0  [0],2'h0}); 
   wire  dcache__tlb_pmp__res_ignore_7  =  dcache__tlb_pmp__io_prv  [1]&~  dcache__tlb_pmp__io_pmp_cfg_l_0  ; 
   wire[5:0]  dcache__tlb_pmp___res_aligned_lsbMask_T_22  =6'h7<<  dcache__tlb_pmp___GEN  ; 
   wire[2:0]  dcache__tlb_pmp__res_aligned_lsbMask_7  =~(  dcache__tlb_pmp___res_aligned_lsbMask_T_22  [2:0]); 
   wire  dcache__tlb_pmp__res_aligned_7  =  dcache__tlb_pmp__io_pmp_cfg_a_0  [1] ? (  dcache__tlb_pmp__res_aligned_lsbMask_7  &~(  dcache__tlb_pmp__io_pmp_mask_0  [2:0]))==3'h0:~((  dcache__tlb_pmp__io_addr  [31:3]^  dcache__tlb_pmp__io_pmp_addr_0  [29:1])==29'h0&  dcache__tlb_pmp__io_pmp_addr_0  [0]&(  dcache__tlb_pmp__io_addr  [2]|  dcache__tlb_pmp__res_aligned_lsbMask_7  [2])); 
  assign   dcache__tlb_pmp__io_r  =  dcache__tlb_pmp__res_hit_7   ?   dcache__tlb_pmp__res_aligned_7  &(  dcache__tlb_pmp__io_pmp_cfg_r_0  |  dcache__tlb_pmp__res_ignore_7  ):  dcache__tlb_pmp__res_hit_6   ?   dcache__tlb_pmp__res_aligned_6  &(  dcache__tlb_pmp__io_pmp_cfg_r_1  |  dcache__tlb_pmp__res_ignore_6  ):  dcache__tlb_pmp__res_hit_5   ?   dcache__tlb_pmp__res_aligned_5  &(  dcache__tlb_pmp__io_pmp_cfg_r_2  |  dcache__tlb_pmp__res_ignore_5  ):  dcache__tlb_pmp__res_hit_4   ?   dcache__tlb_pmp__res_aligned_4  &(  dcache__tlb_pmp__io_pmp_cfg_r_3  |  dcache__tlb_pmp__res_ignore_4  ):  dcache__tlb_pmp__res_hit_3   ?   dcache__tlb_pmp__res_aligned_3  &(  dcache__tlb_pmp__io_pmp_cfg_r_4  |  dcache__tlb_pmp__res_ignore_3  ):  dcache__tlb_pmp__res_hit_2   ?   dcache__tlb_pmp__res_aligned_2  &(  dcache__tlb_pmp__io_pmp_cfg_r_5  |  dcache__tlb_pmp__res_ignore_2  ):  dcache__tlb_pmp__res_hit_1   ?   dcache__tlb_pmp__res_aligned_1  &(  dcache__tlb_pmp__io_pmp_cfg_r_6  |  dcache__tlb_pmp__res_ignore_1  ):  dcache__tlb_pmp__res_hit   ?   dcache__tlb_pmp__res_aligned  &(  dcache__tlb_pmp__io_pmp_cfg_r_7  |  dcache__tlb_pmp__res_ignore  ):  dcache__tlb_pmp__io_prv  [1]; 
  assign   dcache__tlb_pmp__io_w  =  dcache__tlb_pmp__res_hit_7   ?   dcache__tlb_pmp__res_aligned_7  &(  dcache__tlb_pmp__io_pmp_cfg_w_0  |  dcache__tlb_pmp__res_ignore_7  ):  dcache__tlb_pmp__res_hit_6   ?   dcache__tlb_pmp__res_aligned_6  &(  dcache__tlb_pmp__io_pmp_cfg_w_1  |  dcache__tlb_pmp__res_ignore_6  ):  dcache__tlb_pmp__res_hit_5   ?   dcache__tlb_pmp__res_aligned_5  &(  dcache__tlb_pmp__io_pmp_cfg_w_2  |  dcache__tlb_pmp__res_ignore_5  ):  dcache__tlb_pmp__res_hit_4   ?   dcache__tlb_pmp__res_aligned_4  &(  dcache__tlb_pmp__io_pmp_cfg_w_3  |  dcache__tlb_pmp__res_ignore_4  ):  dcache__tlb_pmp__res_hit_3   ?   dcache__tlb_pmp__res_aligned_3  &(  dcache__tlb_pmp__io_pmp_cfg_w_4  |  dcache__tlb_pmp__res_ignore_3  ):  dcache__tlb_pmp__res_hit_2   ?   dcache__tlb_pmp__res_aligned_2  &(  dcache__tlb_pmp__io_pmp_cfg_w_5  |  dcache__tlb_pmp__res_ignore_2  ):  dcache__tlb_pmp__res_hit_1   ?   dcache__tlb_pmp__res_aligned_1  &(  dcache__tlb_pmp__io_pmp_cfg_w_6  |  dcache__tlb_pmp__res_ignore_1  ):  dcache__tlb_pmp__res_hit   ?   dcache__tlb_pmp__res_aligned  &(  dcache__tlb_pmp__io_pmp_cfg_w_7  |  dcache__tlb_pmp__res_ignore  ):  dcache__tlb_pmp__io_prv  [1];
assign dcache__tlb_pmp__io_prv = dcache__s1_tlb_req_prv;
assign dcache__tlb_pmp__io_pmp_cfg_l_0 = dcache__io_ptw_pmp_cfg_l_0;
assign dcache__tlb_pmp__io_pmp_cfg_l_1 = dcache__io_ptw_pmp_cfg_l_1;
assign dcache__tlb_pmp__io_pmp_cfg_l_2 = dcache__io_ptw_pmp_cfg_l_2;
assign dcache__tlb_pmp__io_pmp_cfg_l_3 = dcache__io_ptw_pmp_cfg_l_3;
assign dcache__tlb_pmp__io_pmp_cfg_l_4 = dcache__io_ptw_pmp_cfg_l_4;
assign dcache__tlb_pmp__io_pmp_cfg_l_5 = dcache__io_ptw_pmp_cfg_l_5;
assign dcache__tlb_pmp__io_pmp_cfg_l_6 = dcache__io_ptw_pmp_cfg_l_6;
assign dcache__tlb_pmp__io_pmp_cfg_l_7 = dcache__io_ptw_pmp_cfg_l_7;
assign dcache__tlb_pmp__io_pmp_cfg_a_0 = dcache__io_ptw_pmp_cfg_a_0;
assign dcache__tlb_pmp__io_pmp_cfg_a_1 = dcache__io_ptw_pmp_cfg_a_1;
assign dcache__tlb_pmp__io_pmp_cfg_a_2 = dcache__io_ptw_pmp_cfg_a_2;
assign dcache__tlb_pmp__io_pmp_cfg_a_3 = dcache__io_ptw_pmp_cfg_a_3;
assign dcache__tlb_pmp__io_pmp_cfg_a_4 = dcache__io_ptw_pmp_cfg_a_4;
assign dcache__tlb_pmp__io_pmp_cfg_a_5 = dcache__io_ptw_pmp_cfg_a_5;
assign dcache__tlb_pmp__io_pmp_cfg_a_6 = dcache__io_ptw_pmp_cfg_a_6;
assign dcache__tlb_pmp__io_pmp_cfg_a_7 = dcache__io_ptw_pmp_cfg_a_7;
assign dcache__tlb_pmp__io_pmp_cfg_w_0 = dcache__io_ptw_pmp_cfg_w_0;
assign dcache__tlb_pmp__io_pmp_cfg_w_1 = dcache__io_ptw_pmp_cfg_w_1;
assign dcache__tlb_pmp__io_pmp_cfg_w_2 = dcache__io_ptw_pmp_cfg_w_2;
assign dcache__tlb_pmp__io_pmp_cfg_w_3 = dcache__io_ptw_pmp_cfg_w_3;
assign dcache__tlb_pmp__io_pmp_cfg_w_4 = dcache__io_ptw_pmp_cfg_w_4;
assign dcache__tlb_pmp__io_pmp_cfg_w_5 = dcache__io_ptw_pmp_cfg_w_5;
assign dcache__tlb_pmp__io_pmp_cfg_w_6 = dcache__io_ptw_pmp_cfg_w_6;
assign dcache__tlb_pmp__io_pmp_cfg_w_7 = dcache__io_ptw_pmp_cfg_w_7;
assign dcache__tlb_pmp__io_pmp_cfg_r_0 = dcache__io_ptw_pmp_cfg_r_0;
assign dcache__tlb_pmp__io_pmp_cfg_r_1 = dcache__io_ptw_pmp_cfg_r_1;
assign dcache__tlb_pmp__io_pmp_cfg_r_2 = dcache__io_ptw_pmp_cfg_r_2;
assign dcache__tlb_pmp__io_pmp_cfg_r_3 = dcache__io_ptw_pmp_cfg_r_3;
assign dcache__tlb_pmp__io_pmp_cfg_r_4 = dcache__io_ptw_pmp_cfg_r_4;
assign dcache__tlb_pmp__io_pmp_cfg_r_5 = dcache__io_ptw_pmp_cfg_r_5;
assign dcache__tlb_pmp__io_pmp_cfg_r_6 = dcache__io_ptw_pmp_cfg_r_6;
assign dcache__tlb_pmp__io_pmp_cfg_r_7 = dcache__io_ptw_pmp_cfg_r_7;
assign dcache__tlb_pmp__io_pmp_addr_0 = dcache__io_ptw_pmp_addr_0;
assign dcache__tlb_pmp__io_pmp_addr_1 = dcache__io_ptw_pmp_addr_1;
assign dcache__tlb_pmp__io_pmp_addr_2 = dcache__io_ptw_pmp_addr_2;
assign dcache__tlb_pmp__io_pmp_addr_3 = dcache__io_ptw_pmp_addr_3;
assign dcache__tlb_pmp__io_pmp_addr_4 = dcache__io_ptw_pmp_addr_4;
assign dcache__tlb_pmp__io_pmp_addr_5 = dcache__io_ptw_pmp_addr_5;
assign dcache__tlb_pmp__io_pmp_addr_6 = dcache__io_ptw_pmp_addr_6;
assign dcache__tlb_pmp__io_pmp_addr_7 = dcache__io_ptw_pmp_addr_7;
assign dcache__tlb_pmp__io_pmp_mask_0 = dcache__io_ptw_pmp_mask_0;
assign dcache__tlb_pmp__io_pmp_mask_1 = dcache__io_ptw_pmp_mask_1;
assign dcache__tlb_pmp__io_pmp_mask_2 = dcache__io_ptw_pmp_mask_2;
assign dcache__tlb_pmp__io_pmp_mask_3 = dcache__io_ptw_pmp_mask_3;
assign dcache__tlb_pmp__io_pmp_mask_4 = dcache__io_ptw_pmp_mask_4;
assign dcache__tlb_pmp__io_pmp_mask_5 = dcache__io_ptw_pmp_mask_5;
assign dcache__tlb_pmp__io_pmp_mask_6 = dcache__io_ptw_pmp_mask_6;
assign dcache__tlb_pmp__io_pmp_mask_7 = dcache__io_ptw_pmp_mask_7;
assign dcache__tlb_pmp__io_addr = dcache__s1_tlb_req_vaddr[31:0];
assign dcache__tlb_pmp__io_size = dcache__s1_tlb_req_size;
assign dcache___tlb_pmp_io_r = dcache__tlb_pmp__io_r;
assign dcache___tlb_pmp_io_w = dcache__tlb_pmp__io_w;
  
  
wire  dcache__tlb_entries_barrier__io_x_u;
wire  dcache__tlb_entries_barrier__io_x_ae_ptw;
wire  dcache__tlb_entries_barrier__io_x_ae_final;
wire  dcache__tlb_entries_barrier__io_x_pf;
wire  dcache__tlb_entries_barrier__io_x_gf;
wire  dcache__tlb_entries_barrier__io_x_sw;
wire  dcache__tlb_entries_barrier__io_x_sx;
wire  dcache__tlb_entries_barrier__io_x_sr;
wire  dcache__tlb_entries_barrier__io_x_pw;
wire  dcache__tlb_entries_barrier__io_x_px;
wire  dcache__tlb_entries_barrier__io_x_pr;
wire  dcache__tlb_entries_barrier__io_x_ppp;
wire  dcache__tlb_entries_barrier__io_x_pal;
wire  dcache__tlb_entries_barrier__io_x_paa;
wire  dcache__tlb_entries_barrier__io_x_eff;
wire  dcache__tlb_entries_barrier__io_x_c;
wire  dcache__tlb_entries_barrier__io_y_u;
wire  dcache__tlb_entries_barrier__io_y_ae_ptw;
wire  dcache__tlb_entries_barrier__io_y_ae_final;
wire  dcache__tlb_entries_barrier__io_y_pf;
wire  dcache__tlb_entries_barrier__io_y_gf;
wire  dcache__tlb_entries_barrier__io_y_sw;
wire  dcache__tlb_entries_barrier__io_y_sx;
wire  dcache__tlb_entries_barrier__io_y_sr;
wire  dcache__tlb_entries_barrier__io_y_pw;
wire  dcache__tlb_entries_barrier__io_y_px;
wire  dcache__tlb_entries_barrier__io_y_pr;
wire  dcache__tlb_entries_barrier__io_y_ppp;
wire  dcache__tlb_entries_barrier__io_y_pal;
wire  dcache__tlb_entries_barrier__io_y_paa;
wire  dcache__tlb_entries_barrier__io_y_eff;
wire  dcache__tlb_entries_barrier__io_y_c;
wire  dcache__tlb_entries_barrier_1__io_x_u;
wire  dcache__tlb_entries_barrier_1__io_x_ae_ptw;
wire  dcache__tlb_entries_barrier_1__io_x_ae_final;
wire  dcache__tlb_entries_barrier_1__io_x_pf;
wire  dcache__tlb_entries_barrier_1__io_x_gf;
wire  dcache__tlb_entries_barrier_1__io_x_sw;
wire  dcache__tlb_entries_barrier_1__io_x_sx;
wire  dcache__tlb_entries_barrier_1__io_x_sr;
wire  dcache__tlb_entries_barrier_1__io_x_pw;
wire  dcache__tlb_entries_barrier_1__io_x_px;
wire  dcache__tlb_entries_barrier_1__io_x_pr;
wire  dcache__tlb_entries_barrier_1__io_x_ppp;
wire  dcache__tlb_entries_barrier_1__io_x_pal;
wire  dcache__tlb_entries_barrier_1__io_x_paa;
wire  dcache__tlb_entries_barrier_1__io_x_eff;
wire  dcache__tlb_entries_barrier_1__io_x_c;
wire  dcache__tlb_entries_barrier_1__io_y_u;
wire  dcache__tlb_entries_barrier_1__io_y_ae_ptw;
wire  dcache__tlb_entries_barrier_1__io_y_ae_final;
wire  dcache__tlb_entries_barrier_1__io_y_pf;
wire  dcache__tlb_entries_barrier_1__io_y_gf;
wire  dcache__tlb_entries_barrier_1__io_y_sw;
wire  dcache__tlb_entries_barrier_1__io_y_sx;
wire  dcache__tlb_entries_barrier_1__io_y_sr;
wire  dcache__tlb_entries_barrier_1__io_y_pw;
wire  dcache__tlb_entries_barrier_1__io_y_px;
wire  dcache__tlb_entries_barrier_1__io_y_pr;
wire  dcache__tlb_entries_barrier_1__io_y_ppp;
wire  dcache__tlb_entries_barrier_1__io_y_pal;
wire  dcache__tlb_entries_barrier_1__io_y_paa;
wire  dcache__tlb_entries_barrier_1__io_y_eff;
wire  dcache__tlb_entries_barrier_1__io_y_c;
wire  dcache__tlb_entries_barrier_2__io_x_u;
wire  dcache__tlb_entries_barrier_2__io_x_ae_ptw;
wire  dcache__tlb_entries_barrier_2__io_x_ae_final;
wire  dcache__tlb_entries_barrier_2__io_x_pf;
wire  dcache__tlb_entries_barrier_2__io_x_gf;
wire  dcache__tlb_entries_barrier_2__io_x_sw;
wire  dcache__tlb_entries_barrier_2__io_x_sx;
wire  dcache__tlb_entries_barrier_2__io_x_sr;
wire  dcache__tlb_entries_barrier_2__io_x_pw;
wire  dcache__tlb_entries_barrier_2__io_x_px;
wire  dcache__tlb_entries_barrier_2__io_x_pr;
wire  dcache__tlb_entries_barrier_2__io_x_ppp;
wire  dcache__tlb_entries_barrier_2__io_x_pal;
wire  dcache__tlb_entries_barrier_2__io_x_paa;
wire  dcache__tlb_entries_barrier_2__io_x_eff;
wire  dcache__tlb_entries_barrier_2__io_x_c;
wire  dcache__tlb_entries_barrier_2__io_y_u;
wire  dcache__tlb_entries_barrier_2__io_y_ae_ptw;
wire  dcache__tlb_entries_barrier_2__io_y_ae_final;
wire  dcache__tlb_entries_barrier_2__io_y_pf;
wire  dcache__tlb_entries_barrier_2__io_y_gf;
wire  dcache__tlb_entries_barrier_2__io_y_sw;
wire  dcache__tlb_entries_barrier_2__io_y_sx;
wire  dcache__tlb_entries_barrier_2__io_y_sr;
wire  dcache__tlb_entries_barrier_2__io_y_pw;
wire  dcache__tlb_entries_barrier_2__io_y_px;
wire  dcache__tlb_entries_barrier_2__io_y_pr;
wire  dcache__tlb_entries_barrier_2__io_y_ppp;
wire  dcache__tlb_entries_barrier_2__io_y_pal;
wire  dcache__tlb_entries_barrier_2__io_y_paa;
wire  dcache__tlb_entries_barrier_2__io_y_eff;
wire  dcache__tlb_entries_barrier_2__io_y_c;
wire  dcache__tlb_entries_barrier_3__io_x_u;
wire  dcache__tlb_entries_barrier_3__io_x_ae_ptw;
wire  dcache__tlb_entries_barrier_3__io_x_ae_final;
wire  dcache__tlb_entries_barrier_3__io_x_pf;
wire  dcache__tlb_entries_barrier_3__io_x_gf;
wire  dcache__tlb_entries_barrier_3__io_x_sw;
wire  dcache__tlb_entries_barrier_3__io_x_sx;
wire  dcache__tlb_entries_barrier_3__io_x_sr;
wire  dcache__tlb_entries_barrier_3__io_x_pw;
wire  dcache__tlb_entries_barrier_3__io_x_px;
wire  dcache__tlb_entries_barrier_3__io_x_pr;
wire  dcache__tlb_entries_barrier_3__io_x_ppp;
wire  dcache__tlb_entries_barrier_3__io_x_pal;
wire  dcache__tlb_entries_barrier_3__io_x_paa;
wire  dcache__tlb_entries_barrier_3__io_x_eff;
wire  dcache__tlb_entries_barrier_3__io_x_c;
wire  dcache__tlb_entries_barrier_3__io_y_u;
wire  dcache__tlb_entries_barrier_3__io_y_ae_ptw;
wire  dcache__tlb_entries_barrier_3__io_y_ae_final;
wire  dcache__tlb_entries_barrier_3__io_y_pf;
wire  dcache__tlb_entries_barrier_3__io_y_gf;
wire  dcache__tlb_entries_barrier_3__io_y_sw;
wire  dcache__tlb_entries_barrier_3__io_y_sx;
wire  dcache__tlb_entries_barrier_3__io_y_sr;
wire  dcache__tlb_entries_barrier_3__io_y_pw;
wire  dcache__tlb_entries_barrier_3__io_y_px;
wire  dcache__tlb_entries_barrier_3__io_y_pr;
wire  dcache__tlb_entries_barrier_3__io_y_ppp;
wire  dcache__tlb_entries_barrier_3__io_y_pal;
wire  dcache__tlb_entries_barrier_3__io_y_paa;
wire  dcache__tlb_entries_barrier_3__io_y_eff;
wire  dcache__tlb_entries_barrier_3__io_y_c;
wire  dcache__tlb_entries_barrier_4__io_x_u;
wire  dcache__tlb_entries_barrier_4__io_x_ae_ptw;
wire  dcache__tlb_entries_barrier_4__io_x_ae_final;
wire  dcache__tlb_entries_barrier_4__io_x_pf;
wire  dcache__tlb_entries_barrier_4__io_x_gf;
wire  dcache__tlb_entries_barrier_4__io_x_sw;
wire  dcache__tlb_entries_barrier_4__io_x_sx;
wire  dcache__tlb_entries_barrier_4__io_x_sr;
wire  dcache__tlb_entries_barrier_4__io_x_pw;
wire  dcache__tlb_entries_barrier_4__io_x_px;
wire  dcache__tlb_entries_barrier_4__io_x_pr;
wire  dcache__tlb_entries_barrier_4__io_x_ppp;
wire  dcache__tlb_entries_barrier_4__io_x_pal;
wire  dcache__tlb_entries_barrier_4__io_x_paa;
wire  dcache__tlb_entries_barrier_4__io_x_eff;
wire  dcache__tlb_entries_barrier_4__io_x_c;
wire  dcache__tlb_entries_barrier_4__io_y_u;
wire  dcache__tlb_entries_barrier_4__io_y_ae_ptw;
wire  dcache__tlb_entries_barrier_4__io_y_ae_final;
wire  dcache__tlb_entries_barrier_4__io_y_pf;
wire  dcache__tlb_entries_barrier_4__io_y_gf;
wire  dcache__tlb_entries_barrier_4__io_y_sw;
wire  dcache__tlb_entries_barrier_4__io_y_sx;
wire  dcache__tlb_entries_barrier_4__io_y_sr;
wire  dcache__tlb_entries_barrier_4__io_y_pw;
wire  dcache__tlb_entries_barrier_4__io_y_px;
wire  dcache__tlb_entries_barrier_4__io_y_pr;
wire  dcache__tlb_entries_barrier_4__io_y_ppp;
wire  dcache__tlb_entries_barrier_4__io_y_pal;
wire  dcache__tlb_entries_barrier_4__io_y_paa;
wire  dcache__tlb_entries_barrier_4__io_y_eff;
wire  dcache__tlb_entries_barrier_4__io_y_c;
wire  dcache__tlb_entries_barrier_5__io_x_u;
wire  dcache__tlb_entries_barrier_5__io_x_ae_ptw;
wire  dcache__tlb_entries_barrier_5__io_x_ae_final;
wire  dcache__tlb_entries_barrier_5__io_x_pf;
wire  dcache__tlb_entries_barrier_5__io_x_gf;
wire  dcache__tlb_entries_barrier_5__io_x_sw;
wire  dcache__tlb_entries_barrier_5__io_x_sx;
wire  dcache__tlb_entries_barrier_5__io_x_sr;
wire  dcache__tlb_entries_barrier_5__io_x_pw;
wire  dcache__tlb_entries_barrier_5__io_x_px;
wire  dcache__tlb_entries_barrier_5__io_x_pr;
wire  dcache__tlb_entries_barrier_5__io_x_ppp;
wire  dcache__tlb_entries_barrier_5__io_x_pal;
wire  dcache__tlb_entries_barrier_5__io_x_paa;
wire  dcache__tlb_entries_barrier_5__io_x_eff;
wire  dcache__tlb_entries_barrier_5__io_x_c;
wire  dcache__tlb_entries_barrier_5__io_y_u;
wire  dcache__tlb_entries_barrier_5__io_y_ae_ptw;
wire  dcache__tlb_entries_barrier_5__io_y_ae_final;
wire  dcache__tlb_entries_barrier_5__io_y_pf;
wire  dcache__tlb_entries_barrier_5__io_y_gf;
wire  dcache__tlb_entries_barrier_5__io_y_sw;
wire  dcache__tlb_entries_barrier_5__io_y_sx;
wire  dcache__tlb_entries_barrier_5__io_y_sr;
wire  dcache__tlb_entries_barrier_5__io_y_pw;
wire  dcache__tlb_entries_barrier_5__io_y_px;
wire  dcache__tlb_entries_barrier_5__io_y_pr;
wire  dcache__tlb_entries_barrier_5__io_y_ppp;
wire  dcache__tlb_entries_barrier_5__io_y_pal;
wire  dcache__tlb_entries_barrier_5__io_y_paa;
wire  dcache__tlb_entries_barrier_5__io_y_eff;
wire  dcache__tlb_entries_barrier_5__io_y_c;
wire  dcache__pma_checker_entries_barrier__io_x_u;
wire  dcache__pma_checker_entries_barrier__io_x_ae_ptw;
wire  dcache__pma_checker_entries_barrier__io_x_ae_final;
wire  dcache__pma_checker_entries_barrier__io_x_pf;
wire  dcache__pma_checker_entries_barrier__io_x_gf;
wire  dcache__pma_checker_entries_barrier__io_x_sw;
wire  dcache__pma_checker_entries_barrier__io_x_sx;
wire  dcache__pma_checker_entries_barrier__io_x_sr;
wire  dcache__pma_checker_entries_barrier__io_x_pw;
wire  dcache__pma_checker_entries_barrier__io_x_px;
wire  dcache__pma_checker_entries_barrier__io_x_pr;
wire  dcache__pma_checker_entries_barrier__io_x_ppp;
wire  dcache__pma_checker_entries_barrier__io_x_pal;
wire  dcache__pma_checker_entries_barrier__io_x_paa;
wire  dcache__pma_checker_entries_barrier__io_x_eff;
wire  dcache__pma_checker_entries_barrier__io_x_c;
wire  dcache__pma_checker_entries_barrier__io_y_u;
wire  dcache__pma_checker_entries_barrier__io_y_ae_ptw;
wire  dcache__pma_checker_entries_barrier__io_y_ae_final;
wire  dcache__pma_checker_entries_barrier__io_y_pf;
wire  dcache__pma_checker_entries_barrier__io_y_gf;
wire  dcache__pma_checker_entries_barrier__io_y_sw;
wire  dcache__pma_checker_entries_barrier__io_y_sx;
wire  dcache__pma_checker_entries_barrier__io_y_sr;
wire  dcache__pma_checker_entries_barrier__io_y_pw;
wire  dcache__pma_checker_entries_barrier__io_y_px;
wire  dcache__pma_checker_entries_barrier__io_y_pr;
wire  dcache__pma_checker_entries_barrier__io_y_ppp;
wire  dcache__pma_checker_entries_barrier__io_y_pal;
wire  dcache__pma_checker_entries_barrier__io_y_paa;
wire  dcache__pma_checker_entries_barrier__io_y_eff;
wire  dcache__pma_checker_entries_barrier__io_y_c;
wire  dcache__pma_checker_entries_barrier_1__io_x_u;
wire  dcache__pma_checker_entries_barrier_1__io_x_ae_ptw;
wire  dcache__pma_checker_entries_barrier_1__io_x_ae_final;
wire  dcache__pma_checker_entries_barrier_1__io_x_pf;
wire  dcache__pma_checker_entries_barrier_1__io_x_gf;
wire  dcache__pma_checker_entries_barrier_1__io_x_sw;
wire  dcache__pma_checker_entries_barrier_1__io_x_sx;
wire  dcache__pma_checker_entries_barrier_1__io_x_sr;
wire  dcache__pma_checker_entries_barrier_1__io_x_pw;
wire  dcache__pma_checker_entries_barrier_1__io_x_px;
wire  dcache__pma_checker_entries_barrier_1__io_x_pr;
wire  dcache__pma_checker_entries_barrier_1__io_x_ppp;
wire  dcache__pma_checker_entries_barrier_1__io_x_pal;
wire  dcache__pma_checker_entries_barrier_1__io_x_paa;
wire  dcache__pma_checker_entries_barrier_1__io_x_eff;
wire  dcache__pma_checker_entries_barrier_1__io_x_c;
wire  dcache__pma_checker_entries_barrier_1__io_y_u;
wire  dcache__pma_checker_entries_barrier_1__io_y_ae_ptw;
wire  dcache__pma_checker_entries_barrier_1__io_y_ae_final;
wire  dcache__pma_checker_entries_barrier_1__io_y_pf;
wire  dcache__pma_checker_entries_barrier_1__io_y_gf;
wire  dcache__pma_checker_entries_barrier_1__io_y_sw;
wire  dcache__pma_checker_entries_barrier_1__io_y_sx;
wire  dcache__pma_checker_entries_barrier_1__io_y_sr;
wire  dcache__pma_checker_entries_barrier_1__io_y_pw;
wire  dcache__pma_checker_entries_barrier_1__io_y_px;
wire  dcache__pma_checker_entries_barrier_1__io_y_pr;
wire  dcache__pma_checker_entries_barrier_1__io_y_ppp;
wire  dcache__pma_checker_entries_barrier_1__io_y_pal;
wire  dcache__pma_checker_entries_barrier_1__io_y_paa;
wire  dcache__pma_checker_entries_barrier_1__io_y_eff;
wire  dcache__pma_checker_entries_barrier_1__io_y_c;
wire  dcache__pma_checker_entries_barrier_2__io_x_u;
wire  dcache__pma_checker_entries_barrier_2__io_x_ae_ptw;
wire  dcache__pma_checker_entries_barrier_2__io_x_ae_final;
wire  dcache__pma_checker_entries_barrier_2__io_x_pf;
wire  dcache__pma_checker_entries_barrier_2__io_x_gf;
wire  dcache__pma_checker_entries_barrier_2__io_x_sw;
wire  dcache__pma_checker_entries_barrier_2__io_x_sx;
wire  dcache__pma_checker_entries_barrier_2__io_x_sr;
wire  dcache__pma_checker_entries_barrier_2__io_x_pw;
wire  dcache__pma_checker_entries_barrier_2__io_x_px;
wire  dcache__pma_checker_entries_barrier_2__io_x_pr;
wire  dcache__pma_checker_entries_barrier_2__io_x_ppp;
wire  dcache__pma_checker_entries_barrier_2__io_x_pal;
wire  dcache__pma_checker_entries_barrier_2__io_x_paa;
wire  dcache__pma_checker_entries_barrier_2__io_x_eff;
wire  dcache__pma_checker_entries_barrier_2__io_x_c;
wire  dcache__pma_checker_entries_barrier_2__io_y_u;
wire  dcache__pma_checker_entries_barrier_2__io_y_ae_ptw;
wire  dcache__pma_checker_entries_barrier_2__io_y_ae_final;
wire  dcache__pma_checker_entries_barrier_2__io_y_pf;
wire  dcache__pma_checker_entries_barrier_2__io_y_gf;
wire  dcache__pma_checker_entries_barrier_2__io_y_sw;
wire  dcache__pma_checker_entries_barrier_2__io_y_sx;
wire  dcache__pma_checker_entries_barrier_2__io_y_sr;
wire  dcache__pma_checker_entries_barrier_2__io_y_pw;
wire  dcache__pma_checker_entries_barrier_2__io_y_px;
wire  dcache__pma_checker_entries_barrier_2__io_y_pr;
wire  dcache__pma_checker_entries_barrier_2__io_y_ppp;
wire  dcache__pma_checker_entries_barrier_2__io_y_pal;
wire  dcache__pma_checker_entries_barrier_2__io_y_paa;
wire  dcache__pma_checker_entries_barrier_2__io_y_eff;
wire  dcache__pma_checker_entries_barrier_2__io_y_c;
wire  dcache__pma_checker_entries_barrier_3__io_x_u;
wire  dcache__pma_checker_entries_barrier_3__io_x_ae_ptw;
wire  dcache__pma_checker_entries_barrier_3__io_x_ae_final;
wire  dcache__pma_checker_entries_barrier_3__io_x_pf;
wire  dcache__pma_checker_entries_barrier_3__io_x_gf;
wire  dcache__pma_checker_entries_barrier_3__io_x_sw;
wire  dcache__pma_checker_entries_barrier_3__io_x_sx;
wire  dcache__pma_checker_entries_barrier_3__io_x_sr;
wire  dcache__pma_checker_entries_barrier_3__io_x_pw;
wire  dcache__pma_checker_entries_barrier_3__io_x_px;
wire  dcache__pma_checker_entries_barrier_3__io_x_pr;
wire  dcache__pma_checker_entries_barrier_3__io_x_ppp;
wire  dcache__pma_checker_entries_barrier_3__io_x_pal;
wire  dcache__pma_checker_entries_barrier_3__io_x_paa;
wire  dcache__pma_checker_entries_barrier_3__io_x_eff;
wire  dcache__pma_checker_entries_barrier_3__io_x_c;
wire  dcache__pma_checker_entries_barrier_3__io_y_u;
wire  dcache__pma_checker_entries_barrier_3__io_y_ae_ptw;
wire  dcache__pma_checker_entries_barrier_3__io_y_ae_final;
wire  dcache__pma_checker_entries_barrier_3__io_y_pf;
wire  dcache__pma_checker_entries_barrier_3__io_y_gf;
wire  dcache__pma_checker_entries_barrier_3__io_y_sw;
wire  dcache__pma_checker_entries_barrier_3__io_y_sx;
wire  dcache__pma_checker_entries_barrier_3__io_y_sr;
wire  dcache__pma_checker_entries_barrier_3__io_y_pw;
wire  dcache__pma_checker_entries_barrier_3__io_y_px;
wire  dcache__pma_checker_entries_barrier_3__io_y_pr;
wire  dcache__pma_checker_entries_barrier_3__io_y_ppp;
wire  dcache__pma_checker_entries_barrier_3__io_y_pal;
wire  dcache__pma_checker_entries_barrier_3__io_y_paa;
wire  dcache__pma_checker_entries_barrier_3__io_y_eff;
wire  dcache__pma_checker_entries_barrier_3__io_y_c;
wire  dcache__pma_checker_entries_barrier_4__io_x_u;
wire  dcache__pma_checker_entries_barrier_4__io_x_ae_ptw;
wire  dcache__pma_checker_entries_barrier_4__io_x_ae_final;
wire  dcache__pma_checker_entries_barrier_4__io_x_pf;
wire  dcache__pma_checker_entries_barrier_4__io_x_gf;
wire  dcache__pma_checker_entries_barrier_4__io_x_sw;
wire  dcache__pma_checker_entries_barrier_4__io_x_sx;
wire  dcache__pma_checker_entries_barrier_4__io_x_sr;
wire  dcache__pma_checker_entries_barrier_4__io_x_pw;
wire  dcache__pma_checker_entries_barrier_4__io_x_px;
wire  dcache__pma_checker_entries_barrier_4__io_x_pr;
wire  dcache__pma_checker_entries_barrier_4__io_x_ppp;
wire  dcache__pma_checker_entries_barrier_4__io_x_pal;
wire  dcache__pma_checker_entries_barrier_4__io_x_paa;
wire  dcache__pma_checker_entries_barrier_4__io_x_eff;
wire  dcache__pma_checker_entries_barrier_4__io_x_c;
wire  dcache__pma_checker_entries_barrier_4__io_y_u;
wire  dcache__pma_checker_entries_barrier_4__io_y_ae_ptw;
wire  dcache__pma_checker_entries_barrier_4__io_y_ae_final;
wire  dcache__pma_checker_entries_barrier_4__io_y_pf;
wire  dcache__pma_checker_entries_barrier_4__io_y_gf;
wire  dcache__pma_checker_entries_barrier_4__io_y_sw;
wire  dcache__pma_checker_entries_barrier_4__io_y_sx;
wire  dcache__pma_checker_entries_barrier_4__io_y_sr;
wire  dcache__pma_checker_entries_barrier_4__io_y_pw;
wire  dcache__pma_checker_entries_barrier_4__io_y_px;
wire  dcache__pma_checker_entries_barrier_4__io_y_pr;
wire  dcache__pma_checker_entries_barrier_4__io_y_ppp;
wire  dcache__pma_checker_entries_barrier_4__io_y_pal;
wire  dcache__pma_checker_entries_barrier_4__io_y_paa;
wire  dcache__pma_checker_entries_barrier_4__io_y_eff;
wire  dcache__pma_checker_entries_barrier_4__io_y_c;
 
  assign   dcache__tlb_entries_barrier__io_y_u  =  dcache__tlb_entries_barrier__io_x_u  ; 
  assign   dcache__tlb_entries_barrier__io_y_ae_ptw  =  dcache__tlb_entries_barrier__io_x_ae_ptw  ; 
  assign   dcache__tlb_entries_barrier__io_y_ae_final  =  dcache__tlb_entries_barrier__io_x_ae_final  ; 
  assign   dcache__tlb_entries_barrier__io_y_pf  =  dcache__tlb_entries_barrier__io_x_pf  ; 
  assign   dcache__tlb_entries_barrier__io_y_gf  =  dcache__tlb_entries_barrier__io_x_gf  ; 
  assign   dcache__tlb_entries_barrier__io_y_sw  =  dcache__tlb_entries_barrier__io_x_sw  ; 
  assign   dcache__tlb_entries_barrier__io_y_sx  =  dcache__tlb_entries_barrier__io_x_sx  ; 
  assign   dcache__tlb_entries_barrier__io_y_sr  =  dcache__tlb_entries_barrier__io_x_sr  ; 
  assign   dcache__tlb_entries_barrier__io_y_pw  =  dcache__tlb_entries_barrier__io_x_pw  ; 
  assign   dcache__tlb_entries_barrier__io_y_px  =  dcache__tlb_entries_barrier__io_x_px  ; 
  assign   dcache__tlb_entries_barrier__io_y_pr  =  dcache__tlb_entries_barrier__io_x_pr  ; 
  assign   dcache__tlb_entries_barrier__io_y_ppp  =  dcache__tlb_entries_barrier__io_x_ppp  ; 
  assign   dcache__tlb_entries_barrier__io_y_pal  =  dcache__tlb_entries_barrier__io_x_pal  ; 
  assign   dcache__tlb_entries_barrier__io_y_paa  =  dcache__tlb_entries_barrier__io_x_paa  ; 
  assign   dcache__tlb_entries_barrier__io_y_eff  =  dcache__tlb_entries_barrier__io_x_eff  ; 
  assign   dcache__tlb_entries_barrier__io_y_c  =  dcache__tlb_entries_barrier__io_x_c  ;
  
  
 
  assign   dcache__tlb_entries_barrier_1__io_y_u  =  dcache__tlb_entries_barrier_1__io_x_u  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_ae_ptw  =  dcache__tlb_entries_barrier_1__io_x_ae_ptw  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_ae_final  =  dcache__tlb_entries_barrier_1__io_x_ae_final  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_pf  =  dcache__tlb_entries_barrier_1__io_x_pf  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_gf  =  dcache__tlb_entries_barrier_1__io_x_gf  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_sw  =  dcache__tlb_entries_barrier_1__io_x_sw  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_sx  =  dcache__tlb_entries_barrier_1__io_x_sx  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_sr  =  dcache__tlb_entries_barrier_1__io_x_sr  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_pw  =  dcache__tlb_entries_barrier_1__io_x_pw  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_px  =  dcache__tlb_entries_barrier_1__io_x_px  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_pr  =  dcache__tlb_entries_barrier_1__io_x_pr  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_ppp  =  dcache__tlb_entries_barrier_1__io_x_ppp  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_pal  =  dcache__tlb_entries_barrier_1__io_x_pal  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_paa  =  dcache__tlb_entries_barrier_1__io_x_paa  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_eff  =  dcache__tlb_entries_barrier_1__io_x_eff  ; 
  assign   dcache__tlb_entries_barrier_1__io_y_c  =  dcache__tlb_entries_barrier_1__io_x_c  ;
  
  
 
  assign   dcache__tlb_entries_barrier_2__io_y_u  =  dcache__tlb_entries_barrier_2__io_x_u  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_ae_ptw  =  dcache__tlb_entries_barrier_2__io_x_ae_ptw  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_ae_final  =  dcache__tlb_entries_barrier_2__io_x_ae_final  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_pf  =  dcache__tlb_entries_barrier_2__io_x_pf  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_gf  =  dcache__tlb_entries_barrier_2__io_x_gf  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_sw  =  dcache__tlb_entries_barrier_2__io_x_sw  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_sx  =  dcache__tlb_entries_barrier_2__io_x_sx  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_sr  =  dcache__tlb_entries_barrier_2__io_x_sr  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_pw  =  dcache__tlb_entries_barrier_2__io_x_pw  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_px  =  dcache__tlb_entries_barrier_2__io_x_px  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_pr  =  dcache__tlb_entries_barrier_2__io_x_pr  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_ppp  =  dcache__tlb_entries_barrier_2__io_x_ppp  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_pal  =  dcache__tlb_entries_barrier_2__io_x_pal  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_paa  =  dcache__tlb_entries_barrier_2__io_x_paa  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_eff  =  dcache__tlb_entries_barrier_2__io_x_eff  ; 
  assign   dcache__tlb_entries_barrier_2__io_y_c  =  dcache__tlb_entries_barrier_2__io_x_c  ;
  
  
 
  assign   dcache__tlb_entries_barrier_3__io_y_u  =  dcache__tlb_entries_barrier_3__io_x_u  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_ae_ptw  =  dcache__tlb_entries_barrier_3__io_x_ae_ptw  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_ae_final  =  dcache__tlb_entries_barrier_3__io_x_ae_final  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_pf  =  dcache__tlb_entries_barrier_3__io_x_pf  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_gf  =  dcache__tlb_entries_barrier_3__io_x_gf  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_sw  =  dcache__tlb_entries_barrier_3__io_x_sw  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_sx  =  dcache__tlb_entries_barrier_3__io_x_sx  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_sr  =  dcache__tlb_entries_barrier_3__io_x_sr  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_pw  =  dcache__tlb_entries_barrier_3__io_x_pw  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_px  =  dcache__tlb_entries_barrier_3__io_x_px  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_pr  =  dcache__tlb_entries_barrier_3__io_x_pr  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_ppp  =  dcache__tlb_entries_barrier_3__io_x_ppp  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_pal  =  dcache__tlb_entries_barrier_3__io_x_pal  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_paa  =  dcache__tlb_entries_barrier_3__io_x_paa  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_eff  =  dcache__tlb_entries_barrier_3__io_x_eff  ; 
  assign   dcache__tlb_entries_barrier_3__io_y_c  =  dcache__tlb_entries_barrier_3__io_x_c  ;
  
  
 
  assign   dcache__tlb_entries_barrier_4__io_y_u  =  dcache__tlb_entries_barrier_4__io_x_u  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_ae_ptw  =  dcache__tlb_entries_barrier_4__io_x_ae_ptw  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_ae_final  =  dcache__tlb_entries_barrier_4__io_x_ae_final  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_pf  =  dcache__tlb_entries_barrier_4__io_x_pf  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_gf  =  dcache__tlb_entries_barrier_4__io_x_gf  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_sw  =  dcache__tlb_entries_barrier_4__io_x_sw  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_sx  =  dcache__tlb_entries_barrier_4__io_x_sx  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_sr  =  dcache__tlb_entries_barrier_4__io_x_sr  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_pw  =  dcache__tlb_entries_barrier_4__io_x_pw  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_px  =  dcache__tlb_entries_barrier_4__io_x_px  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_pr  =  dcache__tlb_entries_barrier_4__io_x_pr  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_ppp  =  dcache__tlb_entries_barrier_4__io_x_ppp  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_pal  =  dcache__tlb_entries_barrier_4__io_x_pal  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_paa  =  dcache__tlb_entries_barrier_4__io_x_paa  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_eff  =  dcache__tlb_entries_barrier_4__io_x_eff  ; 
  assign   dcache__tlb_entries_barrier_4__io_y_c  =  dcache__tlb_entries_barrier_4__io_x_c  ;
  
  
 
  assign   dcache__tlb_entries_barrier_5__io_y_u  =  dcache__tlb_entries_barrier_5__io_x_u  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_ae_ptw  =  dcache__tlb_entries_barrier_5__io_x_ae_ptw  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_ae_final  =  dcache__tlb_entries_barrier_5__io_x_ae_final  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_pf  =  dcache__tlb_entries_barrier_5__io_x_pf  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_gf  =  dcache__tlb_entries_barrier_5__io_x_gf  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_sw  =  dcache__tlb_entries_barrier_5__io_x_sw  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_sx  =  dcache__tlb_entries_barrier_5__io_x_sx  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_sr  =  dcache__tlb_entries_barrier_5__io_x_sr  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_pw  =  dcache__tlb_entries_barrier_5__io_x_pw  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_px  =  dcache__tlb_entries_barrier_5__io_x_px  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_pr  =  dcache__tlb_entries_barrier_5__io_x_pr  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_ppp  =  dcache__tlb_entries_barrier_5__io_x_ppp  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_pal  =  dcache__tlb_entries_barrier_5__io_x_pal  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_paa  =  dcache__tlb_entries_barrier_5__io_x_paa  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_eff  =  dcache__tlb_entries_barrier_5__io_x_eff  ; 
  assign   dcache__tlb_entries_barrier_5__io_y_c  =  dcache__tlb_entries_barrier_5__io_x_c  ;
  
  
 
  assign   dcache__pma_checker_entries_barrier__io_y_u  =  dcache__pma_checker_entries_barrier__io_x_u  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_ae_ptw  =  dcache__pma_checker_entries_barrier__io_x_ae_ptw  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_ae_final  =  dcache__pma_checker_entries_barrier__io_x_ae_final  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_pf  =  dcache__pma_checker_entries_barrier__io_x_pf  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_gf  =  dcache__pma_checker_entries_barrier__io_x_gf  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_sw  =  dcache__pma_checker_entries_barrier__io_x_sw  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_sx  =  dcache__pma_checker_entries_barrier__io_x_sx  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_sr  =  dcache__pma_checker_entries_barrier__io_x_sr  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_pw  =  dcache__pma_checker_entries_barrier__io_x_pw  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_px  =  dcache__pma_checker_entries_barrier__io_x_px  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_pr  =  dcache__pma_checker_entries_barrier__io_x_pr  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_ppp  =  dcache__pma_checker_entries_barrier__io_x_ppp  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_pal  =  dcache__pma_checker_entries_barrier__io_x_pal  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_paa  =  dcache__pma_checker_entries_barrier__io_x_paa  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_eff  =  dcache__pma_checker_entries_barrier__io_x_eff  ; 
  assign   dcache__pma_checker_entries_barrier__io_y_c  =  dcache__pma_checker_entries_barrier__io_x_c  ;
  
  
 
  assign   dcache__pma_checker_entries_barrier_1__io_y_u  =  dcache__pma_checker_entries_barrier_1__io_x_u  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_ae_ptw  =  dcache__pma_checker_entries_barrier_1__io_x_ae_ptw  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_ae_final  =  dcache__pma_checker_entries_barrier_1__io_x_ae_final  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_pf  =  dcache__pma_checker_entries_barrier_1__io_x_pf  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_gf  =  dcache__pma_checker_entries_barrier_1__io_x_gf  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_sw  =  dcache__pma_checker_entries_barrier_1__io_x_sw  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_sx  =  dcache__pma_checker_entries_barrier_1__io_x_sx  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_sr  =  dcache__pma_checker_entries_barrier_1__io_x_sr  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_pw  =  dcache__pma_checker_entries_barrier_1__io_x_pw  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_px  =  dcache__pma_checker_entries_barrier_1__io_x_px  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_pr  =  dcache__pma_checker_entries_barrier_1__io_x_pr  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_ppp  =  dcache__pma_checker_entries_barrier_1__io_x_ppp  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_pal  =  dcache__pma_checker_entries_barrier_1__io_x_pal  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_paa  =  dcache__pma_checker_entries_barrier_1__io_x_paa  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_eff  =  dcache__pma_checker_entries_barrier_1__io_x_eff  ; 
  assign   dcache__pma_checker_entries_barrier_1__io_y_c  =  dcache__pma_checker_entries_barrier_1__io_x_c  ;
  
  
 
  assign   dcache__pma_checker_entries_barrier_2__io_y_u  =  dcache__pma_checker_entries_barrier_2__io_x_u  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_ae_ptw  =  dcache__pma_checker_entries_barrier_2__io_x_ae_ptw  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_ae_final  =  dcache__pma_checker_entries_barrier_2__io_x_ae_final  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_pf  =  dcache__pma_checker_entries_barrier_2__io_x_pf  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_gf  =  dcache__pma_checker_entries_barrier_2__io_x_gf  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_sw  =  dcache__pma_checker_entries_barrier_2__io_x_sw  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_sx  =  dcache__pma_checker_entries_barrier_2__io_x_sx  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_sr  =  dcache__pma_checker_entries_barrier_2__io_x_sr  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_pw  =  dcache__pma_checker_entries_barrier_2__io_x_pw  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_px  =  dcache__pma_checker_entries_barrier_2__io_x_px  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_pr  =  dcache__pma_checker_entries_barrier_2__io_x_pr  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_ppp  =  dcache__pma_checker_entries_barrier_2__io_x_ppp  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_pal  =  dcache__pma_checker_entries_barrier_2__io_x_pal  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_paa  =  dcache__pma_checker_entries_barrier_2__io_x_paa  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_eff  =  dcache__pma_checker_entries_barrier_2__io_x_eff  ; 
  assign   dcache__pma_checker_entries_barrier_2__io_y_c  =  dcache__pma_checker_entries_barrier_2__io_x_c  ;
  
  
 
  assign   dcache__pma_checker_entries_barrier_3__io_y_u  =  dcache__pma_checker_entries_barrier_3__io_x_u  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_ae_ptw  =  dcache__pma_checker_entries_barrier_3__io_x_ae_ptw  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_ae_final  =  dcache__pma_checker_entries_barrier_3__io_x_ae_final  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_pf  =  dcache__pma_checker_entries_barrier_3__io_x_pf  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_gf  =  dcache__pma_checker_entries_barrier_3__io_x_gf  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_sw  =  dcache__pma_checker_entries_barrier_3__io_x_sw  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_sx  =  dcache__pma_checker_entries_barrier_3__io_x_sx  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_sr  =  dcache__pma_checker_entries_barrier_3__io_x_sr  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_pw  =  dcache__pma_checker_entries_barrier_3__io_x_pw  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_px  =  dcache__pma_checker_entries_barrier_3__io_x_px  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_pr  =  dcache__pma_checker_entries_barrier_3__io_x_pr  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_ppp  =  dcache__pma_checker_entries_barrier_3__io_x_ppp  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_pal  =  dcache__pma_checker_entries_barrier_3__io_x_pal  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_paa  =  dcache__pma_checker_entries_barrier_3__io_x_paa  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_eff  =  dcache__pma_checker_entries_barrier_3__io_x_eff  ; 
  assign   dcache__pma_checker_entries_barrier_3__io_y_c  =  dcache__pma_checker_entries_barrier_3__io_x_c  ;
  
  
 
  assign   dcache__pma_checker_entries_barrier_4__io_y_u  =  dcache__pma_checker_entries_barrier_4__io_x_u  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_ae_ptw  =  dcache__pma_checker_entries_barrier_4__io_x_ae_ptw  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_ae_final  =  dcache__pma_checker_entries_barrier_4__io_x_ae_final  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_pf  =  dcache__pma_checker_entries_barrier_4__io_x_pf  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_gf  =  dcache__pma_checker_entries_barrier_4__io_x_gf  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_sw  =  dcache__pma_checker_entries_barrier_4__io_x_sw  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_sx  =  dcache__pma_checker_entries_barrier_4__io_x_sx  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_sr  =  dcache__pma_checker_entries_barrier_4__io_x_sr  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_pw  =  dcache__pma_checker_entries_barrier_4__io_x_pw  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_px  =  dcache__pma_checker_entries_barrier_4__io_x_px  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_pr  =  dcache__pma_checker_entries_barrier_4__io_x_pr  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_ppp  =  dcache__pma_checker_entries_barrier_4__io_x_ppp  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_pal  =  dcache__pma_checker_entries_barrier_4__io_x_pal  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_paa  =  dcache__pma_checker_entries_barrier_4__io_x_paa  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_eff  =  dcache__pma_checker_entries_barrier_4__io_x_eff  ; 
  assign   dcache__pma_checker_entries_barrier_4__io_y_c  =  dcache__pma_checker_entries_barrier_4__io_x_c  ;
assign dcache__tlb_entries_barrier__io_x_u = 1'h0;
assign dcache__tlb_entries_barrier__io_x_ae_ptw = 1'h0;
assign dcache__tlb_entries_barrier__io_x_ae_final = 1'h0;
assign dcache__tlb_entries_barrier__io_x_pf = 1'h0;
assign dcache__tlb_entries_barrier__io_x_gf = 1'h0;
assign dcache__tlb_entries_barrier__io_x_sw = 1'h0;
assign dcache__tlb_entries_barrier__io_x_sx = 1'h0;
assign dcache__tlb_entries_barrier__io_x_sr = 1'h0;
assign dcache__tlb_entries_barrier__io_x_pw = 1'h0;
assign dcache__tlb_entries_barrier__io_x_px = 1'h0;
assign dcache__tlb_entries_barrier__io_x_pr = 1'h0;
assign dcache__tlb_entries_barrier__io_x_ppp = 1'h0;
assign dcache__tlb_entries_barrier__io_x_pal = 1'h0;
assign dcache__tlb_entries_barrier__io_x_paa = 1'h0;
assign dcache__tlb_entries_barrier__io_x_eff = 1'h0;
assign dcache__tlb_entries_barrier__io_x_c = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_u = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_ae_ptw = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_ae_final = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_pf = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_gf = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_sw = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_sx = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_sr = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_pw = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_px = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_pr = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_ppp = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_pal = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_paa = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_eff = 1'h0;
assign dcache__tlb_entries_barrier_1__io_x_c = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_u = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_ae_ptw = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_ae_final = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_pf = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_gf = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_sw = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_sx = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_sr = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_pw = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_px = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_pr = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_ppp = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_pal = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_paa = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_eff = 1'h0;
assign dcache__tlb_entries_barrier_2__io_x_c = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_u = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_ae_ptw = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_ae_final = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_pf = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_gf = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_sw = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_sx = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_sr = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_pw = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_px = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_pr = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_ppp = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_pal = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_paa = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_eff = 1'h0;
assign dcache__tlb_entries_barrier_3__io_x_c = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_u = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_ae_ptw = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_ae_final = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_pf = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_gf = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_sw = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_sx = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_sr = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_pw = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_px = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_pr = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_ppp = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_pal = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_paa = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_eff = 1'h0;
assign dcache__tlb_entries_barrier_4__io_x_c = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_u = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_ae_ptw = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_ae_final = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_pf = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_gf = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_sw = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_sx = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_sr = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_pw = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_px = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_pr = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_ppp = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_pal = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_paa = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_eff = 1'h0;
assign dcache__tlb_entries_barrier_5__io_x_c = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_u = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_ae_ptw = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_ae_final = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_pf = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_gf = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_sw = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_sx = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_sr = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_pw = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_px = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_pr = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_ppp = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_pal = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_paa = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_eff = 1'h0;
assign dcache__pma_checker_entries_barrier__io_x_c = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_u = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_ae_ptw = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_ae_final = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_pf = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_gf = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_sw = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_sx = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_sr = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_pw = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_px = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_pr = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_ppp = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_pal = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_paa = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_eff = 1'h0;
assign dcache__pma_checker_entries_barrier_1__io_x_c = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_u = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_ae_ptw = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_ae_final = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_pf = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_gf = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_sw = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_sx = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_sr = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_pw = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_px = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_pr = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_ppp = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_pal = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_paa = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_eff = 1'h0;
assign dcache__pma_checker_entries_barrier_2__io_x_c = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_u = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_ae_ptw = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_ae_final = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_pf = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_gf = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_sw = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_sx = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_sr = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_pw = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_px = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_pr = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_ppp = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_pal = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_paa = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_eff = 1'h0;
assign dcache__pma_checker_entries_barrier_3__io_x_c = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_u = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_ae_ptw = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_ae_final = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_pf = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_gf = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_sw = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_sx = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_sr = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_pw = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_px = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_pr = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_ppp = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_pal = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_paa = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_eff = 1'h0;
assign dcache__pma_checker_entries_barrier_4__io_x_c = 1'h0;
  
  
wire [5:0] dcache__tag_array_0_ext__RW0_addr;
wire  dcache__tag_array_0_ext__RW0_en;
wire  dcache__tag_array_0_ext__RW0_clk;
wire  dcache__tag_array_0_ext__RW0_wmode;
wire [21:0] dcache__tag_array_0_ext__RW0_wdata;
wire [21:0] dcache__tag_array_0_ext__RW0_rdata;
 
   reg[21:0]  dcache__tag_array_0_ext__Memory  [0:63]; 
   reg[5:0]  dcache__tag_array_0_ext___RW0_raddr_d0  ; 
   reg  dcache__tag_array_0_ext___RW0_ren_d0  ; 
   reg  dcache__tag_array_0_ext___RW0_rmode_d0  ; 
  always @( posedge   dcache__tag_array_0_ext__RW0_clk  )
       begin  
          dcache__tag_array_0_ext___RW0_raddr_d0   <=  dcache__tag_array_0_ext__RW0_addr  ; 
          dcache__tag_array_0_ext___RW0_ren_d0   <=  dcache__tag_array_0_ext__RW0_en  ; 
          dcache__tag_array_0_ext___RW0_rmode_d0   <=  dcache__tag_array_0_ext__RW0_wmode  ;
         if (  dcache__tag_array_0_ext__RW0_en  &  dcache__tag_array_0_ext__RW0_wmode  &1'h1) 
             dcache__tag_array_0_ext__Memory   [  dcache__tag_array_0_ext__RW0_addr  ]<=  dcache__tag_array_0_ext__RW0_wdata  ;
       end
  
  assign   dcache__tag_array_0_ext__RW0_rdata  =  dcache__tag_array_0_ext___RW0_ren_d0  &~  dcache__tag_array_0_ext___RW0_rmode_d0   ?   dcache__tag_array_0_ext__Memory  [  dcache__tag_array_0_ext___RW0_raddr_d0  ]:22'bx;
assign dcache__tag_array_0_ext__RW0_addr = dcache__resetting ? dcache__flushCounter:dcache___GEN ? dcache__metaArb_io_in_bits_idx_3:dcache__metaArb_io_in_valid_4 ? dcache__metaArb_io_in_bits_idx_4:dcache__metaArb_io_in_valid_6 ? dcache__metaArb_io_in_bits_idx_6:dcache__metaArb_io_in_bits_idx_7;
assign dcache__tag_array_0_ext__RW0_en = dcache__readEnable|dcache__writeEnable;
assign dcache__tag_array_0_ext__RW0_clk = dcache__clock;
assign dcache__tag_array_0_ext__RW0_wmode = dcache__metaArb_io_out_bits_write;
assign dcache__tag_array_0_ext__RW0_wdata = dcache__resetting ? 22'h0:dcache__metaArb_io_in_valid_2 ? dcache__metaArb_io_in_bits_data_2:dcache__metaArb_io_in_valid_3 ? dcache__metaArb_io_in_bits_data_3:dcache__metaArb_io_in_bits_data_7;
assign dcache___tag_array_0_ext_RW0_rdata = dcache__tag_array_0_ext__RW0_rdata;
  
  
wire  dcache__data__clock;
wire  dcache__data__io_req_valid;
wire [11:0] dcache__data__io_req_bits_addr;
wire  dcache__data__io_req_bits_write;
wire [63:0] dcache__data__io_req_bits_wdata;
wire [7:0] dcache__data__io_req_bits_eccMask;
wire [63:0] dcache__data__io_resp_0;
 
   wire  dcache__data__data_arrays_0_rdata_data_en  ; 
   wire  dcache__data__data_arrays_0_rdata_MPORT_en  ; 
  assign   dcache__data__data_arrays_0_rdata_MPORT_en  =  dcache__data__io_req_valid  &  dcache__data__io_req_bits_write  ; 
  assign   dcache__data__data_arrays_0_rdata_data_en  =  dcache__data__io_req_valid  &~  dcache__data__io_req_bits_write  ;  
  
wire [8:0] dcache__data__data_arrays_0_ext__RW0_addr;
wire  dcache__data__data_arrays_0_ext__RW0_en;
wire  dcache__data__data_arrays_0_ext__RW0_clk;
wire  dcache__data__data_arrays_0_ext__RW0_wmode;
wire [63:0] dcache__data__data_arrays_0_ext__RW0_wdata;
wire [63:0] dcache__data__data_arrays_0_ext__RW0_rdata;
wire [7:0] dcache__data__data_arrays_0_ext__RW0_wmask;
 
   reg[63:0]  dcache__data__data_arrays_0_ext__Memory  [0:511]; 
   reg[8:0]  dcache__data__data_arrays_0_ext___RW0_raddr_d0  ; 
   reg  dcache__data__data_arrays_0_ext___RW0_ren_d0  ; 
   reg  dcache__data__data_arrays_0_ext___RW0_rmode_d0  ; 
  always @( posedge   dcache__data__data_arrays_0_ext__RW0_clk  )
       begin  
          dcache__data__data_arrays_0_ext___RW0_raddr_d0   <=  dcache__data__data_arrays_0_ext__RW0_addr  ; 
          dcache__data__data_arrays_0_ext___RW0_ren_d0   <=  dcache__data__data_arrays_0_ext__RW0_en  ; 
          dcache__data__data_arrays_0_ext___RW0_rmode_d0   <=  dcache__data__data_arrays_0_ext__RW0_wmode  ;
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [0]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h0+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [7:0];
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [1]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h8+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [15:8];
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [2]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h10+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [23:16];
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [3]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h18+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [31:24];
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [4]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h20+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [39:32];
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [5]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h28+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [47:40];
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [6]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h30+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [55:48];
         if (  dcache__data__data_arrays_0_ext__RW0_en  &  dcache__data__data_arrays_0_ext__RW0_wmask  [7]&  dcache__data__data_arrays_0_ext__RW0_wmode  ) 
             dcache__data__data_arrays_0_ext__Memory   [  dcache__data__data_arrays_0_ext__RW0_addr  ][32'h38+:8]<=  dcache__data__data_arrays_0_ext__RW0_wdata  [63:56];
       end
  
  assign   dcache__data__data_arrays_0_ext__RW0_rdata  =  dcache__data__data_arrays_0_ext___RW0_ren_d0  &~  dcache__data__data_arrays_0_ext___RW0_rmode_d0   ?   dcache__data__data_arrays_0_ext__Memory  [  dcache__data__data_arrays_0_ext___RW0_raddr_d0  ]:64'bx;
assign dcache__data__data_arrays_0_ext__RW0_addr = dcache__data__io_req_bits_addr[11:3];
assign dcache__data__data_arrays_0_ext__RW0_en = dcache__data__data_arrays_0_rdata_data_en|dcache__data__data_arrays_0_rdata_MPORT_en;
assign dcache__data__data_arrays_0_ext__RW0_clk = dcache__data__clock;
assign dcache__data__data_arrays_0_ext__RW0_wmode = dcache__data__io_req_bits_write;
assign dcache__data__data_arrays_0_ext__RW0_wdata = dcache__data__io_req_bits_wdata;
assign dcache__data__io_resp_0 = dcache__data__data_arrays_0_ext__RW0_rdata;
assign dcache__data__data_arrays_0_ext__RW0_wmask = dcache__data__io_req_bits_eccMask;

assign dcache__data__clock = dcache__clock;
assign dcache__data__io_req_valid = dcache__dataArb_io_out_valid;
assign dcache__data__io_req_bits_addr = dcache__dataArb_io_in_valid_0 ? dcache___dataArb_io_in_0_bits_wordMask_wordMask_T:dcache__dataArb_io_in_valid_1 ? dcache__dataArb_io_in_bits_addr_1:dcache__dataArb_io_in_valid_2 ? dcache__dataArb_io_in_bits_addr_2:dcache__dataArb_io_in_bits_addr_3;
assign dcache__data__io_req_bits_write = dcache__dataArb_io_in_valid_0 ? dcache__pstore_drain:dcache__dataArb_io_in_valid_1&dcache__dataArb_io_in_bits_write_1;
assign dcache__data__io_req_bits_wdata = dcache__dataArb_io_in_valid_0 ? dcache__dataArb_io_in_bits_wdata_0:dcache__auto_out_d_bits_data;
assign dcache__data__io_req_bits_eccMask = dcache__dataArb_io_in_valid_0 ? dcache__dataArb_io_in_bits_eccMask_0:8'hFF;
assign dcache___data_io_resp_0 = dcache__data__io_resp_0;
  
  
wire [7:0] dcache__amoalus_0__io_mask;
wire [4:0] dcache__amoalus_0__io_cmd;
wire [63:0] dcache__amoalus_0__io_lhs;
wire [63:0] dcache__amoalus_0__io_rhs;
wire [63:0] dcache__amoalus_0__io_out;
 
   wire  dcache__amoalus_0___logic_xor_T_1  =  dcache__amoalus_0__io_cmd  ==5'hA; 
   wire  dcache__amoalus_0__logic_and  =  dcache__amoalus_0___logic_xor_T_1  |  dcache__amoalus_0__io_cmd  ==5'hB; 
   wire  dcache__amoalus_0__logic_xor  =  dcache__amoalus_0__io_cmd  ==5'h9|  dcache__amoalus_0___logic_xor_T_1  ; 
   wire[63:0]  dcache__amoalus_0__adder_out_mask  ={32'hFFFFFFFF,  dcache__amoalus_0__io_mask  [3],31'h7FFFFFFF}; 
   wire[63:0]  dcache__amoalus_0__wmask  ={{8{  dcache__amoalus_0__io_mask  [7]}},{8{  dcache__amoalus_0__io_mask  [6]}},{8{  dcache__amoalus_0__io_mask  [5]}},{8{  dcache__amoalus_0__io_mask  [4]}},{8{  dcache__amoalus_0__io_mask  [3]}},{8{  dcache__amoalus_0__io_mask  [2]}},{8{  dcache__amoalus_0__io_mask  [1]}},{8{  dcache__amoalus_0__io_mask  [0]}}}; 
  assign   dcache__amoalus_0__io_out  =  dcache__amoalus_0__wmask  &(  dcache__amoalus_0__io_cmd  ==5'h8 ? (  dcache__amoalus_0__io_lhs  &  dcache__amoalus_0__adder_out_mask  )+(  dcache__amoalus_0__io_rhs  &  dcache__amoalus_0__adder_out_mask  ):  dcache__amoalus_0__logic_and  |  dcache__amoalus_0__logic_xor   ? (  dcache__amoalus_0__logic_and   ?   dcache__amoalus_0__io_lhs  &  dcache__amoalus_0__io_rhs  :64'h0)|(  dcache__amoalus_0__logic_xor   ?   dcache__amoalus_0__io_lhs  ^  dcache__amoalus_0__io_rhs  :64'h0):((  dcache__amoalus_0__io_mask  [4] ? (  dcache__amoalus_0__io_lhs  [63]==  dcache__amoalus_0__io_rhs  [63] ?   dcache__amoalus_0__io_lhs  [63:32]<  dcache__amoalus_0__io_rhs  [63:32]|  dcache__amoalus_0__io_lhs  [63:32]==  dcache__amoalus_0__io_rhs  [63:32]&  dcache__amoalus_0__io_lhs  [31:0]<  dcache__amoalus_0__io_rhs  [31:0]:  dcache__amoalus_0__io_cmd  [1] ?   dcache__amoalus_0__io_rhs  [63]:  dcache__amoalus_0__io_lhs  [63]):  dcache__amoalus_0__io_lhs  [31]==  dcache__amoalus_0__io_rhs  [31] ?   dcache__amoalus_0__io_lhs  [31:0]<  dcache__amoalus_0__io_rhs  [31:0]:  dcache__amoalus_0__io_cmd  [1] ?   dcache__amoalus_0__io_rhs  [31]:  dcache__amoalus_0__io_lhs  [31]) ?   dcache__amoalus_0__io_cmd  ==5'hC|  dcache__amoalus_0__io_cmd  ==5'hE:  dcache__amoalus_0__io_cmd  ==5'hD|  dcache__amoalus_0__io_cmd  ==5'hF) ?   dcache__amoalus_0__io_lhs  :  dcache__amoalus_0__io_rhs  )|~  dcache__amoalus_0__wmask  &  dcache__amoalus_0__io_lhs  ;
assign dcache__amoalus_0__io_mask = dcache__pstore1_mask;
assign dcache__amoalus_0__io_cmd = dcache__pstore1_cmd;
assign dcache__amoalus_0__io_lhs = dcache__s2_data;
assign dcache__amoalus_0__io_rhs = dcache__pstore1_data;
assign dcache___amoalus_0_io_out = dcache__amoalus_0__io_out;
 
  assign   dcache__auto_out_a_valid  =  dcache__tl_out_a_valid  ; 
  assign   dcache__auto_out_a_bits_opcode  =  dcache__s2_pma_cacheable   ? 3'h6:  dcache__s2_write   ? (  dcache___metaArb_io_in_3_bits_data_c_cat_T_24   ? 3'h1:  dcache__s2_read   ? (  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35   ? 3'h2:  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28   ? 3'h3:3'h0):3'h0):3'h4; 
  assign   dcache__auto_out_a_bits_param  =  dcache__s2_pma_cacheable   ? {1'h0,  dcache__casez_tmp  }:~  dcache__s2_write  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |~  dcache__s2_read   ? 3'h0:  dcache___metaArb_io_in_3_bits_data_c_cat_T_39   ? 3'h3:  dcache___metaArb_io_in_3_bits_data_c_cat_T_38   ? 3'h2:  dcache___metaArb_io_in_3_bits_data_c_cat_T_37   ? 3'h1:  dcache___metaArb_io_in_3_bits_data_c_cat_T_36   ? 3'h0:  dcache___metaArb_io_in_3_bits_data_c_cat_T_35   ? 3'h4:  dcache___metaArb_io_in_3_bits_data_c_cat_T_31   ? 3'h2:  dcache___metaArb_io_in_3_bits_data_c_cat_T_30   ? 3'h1:  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |~  dcache___metaArb_io_in_3_bits_data_c_cat_T_28   ? 3'h0:3'h3; 
  assign   dcache__auto_out_a_bits_size  =  dcache__s2_pma_cacheable   ? 4'h6:  dcache___GEN_16   ? {2'h0,  dcache__s2_req_size  }:4'h0; 
  assign   dcache__auto_out_a_bits_source  =~  dcache__s2_pma_cacheable  &(~  dcache__s2_write  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |~  dcache__s2_read  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  ); 
  assign   dcache__auto_out_a_bits_address  =  dcache__s2_pma_cacheable   ? {  dcache__s2_req_addr  [31:6],6'h0}:  dcache___GEN_16   ?   dcache__s2_req_addr  [31:0]:32'h0; 
  assign   dcache__auto_out_a_bits_mask  =  dcache__s2_pma_cacheable   ? 8'hFF:  dcache__s2_write   ? (  dcache___metaArb_io_in_3_bits_data_c_cat_T_24   ?   dcache__pstore1_mask  :  dcache__s2_read   ?   dcache__atomics_mask  :{  dcache__put_a_mask_acc_5  |  dcache__put_a_mask_eq_5  &  dcache__s2_req_addr  [0],  dcache__put_a_mask_acc_5  |  dcache__put_a_mask_eq_5  &~(  dcache__s2_req_addr  [0]),  dcache__put_a_mask_acc_4  |  dcache__put_a_mask_eq_4  &  dcache__s2_req_addr  [0],  dcache__put_a_mask_acc_4  |  dcache__put_a_mask_eq_4  &~(  dcache__s2_req_addr  [0]),  dcache__put_a_mask_acc_3  |  dcache__put_a_mask_eq_3  &  dcache__s2_req_addr  [0],  dcache__put_a_mask_acc_3  |  dcache__put_a_mask_eq_3  &~(  dcache__s2_req_addr  [0]),  dcache__put_a_mask_acc_2  |  dcache__put_a_mask_eq_2  &  dcache__s2_req_addr  [0],  dcache__put_a_mask_acc_2  |  dcache__put_a_mask_eq_2  &~(  dcache__s2_req_addr  [0])}):{  dcache__get_a_mask_acc_5  |  dcache__get_a_mask_eq_5  &  dcache__s2_req_addr  [0],  dcache__get_a_mask_acc_5  |  dcache__get_a_mask_eq_5  &~(  dcache__s2_req_addr  [0]),  dcache__get_a_mask_acc_4  |  dcache__get_a_mask_eq_4  &  dcache__s2_req_addr  [0],  dcache__get_a_mask_acc_4  |  dcache__get_a_mask_eq_4  &~(  dcache__s2_req_addr  [0]),  dcache__get_a_mask_acc_3  |  dcache__get_a_mask_eq_3  &  dcache__s2_req_addr  [0],  dcache__get_a_mask_acc_3  |  dcache__get_a_mask_eq_3  &~(  dcache__s2_req_addr  [0]),  dcache__get_a_mask_acc_2  |  dcache__get_a_mask_eq_2  &  dcache__s2_req_addr  [0],  dcache__get_a_mask_acc_2  |  dcache__get_a_mask_eq_2  &~(  dcache__s2_req_addr  [0])}; 
  assign   dcache__auto_out_a_bits_data  =  dcache__s2_pma_cacheable  |~  dcache__s2_write  |~(  dcache___metaArb_io_in_3_bits_data_c_cat_T_24  |~  dcache__s2_read  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_39  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_38  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_37  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_36  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_35  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_31  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_30  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_29  |  dcache___metaArb_io_in_3_bits_data_c_cat_T_28  ) ? 64'h0:  dcache__pstore1_data  ; 
  assign   dcache__auto_out_b_ready  =  dcache__nodeOut_b_ready  ; 
  assign   dcache__auto_out_c_valid  =  dcache__nodeOut_c_valid  ; 
  assign   dcache__auto_out_c_bits_opcode  =  dcache__nodeOut_c_bits_opcode  ; 
  assign   dcache__auto_out_c_bits_param  =  dcache___GEN_27   ? ((&  dcache__s2_victim_state_state  )|  dcache__s2_victim_state_state  ==2'h2 ? 3'h1:  dcache__s2_victim_state_state  ==2'h1 ? 3'h2:  dcache__s2_victim_state_state  ==2'h0 ? 3'h5:3'h0):  dcache___inWriteback_T_1  |  dcache___GEN_26  |~(~  dcache__s2_probe  |  dcache__s2_prb_ack_data  |~(|  dcache__s2_probe_state_state  )) ? (  dcache___GEN_13   ? 3'h3:  dcache___GEN_10   ? 3'h4:  dcache___GEN_9   ? 3'h5:  dcache___GEN_8  |  dcache___GEN_7   ? 3'h0:  dcache___GEN_6   ? 3'h4:  dcache___GEN_5   ? 3'h5:  dcache___GEN_4  |  dcache___GEN_3  ==4'hA ? 3'h1:  dcache___GEN_3  ==4'h9 ? 3'h2:  dcache___GEN_3  ==4'h8 ? 3'h5:3'h0):3'h5; 
  assign   dcache__auto_out_c_bits_size  =  dcache__nodeOut_c_bits_size  ; 
  assign   dcache__auto_out_c_bits_source  =  dcache__probe_bits_source  ; 
  assign   dcache__auto_out_c_bits_address  =  dcache__probe_bits_address  ; 
  assign   dcache__auto_out_c_bits_data  =  dcache__s2_data  ; 
  assign   dcache__auto_out_d_ready  =  dcache__nodeOut_d_ready  ; 
  assign   dcache__auto_out_e_valid  =  dcache__nodeOut_e_valid  ; 
  assign   dcache__auto_out_e_bits_sink  =  dcache__auto_out_d_bits_sink  ; 
  assign   dcache__io_cpu_req_ready  =  dcache__io_cpu_req_ready_0  ; 
  assign   dcache__io_cpu_s2_nack  =  dcache__io_cpu_s2_nack_0  ; 
  assign   dcache__io_cpu_resp_valid  =  dcache__s2_valid_hit_pre_data_ecc_and_waw  |  dcache__doUncachedResp  ; 
  assign   dcache__io_cpu_resp_bits_addr  =  dcache__doUncachedResp   ?   dcache__s2_uncached_resp_addr  :  dcache__s2_req_addr  ; 
  assign   dcache__io_cpu_resp_bits_tag  =  dcache__s2_req_tag  ; 
  assign   dcache__io_cpu_resp_bits_cmd  =  dcache__s2_req_cmd  ; 
  assign   dcache__io_cpu_resp_bits_size  =  dcache__s2_req_size  ; 
  assign   dcache__io_cpu_resp_bits_signed  =  dcache__s2_req_signed  ; 
  assign   dcache__io_cpu_resp_bits_dprv  =  dcache__s2_req_dprv  ; 
  assign   dcache__io_cpu_resp_bits_dv  =  dcache__s2_req_dv  ; 
  assign   dcache__io_cpu_resp_bits_data  ={  dcache__s2_req_size  ==2'h0|  dcache__s2_sc   ? {56{  dcache__s2_req_signed  &  dcache__io_cpu_resp_bits_data_zeroed_2  [7]}}:{  dcache__s2_req_size  ==2'h1 ? {48{  dcache__s2_req_signed  &  dcache__io_cpu_resp_bits_data_zeroed_1  [15]}}:{  dcache___io_cpu_resp_bits_data_word_bypass_T_1   ? {32{  dcache__s2_req_signed  &  dcache__io_cpu_resp_bits_data_zeroed  [31]}}:  dcache__s2_data  [63:32],  dcache__io_cpu_resp_bits_data_zeroed  [31:16]},  dcache__io_cpu_resp_bits_data_zeroed_1  [15:8]},  dcache__io_cpu_resp_bits_data_zeroed_2  [7:1],  dcache__io_cpu_resp_bits_data_zeroed_2  [0]|  dcache__s2_sc_fail  }; 
  assign   dcache__io_cpu_resp_bits_mask  =8'h0; 
  assign   dcache__io_cpu_resp_bits_replay  =  dcache__doUncachedResp  ; 
  assign   dcache__io_cpu_resp_bits_has_data  =  dcache__s2_read  ; 
  assign   dcache__io_cpu_resp_bits_data_word_bypass  ={  dcache___io_cpu_resp_bits_data_word_bypass_T_1   ? {32{  dcache__s2_req_signed  &  dcache__io_cpu_resp_bits_data_word_bypass_zeroed  [31]}}:  dcache__s2_data  [63:32],  dcache__io_cpu_resp_bits_data_word_bypass_zeroed  }; 
  assign   dcache__io_cpu_resp_bits_data_raw  =  dcache__s2_data  ; 
  assign   dcache__io_cpu_resp_bits_store_data  =  dcache__pstore1_data  ; 
  assign   dcache__io_cpu_replay_next  =  dcache__io_cpu_replay_next_0  ; 
  assign   dcache__io_cpu_s2_xcpt_ma_ld  =  dcache__io_cpu_s2_xcpt_ma_ld_0  ; 
  assign   dcache__io_cpu_s2_xcpt_ma_st  =  dcache__io_cpu_s2_xcpt_ma_st_0  ; 
  assign   dcache__io_cpu_s2_xcpt_pf_ld  =  dcache__io_cpu_s2_xcpt_pf_ld_0  ; 
  assign   dcache__io_cpu_s2_xcpt_pf_st  =  dcache__io_cpu_s2_xcpt_pf_st_0  ; 
  assign   dcache__io_cpu_s2_xcpt_ae_ld  =  dcache__io_cpu_s2_xcpt_ae_ld_0  ; 
  assign   dcache__io_cpu_s2_xcpt_ae_st  =  dcache__io_cpu_s2_xcpt_ae_st_0  ; 
  assign   dcache__io_cpu_ordered  =~(  dcache__s1_valid  |  dcache__s2_valid  |  dcache__cached_grant_wait  |  dcache__uncachedInFlight_0  ); 
  assign   dcache__io_cpu_perf_release  =(  dcache__io_cpu_perf_release_counter  ==9'h1|  dcache__io_cpu_perf_release_beats1  ==9'h0)&  dcache___io_cpu_perf_release_T  ; 
  assign   dcache__io_cpu_perf_grant  =  dcache__auto_out_d_valid  &  dcache__d_last  ; 
  assign   dcache__io_ptw_req_bits_bits_need_gpa  =1'h0; 
  assign   dcache__io_ptw_req_bits_bits_stage2  =1'h0;
assign dcache__clock = clock;
assign dcache__reset = reset;
assign dcache__auto_out_a_ready = _tlMasterXbar_auto_in_0_a_ready;
assign _dcache_auto_out_a_valid = dcache__auto_out_a_valid;
assign _dcache_auto_out_a_bits_opcode = dcache__auto_out_a_bits_opcode;
assign _dcache_auto_out_a_bits_param = dcache__auto_out_a_bits_param;
assign _dcache_auto_out_a_bits_size = dcache__auto_out_a_bits_size;
assign _dcache_auto_out_a_bits_source = dcache__auto_out_a_bits_source;
assign _dcache_auto_out_a_bits_address = dcache__auto_out_a_bits_address;
assign _dcache_auto_out_a_bits_mask = dcache__auto_out_a_bits_mask;
assign _dcache_auto_out_a_bits_data = dcache__auto_out_a_bits_data;
assign _dcache_auto_out_b_ready = dcache__auto_out_b_ready;
assign dcache__auto_out_b_valid = _tlMasterXbar_auto_in_0_b_valid;
assign dcache__auto_out_b_bits_param = _tlMasterXbar_auto_in_0_b_bits_param;
assign dcache__auto_out_b_bits_size = _tlMasterXbar_auto_in_0_b_bits_size;
assign dcache__auto_out_b_bits_source = _tlMasterXbar_auto_in_0_b_bits_source;
assign dcache__auto_out_b_bits_address = _tlMasterXbar_auto_in_0_b_bits_address;
assign dcache__auto_out_c_ready = _tlMasterXbar_auto_in_0_c_ready;
assign _dcache_auto_out_c_valid = dcache__auto_out_c_valid;
assign _dcache_auto_out_c_bits_opcode = dcache__auto_out_c_bits_opcode;
assign _dcache_auto_out_c_bits_param = dcache__auto_out_c_bits_param;
assign _dcache_auto_out_c_bits_size = dcache__auto_out_c_bits_size;
assign _dcache_auto_out_c_bits_source = dcache__auto_out_c_bits_source;
assign _dcache_auto_out_c_bits_address = dcache__auto_out_c_bits_address;
assign _dcache_auto_out_c_bits_data = dcache__auto_out_c_bits_data;
assign _dcache_auto_out_d_ready = dcache__auto_out_d_ready;
assign dcache__auto_out_d_valid = _tlMasterXbar_auto_in_0_d_valid;
assign dcache__auto_out_d_bits_opcode = _tlMasterXbar_auto_in_0_d_bits_opcode;
assign dcache__auto_out_d_bits_param = _tlMasterXbar_auto_in_0_d_bits_param;
assign dcache__auto_out_d_bits_size = _tlMasterXbar_auto_in_0_d_bits_size;
assign dcache__auto_out_d_bits_source = _tlMasterXbar_auto_in_0_d_bits_source;
assign dcache__auto_out_d_bits_sink = _tlMasterXbar_auto_in_0_d_bits_sink;
assign dcache__auto_out_d_bits_denied = _tlMasterXbar_auto_in_0_d_bits_denied;
assign dcache__auto_out_d_bits_data = _tlMasterXbar_auto_in_0_d_bits_data;
assign dcache__auto_out_e_ready = _tlMasterXbar_auto_in_0_e_ready;
assign _dcache_auto_out_e_valid = dcache__auto_out_e_valid;
assign _dcache_auto_out_e_bits_sink = dcache__auto_out_e_bits_sink;
assign _dcache_io_cpu_req_ready = dcache__io_cpu_req_ready;
assign dcache__io_cpu_req_valid = _dcacheArb_io_mem_req_valid;
assign dcache__io_cpu_req_bits_addr = _dcacheArb_io_mem_req_bits_addr;
assign dcache__io_cpu_req_bits_tag = _dcacheArb_io_mem_req_bits_tag;
assign dcache__io_cpu_req_bits_cmd = _dcacheArb_io_mem_req_bits_cmd;
assign dcache__io_cpu_req_bits_size = _dcacheArb_io_mem_req_bits_size;
assign dcache__io_cpu_req_bits_signed = _dcacheArb_io_mem_req_bits_signed;
assign dcache__io_cpu_req_bits_dv = _dcacheArb_io_mem_req_bits_dv;
assign dcache__io_cpu_s1_kill = _dcacheArb_io_mem_s1_kill;
assign dcache__io_cpu_s1_data_data = _dcacheArb_io_mem_s1_data_data;
assign dcache__io_cpu_s1_data_mask = 8'h0;
assign _dcache_io_cpu_s2_nack = dcache__io_cpu_s2_nack;
assign _dcache_io_cpu_resp_valid = dcache__io_cpu_resp_valid;
assign _dcache_io_cpu_resp_bits_tag = dcache__io_cpu_resp_bits_tag;
assign _dcache_io_cpu_resp_bits_data = dcache__io_cpu_resp_bits_data;
assign _dcache_io_cpu_resp_bits_replay = dcache__io_cpu_resp_bits_replay;
assign _dcache_io_cpu_resp_bits_has_data = dcache__io_cpu_resp_bits_has_data;
assign _dcache_io_cpu_resp_bits_data_word_bypass = dcache__io_cpu_resp_bits_data_word_bypass;
assign _dcache_io_cpu_replay_next = dcache__io_cpu_replay_next;
assign _dcache_io_cpu_s2_xcpt_ma_ld = dcache__io_cpu_s2_xcpt_ma_ld;
assign _dcache_io_cpu_s2_xcpt_ma_st = dcache__io_cpu_s2_xcpt_ma_st;
assign _dcache_io_cpu_s2_xcpt_pf_ld = dcache__io_cpu_s2_xcpt_pf_ld;
assign _dcache_io_cpu_s2_xcpt_pf_st = dcache__io_cpu_s2_xcpt_pf_st;
assign _dcache_io_cpu_s2_xcpt_ae_ld = dcache__io_cpu_s2_xcpt_ae_ld;
assign _dcache_io_cpu_s2_xcpt_ae_st = dcache__io_cpu_s2_xcpt_ae_st;
assign _dcache_io_cpu_ordered = dcache__io_cpu_ordered;
assign _dcache_io_cpu_perf_release = dcache__io_cpu_perf_release;
assign _dcache_io_cpu_perf_grant = dcache__io_cpu_perf_grant;
assign _dcache_io_ptw_req_bits_bits_need_gpa = dcache__io_ptw_req_bits_bits_need_gpa;
assign _dcache_io_ptw_req_bits_bits_stage2 = dcache__io_ptw_req_bits_bits_stage2;
assign dcache__io_ptw_status_debug = _ptw_io_requestor_0_status_debug;
assign dcache__io_ptw_pmp_cfg_l_0 = _ptw_io_requestor_0_pmp_cfg_l_0;
assign dcache__io_ptw_pmp_cfg_l_1 = _ptw_io_requestor_0_pmp_cfg_l_1;
assign dcache__io_ptw_pmp_cfg_l_2 = _ptw_io_requestor_0_pmp_cfg_l_2;
assign dcache__io_ptw_pmp_cfg_l_3 = _ptw_io_requestor_0_pmp_cfg_l_3;
assign dcache__io_ptw_pmp_cfg_l_4 = _ptw_io_requestor_0_pmp_cfg_l_4;
assign dcache__io_ptw_pmp_cfg_l_5 = _ptw_io_requestor_0_pmp_cfg_l_5;
assign dcache__io_ptw_pmp_cfg_l_6 = _ptw_io_requestor_0_pmp_cfg_l_6;
assign dcache__io_ptw_pmp_cfg_l_7 = _ptw_io_requestor_0_pmp_cfg_l_7;
assign dcache__io_ptw_pmp_cfg_a_0 = _ptw_io_requestor_0_pmp_cfg_a_0;
assign dcache__io_ptw_pmp_cfg_a_1 = _ptw_io_requestor_0_pmp_cfg_a_1;
assign dcache__io_ptw_pmp_cfg_a_2 = _ptw_io_requestor_0_pmp_cfg_a_2;
assign dcache__io_ptw_pmp_cfg_a_3 = _ptw_io_requestor_0_pmp_cfg_a_3;
assign dcache__io_ptw_pmp_cfg_a_4 = _ptw_io_requestor_0_pmp_cfg_a_4;
assign dcache__io_ptw_pmp_cfg_a_5 = _ptw_io_requestor_0_pmp_cfg_a_5;
assign dcache__io_ptw_pmp_cfg_a_6 = _ptw_io_requestor_0_pmp_cfg_a_6;
assign dcache__io_ptw_pmp_cfg_a_7 = _ptw_io_requestor_0_pmp_cfg_a_7;
assign dcache__io_ptw_pmp_cfg_w_0 = _ptw_io_requestor_0_pmp_cfg_w_0;
assign dcache__io_ptw_pmp_cfg_w_1 = _ptw_io_requestor_0_pmp_cfg_w_1;
assign dcache__io_ptw_pmp_cfg_w_2 = _ptw_io_requestor_0_pmp_cfg_w_2;
assign dcache__io_ptw_pmp_cfg_w_3 = _ptw_io_requestor_0_pmp_cfg_w_3;
assign dcache__io_ptw_pmp_cfg_w_4 = _ptw_io_requestor_0_pmp_cfg_w_4;
assign dcache__io_ptw_pmp_cfg_w_5 = _ptw_io_requestor_0_pmp_cfg_w_5;
assign dcache__io_ptw_pmp_cfg_w_6 = _ptw_io_requestor_0_pmp_cfg_w_6;
assign dcache__io_ptw_pmp_cfg_w_7 = _ptw_io_requestor_0_pmp_cfg_w_7;
assign dcache__io_ptw_pmp_cfg_r_0 = _ptw_io_requestor_0_pmp_cfg_r_0;
assign dcache__io_ptw_pmp_cfg_r_1 = _ptw_io_requestor_0_pmp_cfg_r_1;
assign dcache__io_ptw_pmp_cfg_r_2 = _ptw_io_requestor_0_pmp_cfg_r_2;
assign dcache__io_ptw_pmp_cfg_r_3 = _ptw_io_requestor_0_pmp_cfg_r_3;
assign dcache__io_ptw_pmp_cfg_r_4 = _ptw_io_requestor_0_pmp_cfg_r_4;
assign dcache__io_ptw_pmp_cfg_r_5 = _ptw_io_requestor_0_pmp_cfg_r_5;
assign dcache__io_ptw_pmp_cfg_r_6 = _ptw_io_requestor_0_pmp_cfg_r_6;
assign dcache__io_ptw_pmp_cfg_r_7 = _ptw_io_requestor_0_pmp_cfg_r_7;
assign dcache__io_ptw_pmp_addr_0 = _ptw_io_requestor_0_pmp_addr_0;
assign dcache__io_ptw_pmp_addr_1 = _ptw_io_requestor_0_pmp_addr_1;
assign dcache__io_ptw_pmp_addr_2 = _ptw_io_requestor_0_pmp_addr_2;
assign dcache__io_ptw_pmp_addr_3 = _ptw_io_requestor_0_pmp_addr_3;
assign dcache__io_ptw_pmp_addr_4 = _ptw_io_requestor_0_pmp_addr_4;
assign dcache__io_ptw_pmp_addr_5 = _ptw_io_requestor_0_pmp_addr_5;
assign dcache__io_ptw_pmp_addr_6 = _ptw_io_requestor_0_pmp_addr_6;
assign dcache__io_ptw_pmp_addr_7 = _ptw_io_requestor_0_pmp_addr_7;
assign dcache__io_ptw_pmp_mask_0 = _ptw_io_requestor_0_pmp_mask_0;
assign dcache__io_ptw_pmp_mask_1 = _ptw_io_requestor_0_pmp_mask_1;
assign dcache__io_ptw_pmp_mask_2 = _ptw_io_requestor_0_pmp_mask_2;
assign dcache__io_ptw_pmp_mask_3 = _ptw_io_requestor_0_pmp_mask_3;
assign dcache__io_ptw_pmp_mask_4 = _ptw_io_requestor_0_pmp_mask_4;
assign dcache__io_ptw_pmp_mask_5 = _ptw_io_requestor_0_pmp_mask_5;
assign dcache__io_ptw_pmp_mask_6 = _ptw_io_requestor_0_pmp_mask_6;
assign dcache__io_ptw_pmp_mask_7 = _ptw_io_requestor_0_pmp_mask_7;
 
  
wire  frontend__clock;
wire  frontend__reset;
wire  frontend__auto_icache_master_out_a_ready;
wire  frontend__auto_icache_master_out_a_valid;
wire [31:0] frontend__auto_icache_master_out_a_bits_address;
wire  frontend__auto_icache_master_out_d_valid;
wire [2:0] frontend__auto_icache_master_out_d_bits_opcode;
wire [3:0] frontend__auto_icache_master_out_d_bits_size;
wire [63:0] frontend__auto_icache_master_out_d_bits_data;
wire  frontend__auto_icache_master_out_d_bits_corrupt;
wire  frontend__io_cpu_might_request;
wire  frontend__io_cpu_req_valid;
wire [33:0] frontend__io_cpu_req_bits_pc;
wire  frontend__io_cpu_req_bits_speculative;
wire  frontend__io_cpu_resp_ready;
wire  frontend__io_cpu_resp_valid;
wire [33:0] frontend__io_cpu_resp_bits_pc;
wire [31:0] frontend__io_cpu_resp_bits_data;
wire  frontend__io_cpu_resp_bits_xcpt_pf_inst;
wire  frontend__io_cpu_resp_bits_xcpt_gf_inst;
wire  frontend__io_cpu_resp_bits_xcpt_ae_inst;
wire  frontend__io_cpu_resp_bits_replay;
wire  frontend__io_cpu_btb_update_valid;
wire  frontend__io_cpu_bht_update_valid;
wire  frontend__io_cpu_flush_icache;
wire  frontend__io_ptw_req_bits_bits_need_gpa;
wire  frontend__io_ptw_req_bits_bits_stage2;
wire  frontend__io_ptw_status_debug;
wire  frontend__io_ptw_pmp_cfg_l_0;
wire  frontend__io_ptw_pmp_cfg_l_1;
wire  frontend__io_ptw_pmp_cfg_l_2;
wire  frontend__io_ptw_pmp_cfg_l_3;
wire  frontend__io_ptw_pmp_cfg_l_4;
wire  frontend__io_ptw_pmp_cfg_l_5;
wire  frontend__io_ptw_pmp_cfg_l_6;
wire  frontend__io_ptw_pmp_cfg_l_7;
wire [1:0] frontend__io_ptw_pmp_cfg_a_0;
wire [1:0] frontend__io_ptw_pmp_cfg_a_1;
wire [1:0] frontend__io_ptw_pmp_cfg_a_2;
wire [1:0] frontend__io_ptw_pmp_cfg_a_3;
wire [1:0] frontend__io_ptw_pmp_cfg_a_4;
wire [1:0] frontend__io_ptw_pmp_cfg_a_5;
wire [1:0] frontend__io_ptw_pmp_cfg_a_6;
wire [1:0] frontend__io_ptw_pmp_cfg_a_7;
wire  frontend__io_ptw_pmp_cfg_x_0;
wire  frontend__io_ptw_pmp_cfg_x_1;
wire  frontend__io_ptw_pmp_cfg_x_2;
wire  frontend__io_ptw_pmp_cfg_x_3;
wire  frontend__io_ptw_pmp_cfg_x_4;
wire  frontend__io_ptw_pmp_cfg_x_5;
wire  frontend__io_ptw_pmp_cfg_x_6;
wire  frontend__io_ptw_pmp_cfg_x_7;
wire [29:0] frontend__io_ptw_pmp_addr_0;
wire [29:0] frontend__io_ptw_pmp_addr_1;
wire [29:0] frontend__io_ptw_pmp_addr_2;
wire [29:0] frontend__io_ptw_pmp_addr_3;
wire [29:0] frontend__io_ptw_pmp_addr_4;
wire [29:0] frontend__io_ptw_pmp_addr_5;
wire [29:0] frontend__io_ptw_pmp_addr_6;
wire [29:0] frontend__io_ptw_pmp_addr_7;
wire [31:0] frontend__io_ptw_pmp_mask_0;
wire [31:0] frontend__io_ptw_pmp_mask_1;
wire [31:0] frontend__io_ptw_pmp_mask_2;
wire [31:0] frontend__io_ptw_pmp_mask_3;
wire [31:0] frontend__io_ptw_pmp_mask_4;
wire [31:0] frontend__io_ptw_pmp_mask_5;
wire [31:0] frontend__io_ptw_pmp_mask_6;
wire [31:0] frontend__io_ptw_pmp_mask_7;
wire [63:0] frontend__io_ptw_customCSRs_csrs_0_value;
 
   wire[32:0]  frontend___io_cpu_npc_T  ; 
   wire  frontend__fq_io_enq_valid  ; 
   wire[31:0]  frontend___tlb_io_resp_paddr  ; 
   wire  frontend___tlb_io_resp_pf_inst  ; 
   wire  frontend___tlb_io_resp_ae_inst  ; 
   wire  frontend___tlb_io_resp_cacheable  ; 
   wire  frontend___fq_io_enq_ready  ; 
   wire[4:0]  frontend___fq_io_mask  ; 
   wire  frontend___icache_io_resp_valid  ; 
   wire[31:0]  frontend___icache_io_resp_bits_data  ; 
   wire  frontend___icache_io_resp_bits_ae  ; 
   reg  frontend__s1_valid  ; 
   reg  frontend__s2_valid  ; 
   wire  frontend__s0_valid  =  frontend__io_cpu_req_valid  |~(  frontend___fq_io_mask  [2])|~(  frontend___fq_io_mask  [3])&(~  frontend__s1_valid  |~  frontend__s2_valid  )|~(  frontend___fq_io_mask  [4])&~  frontend__s1_valid  &~  frontend__s2_valid  ; 
   reg[33:0]  frontend__s1_pc  ; 
   reg  frontend__s1_speculative  ; 
   reg[33:0]  frontend__s2_pc  ; 
   reg  frontend__s2_tlb_resp_pf_inst  ; 
   reg  frontend__s2_tlb_resp_ae_inst  ; 
   reg  frontend__s2_tlb_resp_cacheable  ; 
   wire  frontend___s2_xcpt_T  =  frontend__s2_tlb_resp_ae_inst  |  frontend__s2_tlb_resp_pf_inst  ; 
   reg  frontend__s2_speculative  ; 
   wire[33:0]  frontend__predicted_npc  ={  frontend__s1_pc  [33:2],2'h0}+34'h4; 
   reg  frontend__s2_replay_REG  ; 
   wire  frontend__s2_replay  =  frontend__s2_valid  &~(  frontend___fq_io_enq_ready  &  frontend__fq_io_enq_valid  )|  frontend__s2_replay_REG  ; 
   wire  frontend__icache_io_s2_kill  =  frontend__s2_speculative  &~(  frontend__s2_tlb_resp_cacheable  &~(  frontend__io_ptw_customCSRs_csrs_0_value  [3]))|  frontend___s2_xcpt_T  ; 
   reg  frontend__fq_io_enq_valid_REG  ; 
  assign   frontend__fq_io_enq_valid  =  frontend__fq_io_enq_valid_REG  &  frontend__s2_valid  &(  frontend___icache_io_resp_valid  |  frontend__icache_io_s2_kill  ); 
  assign   frontend___io_cpu_npc_T  =  frontend__io_cpu_req_valid   ?   frontend__io_cpu_req_bits_pc  [33:1]:  frontend__s2_replay   ?   frontend__s2_pc  [33:1]:  frontend__predicted_npc  [33:1]; 
  always @( posedge   frontend__clock  )
       begin 
         if (~  frontend__reset  &~(~(  frontend__io_cpu_req_valid  |  frontend__io_cpu_flush_icache  |  frontend__io_cpu_bht_update_valid  |  frontend__io_cpu_btb_update_valid  )|  frontend__io_cpu_might_request  ))
            begin 
              if (1)$display("Assertion failed\n    at Frontend.scala:92 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n");
              if (1)$display("");
            end 
         if (~  frontend__reset  &  frontend__s2_speculative  &  frontend__io_ptw_customCSRs_csrs_0_value  [3]&~  frontend__icache_io_s2_kill  )
            begin 
              if (1)$display("Assertion failed\n    at Frontend.scala:190 assert(!(s2_speculative && io.ptw.customCSRs.asInstanceOf[RocketCustomCSRs].disableSpeculativeICacheRefill && !icache.io.s2_kill))\n");
              if (1)$display("");
            end 
       end
  
  always @( posedge   frontend__clock  )
       begin  
          frontend__s1_valid   <=  frontend__s0_valid  ; 
          frontend__s1_pc   <={  frontend___io_cpu_npc_T  ,1'h0};
         if (  frontend__io_cpu_req_valid  ) 
             frontend__s1_speculative   <=  frontend__io_cpu_req_bits_speculative  ;
          else 
            if (  frontend__s2_replay  ) 
                frontend__s1_speculative   <=  frontend__s2_speculative  ;
             else  
                frontend__s1_speculative   <=  frontend__s1_speculative  |  frontend__s2_valid  &~  frontend__s2_speculative  ;
         if (~  frontend__s2_replay  )
            begin  
               frontend__s2_tlb_resp_pf_inst   <=  frontend___tlb_io_resp_pf_inst  ; 
               frontend__s2_tlb_resp_ae_inst   <=  frontend___tlb_io_resp_ae_inst  ; 
               frontend__s2_tlb_resp_cacheable   <=  frontend___tlb_io_resp_cacheable  ;
            end  
          frontend__fq_io_enq_valid_REG   <=  frontend__s1_valid  ;
         if (  frontend__reset  )
            begin  
               frontend__s2_valid   <=1'h0; 
               frontend__s2_pc   <=34'h10040; 
               frontend__s2_speculative   <=1'h0; 
               frontend__s2_replay_REG   <=1'h1;
            end 
          else 
            begin  
               frontend__s2_valid   <=~  frontend__s2_replay  &~  frontend__io_cpu_req_valid  ;
              if (~  frontend__s2_replay  )
                 begin  
                    frontend__s2_pc   <=  frontend__s1_pc  ; 
                    frontend__s2_speculative   <=  frontend__s1_speculative  ;
                 end  
               frontend__s2_replay_REG   <=  frontend__s2_replay  &~  frontend__s0_valid  ;
            end 
       end
   
  
wire  frontend__icache__clock;
wire  frontend__icache__reset;
wire  frontend__icache__auto_master_out_a_ready;
wire  frontend__icache__auto_master_out_a_valid;
wire [31:0] frontend__icache__auto_master_out_a_bits_address;
wire  frontend__icache__auto_master_out_d_valid;
wire [2:0] frontend__icache__auto_master_out_d_bits_opcode;
wire [3:0] frontend__icache__auto_master_out_d_bits_size;
wire [63:0] frontend__icache__auto_master_out_d_bits_data;
wire  frontend__icache__auto_master_out_d_bits_corrupt;
wire  frontend__icache__io_req_valid;
wire [32:0] frontend__icache__io_req_bits_addr;
wire [31:0] frontend__icache__io_s1_paddr;
wire  frontend__icache__io_s1_kill;
wire  frontend__icache__io_s2_kill;
wire  frontend__icache__io_resp_valid;
wire [31:0] frontend__icache__io_resp_bits_data;
wire  frontend__icache__io_resp_bits_ae;
wire  frontend__icache__io_invalidate;
 
   wire  frontend__icache__readEnable  ; 
   wire  frontend__icache__writeEnable  ; 
   wire  frontend__icache__readEnable_0  ; 
   wire  frontend__icache__wen  ; 
   wire  frontend__icache__readEnable_1  ; 
   wire[5:0]  frontend__icache___tag_rdata_T  ; 
   wire  frontend__icache__io_req_ready  ; 
   wire[31:0]  frontend__icache___data_arrays_1_0_ext_RW0_rdata  ; 
   wire[31:0]  frontend__icache___data_arrays_0_0_ext_RW0_rdata  ; 
   wire[20:0]  frontend__icache___tag_array_0_ext_RW0_rdata  ; 
   wire  frontend__icache__s0_valid  =  frontend__icache__io_req_ready  &  frontend__icache__io_req_valid  ; 
   reg  frontend__icache__s1_valid  ; 
   reg  frontend__icache__s2_valid  ; 
   reg  frontend__icache__s2_hit  ; 
   reg  frontend__icache__invalidated  ; 
   reg  frontend__icache__refill_valid  ; 
   wire  frontend__icache__s2_miss  =  frontend__icache__s2_valid  &~  frontend__icache__s2_hit  &~  frontend__icache__io_s2_kill  ; 
   reg  frontend__icache__s2_request_refill_REG  ; 
   wire  frontend__icache__s2_request_refill  =  frontend__icache__s2_miss  &  frontend__icache__s2_request_refill_REG  ; 
   reg[31:0]  frontend__icache__refill_paddr  ; 
   wire  frontend__icache__refill_one_beat  =  frontend__icache__auto_master_out_d_valid  &  frontend__icache__auto_master_out_d_bits_opcode  [0]; 
  assign   frontend__icache__io_req_ready  =~  frontend__icache__refill_one_beat  ; 
   wire[26:0]  frontend__icache___beats1_decode_T_1  =27'hFFF<<  frontend__icache__auto_master_out_d_bits_size  ; 
   wire[8:0]  frontend__icache__beats1  =  frontend__icache__auto_master_out_d_bits_opcode  [0] ? ~(  frontend__icache___beats1_decode_T_1  [11:3]):9'h0; 
   reg[8:0]  frontend__icache__counter  ; 
   wire[8:0]  frontend__icache___counter1_T  =  frontend__icache__counter  -9'h1; 
   wire[8:0]  frontend__icache__refill_cnt  =  frontend__icache__beats1  &~  frontend__icache___counter1_T  ; 
   wire  frontend__icache__writeEnable_0  =  frontend__icache__refill_one_beat  &(  frontend__icache__counter  ==9'h1|  frontend__icache__beats1  ==9'h0)&  frontend__icache__auto_master_out_d_valid  ; 
  assign   frontend__icache___tag_rdata_T  =  frontend__icache__io_req_bits_addr  [11:6]; 
  assign   frontend__icache__readEnable_1  =~  frontend__icache__writeEnable_0  &  frontend__icache__s0_valid  ; 
   reg  frontend__icache__accruedRefillError  ; 
   wire  frontend__icache__refillError  =  frontend__icache__auto_master_out_d_bits_corrupt  |(|  frontend__icache__refill_cnt  )&  frontend__icache__accruedRefillError  ; 
   reg[63:0]  frontend__icache__vb_array  ; 
   wire[63:0]  frontend__icache___s1_vb_T_1  =  frontend__icache__vb_array  >>  frontend__icache__io_s1_paddr  [11:6]; 
   wire  frontend__icache__s1_hit  =  frontend__icache___s1_vb_T_1  [0]&  frontend__icache___tag_array_0_ext_RW0_rdata  [19:0]==  frontend__icache__io_s1_paddr  [31:12]; 
  assign   frontend__icache__wen  =  frontend__icache__refill_one_beat  &~  frontend__icache__invalidated  ; 
   wire[8:0]  frontend__icache___mem_idx_T_6  ={  frontend__icache__refill_paddr  [11:6],3'h0}; 
  assign   frontend__icache__readEnable_0  =~  frontend__icache__wen  &  frontend__icache__s0_valid  &~(  frontend__icache__io_req_bits_addr  [2]); 
  assign   frontend__icache__writeEnable  =  frontend__icache__refill_one_beat  &~  frontend__icache__invalidated  ; 
  assign   frontend__icache__readEnable  =~  frontend__icache__writeEnable  &  frontend__icache__s0_valid  &  frontend__icache__io_req_bits_addr  [2]; 
   reg[31:0]  frontend__icache__s2_dout_0  ; 
   reg  frontend__icache__s2_tl_error  ; 
   wire[127:0]  frontend__icache___vb_array_T_3  =128'h1<<  frontend__icache__refill_paddr  [11:6]; 
   wire  frontend__icache___s1_can_request_refill_T  =  frontend__icache__s2_miss  |  frontend__icache__refill_valid  ; 
  always @( posedge   frontend__icache__clock  )
       begin 
         if (  frontend__icache__reset  )
            begin  
               frontend__icache__s1_valid   <=1'h0; 
               frontend__icache__s2_valid   <=1'h0; 
               frontend__icache__refill_valid   <=1'h0; 
               frontend__icache__counter   <=9'h0; 
               frontend__icache__vb_array   <=64'h0;
            end 
          else 
            begin  
               frontend__icache__s1_valid   <=  frontend__icache__s0_valid  ; 
               frontend__icache__s2_valid   <=  frontend__icache__s1_valid  &~  frontend__icache__io_s1_kill  ; 
               frontend__icache__refill_valid   <=~  frontend__icache__writeEnable_0  &(  frontend__icache__auto_master_out_a_ready  &  frontend__icache__s2_request_refill  |  frontend__icache__refill_valid  );
              if (  frontend__icache__auto_master_out_d_valid  )
                 begin 
                   if (  frontend__icache__counter  ==9'h0) 
                       frontend__icache__counter   <=  frontend__icache__beats1  ;
                    else  
                       frontend__icache__counter   <=  frontend__icache___counter1_T  ;
                 end 
              if (  frontend__icache__io_invalidate  ) 
                  frontend__icache__vb_array   <=64'h0;
               else 
                 if (  frontend__icache__refill_one_beat  ) 
                     frontend__icache__vb_array   <=  frontend__icache__writeEnable_0  &~  frontend__icache__invalidated   ?   frontend__icache__vb_array  |  frontend__icache___vb_array_T_3  [63:0]:~(~  frontend__icache__vb_array  |  frontend__icache___vb_array_T_3  [63:0]);
            end  
          frontend__icache__s2_hit   <=  frontend__icache__s1_hit  ; 
          frontend__icache__invalidated   <=  frontend__icache__refill_valid  &(  frontend__icache__io_invalidate  |  frontend__icache__invalidated  ); 
          frontend__icache__s2_request_refill_REG   <=~  frontend__icache___s1_can_request_refill_T  ;
         if (  frontend__icache__s1_valid  &~  frontend__icache___s1_can_request_refill_T  ) 
             frontend__icache__refill_paddr   <=  frontend__icache__io_s1_paddr  ;
         if (  frontend__icache__refill_one_beat  ) 
             frontend__icache__accruedRefillError   <=  frontend__icache__refillError  ;
         if (  frontend__icache__s1_valid  )
            begin  
               frontend__icache__s2_dout_0   <=  frontend__icache__io_s1_paddr  [2] ?   frontend__icache___data_arrays_1_0_ext_RW0_rdata  :  frontend__icache___data_arrays_0_0_ext_RW0_rdata  ; 
               frontend__icache__s2_tl_error   <=  frontend__icache__s1_hit  &  frontend__icache___tag_array_0_ext_RW0_rdata  [20];
            end 
       end
   
  
wire [5:0] frontend__icache__tag_array_0_ext__RW0_addr;
wire  frontend__icache__tag_array_0_ext__RW0_en;
wire  frontend__icache__tag_array_0_ext__RW0_clk;
wire  frontend__icache__tag_array_0_ext__RW0_wmode;
wire [20:0] frontend__icache__tag_array_0_ext__RW0_wdata;
wire [20:0] frontend__icache__tag_array_0_ext__RW0_rdata;
 
   reg[20:0]  frontend__icache__tag_array_0_ext__Memory  [0:63]; 
   reg[5:0]  frontend__icache__tag_array_0_ext___RW0_raddr_d0  ; 
   reg  frontend__icache__tag_array_0_ext___RW0_ren_d0  ; 
   reg  frontend__icache__tag_array_0_ext___RW0_rmode_d0  ; 
  always @( posedge   frontend__icache__tag_array_0_ext__RW0_clk  )
       begin  
          frontend__icache__tag_array_0_ext___RW0_raddr_d0   <=  frontend__icache__tag_array_0_ext__RW0_addr  ; 
          frontend__icache__tag_array_0_ext___RW0_ren_d0   <=  frontend__icache__tag_array_0_ext__RW0_en  ; 
          frontend__icache__tag_array_0_ext___RW0_rmode_d0   <=  frontend__icache__tag_array_0_ext__RW0_wmode  ;
         if (  frontend__icache__tag_array_0_ext__RW0_en  &  frontend__icache__tag_array_0_ext__RW0_wmode  &1'h1) 
             frontend__icache__tag_array_0_ext__Memory   [  frontend__icache__tag_array_0_ext__RW0_addr  ]<=  frontend__icache__tag_array_0_ext__RW0_wdata  ;
       end
  
  assign   frontend__icache__tag_array_0_ext__RW0_rdata  =  frontend__icache__tag_array_0_ext___RW0_ren_d0  &~  frontend__icache__tag_array_0_ext___RW0_rmode_d0   ?   frontend__icache__tag_array_0_ext__Memory  [  frontend__icache__tag_array_0_ext___RW0_raddr_d0  ]:21'bx;
assign frontend__icache__tag_array_0_ext__RW0_addr = frontend__icache__writeEnable_0 ? frontend__icache__refill_paddr[11:6]:frontend__icache___tag_rdata_T;
assign frontend__icache__tag_array_0_ext__RW0_en = frontend__icache__readEnable_1|frontend__icache__writeEnable_0;
assign frontend__icache__tag_array_0_ext__RW0_clk = frontend__icache__clock;
assign frontend__icache__tag_array_0_ext__RW0_wmode = frontend__icache__refill_one_beat;
assign frontend__icache__tag_array_0_ext__RW0_wdata = {frontend__icache__refillError,frontend__icache__refill_paddr[31:12]};
assign frontend__icache___tag_array_0_ext_RW0_rdata = frontend__icache__tag_array_0_ext__RW0_rdata;
  
  
wire [8:0] frontend__icache__data_arrays_0_0_ext__RW0_addr;
wire  frontend__icache__data_arrays_0_0_ext__RW0_en;
wire  frontend__icache__data_arrays_0_0_ext__RW0_clk;
wire  frontend__icache__data_arrays_0_0_ext__RW0_wmode;
wire [31:0] frontend__icache__data_arrays_0_0_ext__RW0_wdata;
wire [31:0] frontend__icache__data_arrays_0_0_ext__RW0_rdata;
wire [8:0] frontend__icache__data_arrays_1_0_ext__RW0_addr;
wire  frontend__icache__data_arrays_1_0_ext__RW0_en;
wire  frontend__icache__data_arrays_1_0_ext__RW0_clk;
wire  frontend__icache__data_arrays_1_0_ext__RW0_wmode;
wire [31:0] frontend__icache__data_arrays_1_0_ext__RW0_wdata;
wire [31:0] frontend__icache__data_arrays_1_0_ext__RW0_rdata;
 
   reg[31:0]  frontend__icache__data_arrays_0_0_ext__Memory  [0:511]; 
   reg[8:0]  frontend__icache__data_arrays_0_0_ext___RW0_raddr_d0  ; 
   reg  frontend__icache__data_arrays_0_0_ext___RW0_ren_d0  ; 
   reg  frontend__icache__data_arrays_0_0_ext___RW0_rmode_d0  ; 
  always @( posedge   frontend__icache__data_arrays_0_0_ext__RW0_clk  )
       begin  
          frontend__icache__data_arrays_0_0_ext___RW0_raddr_d0   <=  frontend__icache__data_arrays_0_0_ext__RW0_addr  ; 
          frontend__icache__data_arrays_0_0_ext___RW0_ren_d0   <=  frontend__icache__data_arrays_0_0_ext__RW0_en  ; 
          frontend__icache__data_arrays_0_0_ext___RW0_rmode_d0   <=  frontend__icache__data_arrays_0_0_ext__RW0_wmode  ;
         if (  frontend__icache__data_arrays_0_0_ext__RW0_en  &  frontend__icache__data_arrays_0_0_ext__RW0_wmode  &1'h1) 
             frontend__icache__data_arrays_0_0_ext__Memory   [  frontend__icache__data_arrays_0_0_ext__RW0_addr  ]<=  frontend__icache__data_arrays_0_0_ext__RW0_wdata  ;
       end
  
  assign   frontend__icache__data_arrays_0_0_ext__RW0_rdata  =  frontend__icache__data_arrays_0_0_ext___RW0_ren_d0  &~  frontend__icache__data_arrays_0_0_ext___RW0_rmode_d0   ?   frontend__icache__data_arrays_0_0_ext__Memory  [  frontend__icache__data_arrays_0_0_ext___RW0_raddr_d0  ]:32'bx;
  
  
 
   reg[31:0]  frontend__icache__data_arrays_1_0_ext__Memory  [0:511]; 
   reg[8:0]  frontend__icache__data_arrays_1_0_ext___RW0_raddr_d0  ; 
   reg  frontend__icache__data_arrays_1_0_ext___RW0_ren_d0  ; 
   reg  frontend__icache__data_arrays_1_0_ext___RW0_rmode_d0  ; 
  always @( posedge   frontend__icache__data_arrays_1_0_ext__RW0_clk  )
       begin  
          frontend__icache__data_arrays_1_0_ext___RW0_raddr_d0   <=  frontend__icache__data_arrays_1_0_ext__RW0_addr  ; 
          frontend__icache__data_arrays_1_0_ext___RW0_ren_d0   <=  frontend__icache__data_arrays_1_0_ext__RW0_en  ; 
          frontend__icache__data_arrays_1_0_ext___RW0_rmode_d0   <=  frontend__icache__data_arrays_1_0_ext__RW0_wmode  ;
         if (  frontend__icache__data_arrays_1_0_ext__RW0_en  &  frontend__icache__data_arrays_1_0_ext__RW0_wmode  &1'h1) 
             frontend__icache__data_arrays_1_0_ext__Memory   [  frontend__icache__data_arrays_1_0_ext__RW0_addr  ]<=  frontend__icache__data_arrays_1_0_ext__RW0_wdata  ;
       end
  
  assign   frontend__icache__data_arrays_1_0_ext__RW0_rdata  =  frontend__icache__data_arrays_1_0_ext___RW0_ren_d0  &~  frontend__icache__data_arrays_1_0_ext___RW0_rmode_d0   ?   frontend__icache__data_arrays_1_0_ext__Memory  [  frontend__icache__data_arrays_1_0_ext___RW0_raddr_d0  ]:32'bx;
assign frontend__icache__data_arrays_0_0_ext__RW0_addr = frontend__icache__refill_one_beat ? frontend__icache___mem_idx_T_6|frontend__icache__refill_cnt:frontend__icache__io_req_bits_addr[11:3];
assign frontend__icache__data_arrays_0_0_ext__RW0_en = frontend__icache__readEnable_0|frontend__icache__wen;
assign frontend__icache__data_arrays_0_0_ext__RW0_clk = frontend__icache__clock;
assign frontend__icache__data_arrays_0_0_ext__RW0_wmode = frontend__icache__refill_one_beat;
assign frontend__icache__data_arrays_0_0_ext__RW0_wdata = frontend__icache__auto_master_out_d_bits_data[31:0];
assign frontend__icache___data_arrays_0_0_ext_RW0_rdata = frontend__icache__data_arrays_0_0_ext__RW0_rdata;
assign frontend__icache__data_arrays_1_0_ext__RW0_addr = frontend__icache__refill_one_beat ? frontend__icache___mem_idx_T_6|frontend__icache__refill_cnt:frontend__icache__io_req_bits_addr[11:3];
assign frontend__icache__data_arrays_1_0_ext__RW0_en = frontend__icache__readEnable|frontend__icache__writeEnable;
assign frontend__icache__data_arrays_1_0_ext__RW0_clk = frontend__icache__clock;
assign frontend__icache__data_arrays_1_0_ext__RW0_wmode = frontend__icache__refill_one_beat;
assign frontend__icache__data_arrays_1_0_ext__RW0_wdata = frontend__icache__auto_master_out_d_bits_data[63:32];
assign frontend__icache___data_arrays_1_0_ext_RW0_rdata = frontend__icache__data_arrays_1_0_ext__RW0_rdata;
 
  assign   frontend__icache__auto_master_out_a_valid  =  frontend__icache__s2_request_refill  ; 
  assign   frontend__icache__auto_master_out_a_bits_address  ={  frontend__icache__refill_paddr  [31:6],6'h0}; 
  assign   frontend__icache__io_resp_valid  =  frontend__icache__s2_valid  &  frontend__icache__s2_hit  ; 
  assign   frontend__icache__io_resp_bits_data  =  frontend__icache__s2_dout_0  ; 
  assign   frontend__icache__io_resp_bits_ae  =  frontend__icache__s2_tl_error  ;
assign frontend__icache__clock = frontend__clock;
assign frontend__icache__reset = frontend__reset;
assign frontend__icache__auto_master_out_a_ready = frontend__auto_icache_master_out_a_ready;
assign frontend__auto_icache_master_out_a_valid = frontend__icache__auto_master_out_a_valid;
assign frontend__auto_icache_master_out_a_bits_address = frontend__icache__auto_master_out_a_bits_address;
assign frontend__icache__auto_master_out_d_valid = frontend__auto_icache_master_out_d_valid;
assign frontend__icache__auto_master_out_d_bits_opcode = frontend__auto_icache_master_out_d_bits_opcode;
assign frontend__icache__auto_master_out_d_bits_size = frontend__auto_icache_master_out_d_bits_size;
assign frontend__icache__auto_master_out_d_bits_data = frontend__auto_icache_master_out_d_bits_data;
assign frontend__icache__auto_master_out_d_bits_corrupt = frontend__auto_icache_master_out_d_bits_corrupt;
assign frontend__icache__io_req_valid = frontend__s0_valid;
assign frontend__icache__io_req_bits_addr = {frontend___io_cpu_npc_T[31:0],1'h0};
assign frontend__icache__io_s1_paddr = frontend___tlb_io_resp_paddr;
assign frontend__icache__io_s1_kill = frontend__io_cpu_req_valid|frontend__s2_replay;
assign frontend__icache__io_s2_kill = frontend__icache_io_s2_kill;
assign frontend___icache_io_resp_valid = frontend__icache__io_resp_valid;
assign frontend___icache_io_resp_bits_data = frontend__icache__io_resp_bits_data;
assign frontend___icache_io_resp_bits_ae = frontend__icache__io_resp_bits_ae;
assign frontend__icache__io_invalidate = frontend__io_cpu_flush_icache;
  
  
wire  frontend__fq__clock;
wire  frontend__fq__reset;
wire  frontend__fq__io_enq_ready;
wire  frontend__fq__io_enq_valid;
wire [33:0] frontend__fq__io_enq_bits_pc;
wire [31:0] frontend__fq__io_enq_bits_data;
wire  frontend__fq__io_enq_bits_xcpt_pf_inst;
wire  frontend__fq__io_enq_bits_xcpt_ae_inst;
wire  frontend__fq__io_enq_bits_replay;
wire  frontend__fq__io_deq_ready;
wire  frontend__fq__io_deq_valid;
wire [33:0] frontend__fq__io_deq_bits_pc;
wire [31:0] frontend__fq__io_deq_bits_data;
wire  frontend__fq__io_deq_bits_xcpt_pf_inst;
wire  frontend__fq__io_deq_bits_xcpt_gf_inst;
wire  frontend__fq__io_deq_bits_xcpt_ae_inst;
wire  frontend__fq__io_deq_bits_replay;
wire [4:0] frontend__fq__io_mask;
 
   reg  frontend__fq__valid_0  ; 
   reg  frontend__fq__valid_1  ; 
   reg  frontend__fq__valid_2  ; 
   reg  frontend__fq__valid_3  ; 
   reg  frontend__fq__valid_4  ; 
   reg[33:0]  frontend__fq__elts_pc_0  ; 
   reg[33:0]  frontend__fq__elts_pc_1  ; 
   reg[33:0]  frontend__fq__elts_pc_2  ; 
   reg[33:0]  frontend__fq__elts_pc_3  ; 
   reg[33:0]  frontend__fq__elts_pc_4  ; 
   reg[31:0]  frontend__fq__elts_data_0  ; 
   reg[31:0]  frontend__fq__elts_data_1  ; 
   reg[31:0]  frontend__fq__elts_data_2  ; 
   reg[31:0]  frontend__fq__elts_data_3  ; 
   reg[31:0]  frontend__fq__elts_data_4  ; 
   reg  frontend__fq__elts_xcpt_pf_inst_0  ; 
   reg  frontend__fq__elts_xcpt_pf_inst_1  ; 
   reg  frontend__fq__elts_xcpt_pf_inst_2  ; 
   reg  frontend__fq__elts_xcpt_pf_inst_3  ; 
   reg  frontend__fq__elts_xcpt_pf_inst_4  ; 
   reg  frontend__fq__elts_xcpt_gf_inst_0  ; 
   reg  frontend__fq__elts_xcpt_gf_inst_1  ; 
   reg  frontend__fq__elts_xcpt_gf_inst_2  ; 
   reg  frontend__fq__elts_xcpt_gf_inst_3  ; 
   reg  frontend__fq__elts_xcpt_gf_inst_4  ; 
   reg  frontend__fq__elts_xcpt_ae_inst_0  ; 
   reg  frontend__fq__elts_xcpt_ae_inst_1  ; 
   reg  frontend__fq__elts_xcpt_ae_inst_2  ; 
   reg  frontend__fq__elts_xcpt_ae_inst_3  ; 
   reg  frontend__fq__elts_xcpt_ae_inst_4  ; 
   reg  frontend__fq__elts_replay_0  ; 
   reg  frontend__fq__elts_replay_1  ; 
   reg  frontend__fq__elts_replay_2  ; 
   reg  frontend__fq__elts_replay_3  ; 
   reg  frontend__fq__elts_replay_4  ; 
   wire  frontend__fq___valid_4_T_4  =~  frontend__fq__valid_4  &  frontend__fq__io_enq_valid  ; 
   wire  frontend__fq__wen_4  =  frontend__fq__io_deq_ready   ?   frontend__fq___valid_4_T_4  &  frontend__fq__valid_4  :  frontend__fq___valid_4_T_4  &  frontend__fq__valid_3  &~  frontend__fq__valid_4  ; 
  always @( posedge   frontend__fq__clock  )
       begin 
         if (  frontend__fq__reset  )
            begin  
               frontend__fq__valid_0   <=1'h0; 
               frontend__fq__valid_1   <=1'h0; 
               frontend__fq__valid_2   <=1'h0; 
               frontend__fq__valid_3   <=1'h0; 
               frontend__fq__valid_4   <=1'h0;
            end 
          else 
            if (  frontend__fq__io_deq_ready  )
               begin  
                  frontend__fq__valid_0   <=  frontend__fq__valid_1  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_0  ; 
                  frontend__fq__valid_1   <=  frontend__fq__valid_2  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_1  ; 
                  frontend__fq__valid_2   <=  frontend__fq__valid_3  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_2  ; 
                  frontend__fq__valid_3   <=  frontend__fq__valid_4  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_3  ; 
                  frontend__fq__valid_4   <=  frontend__fq___valid_4_T_4  &  frontend__fq__valid_4  ;
               end 
             else 
               begin  
                  frontend__fq__valid_0   <=  frontend__fq___valid_4_T_4  |  frontend__fq__valid_0  ; 
                  frontend__fq__valid_1   <=  frontend__fq___valid_4_T_4  &  frontend__fq__valid_0  |  frontend__fq__valid_1  ; 
                  frontend__fq__valid_2   <=  frontend__fq___valid_4_T_4  &  frontend__fq__valid_1  |  frontend__fq__valid_2  ; 
                  frontend__fq__valid_3   <=  frontend__fq___valid_4_T_4  &  frontend__fq__valid_2  |  frontend__fq__valid_3  ; 
                  frontend__fq__valid_4   <=  frontend__fq___valid_4_T_4  &  frontend__fq__valid_3  |  frontend__fq__valid_4  ;
               end 
         if (  frontend__fq__io_deq_ready   ?   frontend__fq__valid_1  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_0  :  frontend__fq___valid_4_T_4  &~  frontend__fq__valid_0  )
            begin  
               frontend__fq__elts_pc_0   <=  frontend__fq__valid_1   ?   frontend__fq__elts_pc_1  :  frontend__fq__io_enq_bits_pc  ; 
               frontend__fq__elts_data_0   <=  frontend__fq__valid_1   ?   frontend__fq__elts_data_1  :  frontend__fq__io_enq_bits_data  ; 
               frontend__fq__elts_xcpt_pf_inst_0   <=  frontend__fq__valid_1   ?   frontend__fq__elts_xcpt_pf_inst_1  :  frontend__fq__io_enq_bits_xcpt_pf_inst  ; 
               frontend__fq__elts_xcpt_gf_inst_0   <=  frontend__fq__valid_1  &  frontend__fq__elts_xcpt_gf_inst_1  ; 
               frontend__fq__elts_xcpt_ae_inst_0   <=  frontend__fq__valid_1   ?   frontend__fq__elts_xcpt_ae_inst_1  :  frontend__fq__io_enq_bits_xcpt_ae_inst  ; 
               frontend__fq__elts_replay_0   <=  frontend__fq__valid_1   ?   frontend__fq__elts_replay_1  :  frontend__fq__io_enq_bits_replay  ;
            end 
         if (  frontend__fq__io_deq_ready   ?   frontend__fq__valid_2  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_1  :  frontend__fq___valid_4_T_4  &  frontend__fq__valid_0  &~  frontend__fq__valid_1  )
            begin  
               frontend__fq__elts_pc_1   <=  frontend__fq__valid_2   ?   frontend__fq__elts_pc_2  :  frontend__fq__io_enq_bits_pc  ; 
               frontend__fq__elts_data_1   <=  frontend__fq__valid_2   ?   frontend__fq__elts_data_2  :  frontend__fq__io_enq_bits_data  ; 
               frontend__fq__elts_xcpt_pf_inst_1   <=  frontend__fq__valid_2   ?   frontend__fq__elts_xcpt_pf_inst_2  :  frontend__fq__io_enq_bits_xcpt_pf_inst  ; 
               frontend__fq__elts_xcpt_gf_inst_1   <=  frontend__fq__valid_2  &  frontend__fq__elts_xcpt_gf_inst_2  ; 
               frontend__fq__elts_xcpt_ae_inst_1   <=  frontend__fq__valid_2   ?   frontend__fq__elts_xcpt_ae_inst_2  :  frontend__fq__io_enq_bits_xcpt_ae_inst  ; 
               frontend__fq__elts_replay_1   <=  frontend__fq__valid_2   ?   frontend__fq__elts_replay_2  :  frontend__fq__io_enq_bits_replay  ;
            end 
         if (  frontend__fq__io_deq_ready   ?   frontend__fq__valid_3  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_2  :  frontend__fq___valid_4_T_4  &  frontend__fq__valid_1  &~  frontend__fq__valid_2  )
            begin  
               frontend__fq__elts_pc_2   <=  frontend__fq__valid_3   ?   frontend__fq__elts_pc_3  :  frontend__fq__io_enq_bits_pc  ; 
               frontend__fq__elts_data_2   <=  frontend__fq__valid_3   ?   frontend__fq__elts_data_3  :  frontend__fq__io_enq_bits_data  ; 
               frontend__fq__elts_xcpt_pf_inst_2   <=  frontend__fq__valid_3   ?   frontend__fq__elts_xcpt_pf_inst_3  :  frontend__fq__io_enq_bits_xcpt_pf_inst  ; 
               frontend__fq__elts_xcpt_gf_inst_2   <=  frontend__fq__valid_3  &  frontend__fq__elts_xcpt_gf_inst_3  ; 
               frontend__fq__elts_xcpt_ae_inst_2   <=  frontend__fq__valid_3   ?   frontend__fq__elts_xcpt_ae_inst_3  :  frontend__fq__io_enq_bits_xcpt_ae_inst  ; 
               frontend__fq__elts_replay_2   <=  frontend__fq__valid_3   ?   frontend__fq__elts_replay_3  :  frontend__fq__io_enq_bits_replay  ;
            end 
         if (  frontend__fq__io_deq_ready   ?   frontend__fq__valid_4  |  frontend__fq___valid_4_T_4  &  frontend__fq__valid_3  :  frontend__fq___valid_4_T_4  &  frontend__fq__valid_2  &~  frontend__fq__valid_3  )
            begin  
               frontend__fq__elts_pc_3   <=  frontend__fq__valid_4   ?   frontend__fq__elts_pc_4  :  frontend__fq__io_enq_bits_pc  ; 
               frontend__fq__elts_data_3   <=  frontend__fq__valid_4   ?   frontend__fq__elts_data_4  :  frontend__fq__io_enq_bits_data  ; 
               frontend__fq__elts_xcpt_pf_inst_3   <=  frontend__fq__valid_4   ?   frontend__fq__elts_xcpt_pf_inst_4  :  frontend__fq__io_enq_bits_xcpt_pf_inst  ; 
               frontend__fq__elts_xcpt_gf_inst_3   <=  frontend__fq__valid_4  &  frontend__fq__elts_xcpt_gf_inst_4  ; 
               frontend__fq__elts_xcpt_ae_inst_3   <=  frontend__fq__valid_4   ?   frontend__fq__elts_xcpt_ae_inst_4  :  frontend__fq__io_enq_bits_xcpt_ae_inst  ; 
               frontend__fq__elts_replay_3   <=  frontend__fq__valid_4   ?   frontend__fq__elts_replay_4  :  frontend__fq__io_enq_bits_replay  ;
            end 
         if (  frontend__fq__wen_4  )
            begin  
               frontend__fq__elts_pc_4   <=  frontend__fq__io_enq_bits_pc  ; 
               frontend__fq__elts_data_4   <=  frontend__fq__io_enq_bits_data  ; 
               frontend__fq__elts_xcpt_pf_inst_4   <=  frontend__fq__io_enq_bits_xcpt_pf_inst  ; 
               frontend__fq__elts_xcpt_ae_inst_4   <=  frontend__fq__io_enq_bits_xcpt_ae_inst  ; 
               frontend__fq__elts_replay_4   <=  frontend__fq__io_enq_bits_replay  ;
            end  
          frontend__fq__elts_xcpt_gf_inst_4   <=~  frontend__fq__wen_4  &  frontend__fq__elts_xcpt_gf_inst_4  ;
       end
  
  assign   frontend__fq__io_enq_ready  =~  frontend__fq__valid_4  ; 
  assign   frontend__fq__io_deq_valid  =  frontend__fq__io_enq_valid  |  frontend__fq__valid_0  ; 
  assign   frontend__fq__io_deq_bits_pc  =  frontend__fq__valid_0   ?   frontend__fq__elts_pc_0  :  frontend__fq__io_enq_bits_pc  ; 
  assign   frontend__fq__io_deq_bits_data  =  frontend__fq__valid_0   ?   frontend__fq__elts_data_0  :  frontend__fq__io_enq_bits_data  ; 
  assign   frontend__fq__io_deq_bits_xcpt_pf_inst  =  frontend__fq__valid_0   ?   frontend__fq__elts_xcpt_pf_inst_0  :  frontend__fq__io_enq_bits_xcpt_pf_inst  ; 
  assign   frontend__fq__io_deq_bits_xcpt_gf_inst  =  frontend__fq__valid_0  &  frontend__fq__elts_xcpt_gf_inst_0  ; 
  assign   frontend__fq__io_deq_bits_xcpt_ae_inst  =  frontend__fq__valid_0   ?   frontend__fq__elts_xcpt_ae_inst_0  :  frontend__fq__io_enq_bits_xcpt_ae_inst  ; 
  assign   frontend__fq__io_deq_bits_replay  =  frontend__fq__valid_0   ?   frontend__fq__elts_replay_0  :  frontend__fq__io_enq_bits_replay  ; 
  assign   frontend__fq__io_mask  ={  frontend__fq__valid_4  ,  frontend__fq__valid_3  ,  frontend__fq__valid_2  ,  frontend__fq__valid_1  ,  frontend__fq__valid_0  };
assign frontend__fq__clock = frontend__clock;
assign frontend__fq__reset = frontend__reset|frontend__io_cpu_req_valid;
assign frontend___fq_io_enq_ready = frontend__fq__io_enq_ready;
assign frontend__fq__io_enq_valid = frontend__fq_io_enq_valid;
assign frontend__fq__io_enq_bits_pc = frontend__s2_pc;
assign frontend__fq__io_enq_bits_data = frontend___icache_io_resp_bits_data;
assign frontend__fq__io_enq_bits_xcpt_pf_inst = frontend__s2_tlb_resp_pf_inst;
assign frontend__fq__io_enq_bits_xcpt_ae_inst = frontend___icache_io_resp_valid&frontend___icache_io_resp_bits_ae|frontend__s2_tlb_resp_ae_inst;
assign frontend__fq__io_enq_bits_replay = frontend__icache_io_s2_kill&~frontend___icache_io_resp_valid&~frontend___s2_xcpt_T;
assign frontend__fq__io_deq_ready = frontend__io_cpu_resp_ready;
assign frontend__io_cpu_resp_valid = frontend__fq__io_deq_valid;
assign frontend__io_cpu_resp_bits_pc = frontend__fq__io_deq_bits_pc;
assign frontend__io_cpu_resp_bits_data = frontend__fq__io_deq_bits_data;
assign frontend__io_cpu_resp_bits_xcpt_pf_inst = frontend__fq__io_deq_bits_xcpt_pf_inst;
assign frontend__io_cpu_resp_bits_xcpt_gf_inst = frontend__fq__io_deq_bits_xcpt_gf_inst;
assign frontend__io_cpu_resp_bits_xcpt_ae_inst = frontend__fq__io_deq_bits_xcpt_ae_inst;
assign frontend__io_cpu_resp_bits_replay = frontend__fq__io_deq_bits_replay;
assign frontend___fq_io_mask = frontend__fq__io_mask;
  
  
wire [33:0] frontend__tlb__io_req_bits_vaddr;
wire [31:0] frontend__tlb__io_resp_paddr;
wire  frontend__tlb__io_resp_pf_inst;
wire  frontend__tlb__io_resp_ae_inst;
wire  frontend__tlb__io_resp_cacheable;
wire  frontend__tlb__io_ptw_req_bits_bits_need_gpa;
wire  frontend__tlb__io_ptw_req_bits_bits_stage2;
wire  frontend__tlb__io_ptw_status_debug;
wire  frontend__tlb__io_ptw_pmp_cfg_l_0;
wire  frontend__tlb__io_ptw_pmp_cfg_l_1;
wire  frontend__tlb__io_ptw_pmp_cfg_l_2;
wire  frontend__tlb__io_ptw_pmp_cfg_l_3;
wire  frontend__tlb__io_ptw_pmp_cfg_l_4;
wire  frontend__tlb__io_ptw_pmp_cfg_l_5;
wire  frontend__tlb__io_ptw_pmp_cfg_l_6;
wire  frontend__tlb__io_ptw_pmp_cfg_l_7;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_0;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_1;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_2;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_3;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_4;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_5;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_6;
wire [1:0] frontend__tlb__io_ptw_pmp_cfg_a_7;
wire  frontend__tlb__io_ptw_pmp_cfg_x_0;
wire  frontend__tlb__io_ptw_pmp_cfg_x_1;
wire  frontend__tlb__io_ptw_pmp_cfg_x_2;
wire  frontend__tlb__io_ptw_pmp_cfg_x_3;
wire  frontend__tlb__io_ptw_pmp_cfg_x_4;
wire  frontend__tlb__io_ptw_pmp_cfg_x_5;
wire  frontend__tlb__io_ptw_pmp_cfg_x_6;
wire  frontend__tlb__io_ptw_pmp_cfg_x_7;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_0;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_1;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_2;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_3;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_4;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_5;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_6;
wire [29:0] frontend__tlb__io_ptw_pmp_addr_7;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_0;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_1;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_2;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_3;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_4;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_5;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_6;
wire [31:0] frontend__tlb__io_ptw_pmp_mask_7;
 
   wire  frontend__tlb___pmp_io_x  ; 
   wire[3:0]  frontend__tlb___GEN  =  frontend__tlb__io_req_bits_vaddr  [31:28]^4'h8; 
   wire  frontend__tlb__legal_address  ={  frontend__tlb__io_req_bits_vaddr  [33:14],~(  frontend__tlb__io_req_bits_vaddr  [13:12])}==22'h0|{  frontend__tlb__io_req_bits_vaddr  [33:28],~(  frontend__tlb__io_req_bits_vaddr  [27:26])}==8'h0|{  frontend__tlb__io_req_bits_vaddr  [33:26],  frontend__tlb__io_req_bits_vaddr  [25:16]^10'h200}==18'h0|~(|(  frontend__tlb__io_req_bits_vaddr  [33:12]))|{  frontend__tlb__io_req_bits_vaddr  [33:17],~(  frontend__tlb__io_req_bits_vaddr  [16])}==18'h0|{  frontend__tlb__io_req_bits_vaddr  [33:32],  frontend__tlb___GEN  }==6'h0|{  frontend__tlb__io_req_bits_vaddr  [33:31],~(  frontend__tlb__io_req_bits_vaddr  [30:29])}==5'h0;  
  
wire [1:0] frontend__tlb__pmp__io_prv;
wire  frontend__tlb__pmp__io_pmp_cfg_l_0;
wire  frontend__tlb__pmp__io_pmp_cfg_l_1;
wire  frontend__tlb__pmp__io_pmp_cfg_l_2;
wire  frontend__tlb__pmp__io_pmp_cfg_l_3;
wire  frontend__tlb__pmp__io_pmp_cfg_l_4;
wire  frontend__tlb__pmp__io_pmp_cfg_l_5;
wire  frontend__tlb__pmp__io_pmp_cfg_l_6;
wire  frontend__tlb__pmp__io_pmp_cfg_l_7;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_0;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_1;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_2;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_3;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_4;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_5;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_6;
wire [1:0] frontend__tlb__pmp__io_pmp_cfg_a_7;
wire  frontend__tlb__pmp__io_pmp_cfg_x_0;
wire  frontend__tlb__pmp__io_pmp_cfg_x_1;
wire  frontend__tlb__pmp__io_pmp_cfg_x_2;
wire  frontend__tlb__pmp__io_pmp_cfg_x_3;
wire  frontend__tlb__pmp__io_pmp_cfg_x_4;
wire  frontend__tlb__pmp__io_pmp_cfg_x_5;
wire  frontend__tlb__pmp__io_pmp_cfg_x_6;
wire  frontend__tlb__pmp__io_pmp_cfg_x_7;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_0;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_1;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_2;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_3;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_4;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_5;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_6;
wire [29:0] frontend__tlb__pmp__io_pmp_addr_7;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_0;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_1;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_2;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_3;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_4;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_5;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_6;
wire [31:0] frontend__tlb__pmp__io_pmp_mask_7;
wire [31:0] frontend__tlb__pmp__io_addr;
wire  frontend__tlb__pmp__io_x;
 
  assign   frontend__tlb__pmp__io_x  =(  frontend__tlb__pmp__io_pmp_cfg_a_0  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_0  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_0  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_0  [0]&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_0  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_0  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_0  :(  frontend__tlb__pmp__io_pmp_cfg_a_1  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_1  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_1  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_1  [0]&  frontend__tlb__pmp__io_addr  >={  frontend__tlb__pmp__io_pmp_addr_0  ,2'h0}&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_1  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_1  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_1  :(  frontend__tlb__pmp__io_pmp_cfg_a_2  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_2  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_2  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_2  [0]&  frontend__tlb__pmp__io_addr  >={  frontend__tlb__pmp__io_pmp_addr_1  ,2'h0}&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_2  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_2  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_2  :(  frontend__tlb__pmp__io_pmp_cfg_a_3  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_3  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_3  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_3  [0]&  frontend__tlb__pmp__io_addr  >={  frontend__tlb__pmp__io_pmp_addr_2  ,2'h0}&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_3  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_3  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_3  :(  frontend__tlb__pmp__io_pmp_cfg_a_4  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_4  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_4  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_4  [0]&  frontend__tlb__pmp__io_addr  >={  frontend__tlb__pmp__io_pmp_addr_3  ,2'h0}&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_4  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_4  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_4  :(  frontend__tlb__pmp__io_pmp_cfg_a_5  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_5  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_5  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_5  [0]&  frontend__tlb__pmp__io_addr  >={  frontend__tlb__pmp__io_pmp_addr_4  ,2'h0}&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_5  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_5  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_5  :(  frontend__tlb__pmp__io_pmp_cfg_a_6  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_6  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_6  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_6  [0]&  frontend__tlb__pmp__io_addr  >={  frontend__tlb__pmp__io_pmp_addr_5  ,2'h0}&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_6  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_6  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_6  :(  frontend__tlb__pmp__io_pmp_cfg_a_7  [1] ? ((  frontend__tlb__pmp__io_addr  ^{  frontend__tlb__pmp__io_pmp_addr_7  ,2'h0})&~  frontend__tlb__pmp__io_pmp_mask_7  )==32'h0:  frontend__tlb__pmp__io_pmp_cfg_a_7  [0]&  frontend__tlb__pmp__io_addr  >={  frontend__tlb__pmp__io_pmp_addr_6  ,2'h0}&  frontend__tlb__pmp__io_addr  <{  frontend__tlb__pmp__io_pmp_addr_7  ,2'h0}) ?   frontend__tlb__pmp__io_pmp_cfg_x_7  |  frontend__tlb__pmp__io_prv  [1]&~  frontend__tlb__pmp__io_pmp_cfg_l_7  :  frontend__tlb__pmp__io_prv  [1];
assign frontend__tlb__pmp__io_prv = 2'h3;
assign frontend__tlb__pmp__io_pmp_cfg_l_0 = frontend__tlb__io_ptw_pmp_cfg_l_0;
assign frontend__tlb__pmp__io_pmp_cfg_l_1 = frontend__tlb__io_ptw_pmp_cfg_l_1;
assign frontend__tlb__pmp__io_pmp_cfg_l_2 = frontend__tlb__io_ptw_pmp_cfg_l_2;
assign frontend__tlb__pmp__io_pmp_cfg_l_3 = frontend__tlb__io_ptw_pmp_cfg_l_3;
assign frontend__tlb__pmp__io_pmp_cfg_l_4 = frontend__tlb__io_ptw_pmp_cfg_l_4;
assign frontend__tlb__pmp__io_pmp_cfg_l_5 = frontend__tlb__io_ptw_pmp_cfg_l_5;
assign frontend__tlb__pmp__io_pmp_cfg_l_6 = frontend__tlb__io_ptw_pmp_cfg_l_6;
assign frontend__tlb__pmp__io_pmp_cfg_l_7 = frontend__tlb__io_ptw_pmp_cfg_l_7;
assign frontend__tlb__pmp__io_pmp_cfg_a_0 = frontend__tlb__io_ptw_pmp_cfg_a_0;
assign frontend__tlb__pmp__io_pmp_cfg_a_1 = frontend__tlb__io_ptw_pmp_cfg_a_1;
assign frontend__tlb__pmp__io_pmp_cfg_a_2 = frontend__tlb__io_ptw_pmp_cfg_a_2;
assign frontend__tlb__pmp__io_pmp_cfg_a_3 = frontend__tlb__io_ptw_pmp_cfg_a_3;
assign frontend__tlb__pmp__io_pmp_cfg_a_4 = frontend__tlb__io_ptw_pmp_cfg_a_4;
assign frontend__tlb__pmp__io_pmp_cfg_a_5 = frontend__tlb__io_ptw_pmp_cfg_a_5;
assign frontend__tlb__pmp__io_pmp_cfg_a_6 = frontend__tlb__io_ptw_pmp_cfg_a_6;
assign frontend__tlb__pmp__io_pmp_cfg_a_7 = frontend__tlb__io_ptw_pmp_cfg_a_7;
assign frontend__tlb__pmp__io_pmp_cfg_x_0 = frontend__tlb__io_ptw_pmp_cfg_x_0;
assign frontend__tlb__pmp__io_pmp_cfg_x_1 = frontend__tlb__io_ptw_pmp_cfg_x_1;
assign frontend__tlb__pmp__io_pmp_cfg_x_2 = frontend__tlb__io_ptw_pmp_cfg_x_2;
assign frontend__tlb__pmp__io_pmp_cfg_x_3 = frontend__tlb__io_ptw_pmp_cfg_x_3;
assign frontend__tlb__pmp__io_pmp_cfg_x_4 = frontend__tlb__io_ptw_pmp_cfg_x_4;
assign frontend__tlb__pmp__io_pmp_cfg_x_5 = frontend__tlb__io_ptw_pmp_cfg_x_5;
assign frontend__tlb__pmp__io_pmp_cfg_x_6 = frontend__tlb__io_ptw_pmp_cfg_x_6;
assign frontend__tlb__pmp__io_pmp_cfg_x_7 = frontend__tlb__io_ptw_pmp_cfg_x_7;
assign frontend__tlb__pmp__io_pmp_addr_0 = frontend__tlb__io_ptw_pmp_addr_0;
assign frontend__tlb__pmp__io_pmp_addr_1 = frontend__tlb__io_ptw_pmp_addr_1;
assign frontend__tlb__pmp__io_pmp_addr_2 = frontend__tlb__io_ptw_pmp_addr_2;
assign frontend__tlb__pmp__io_pmp_addr_3 = frontend__tlb__io_ptw_pmp_addr_3;
assign frontend__tlb__pmp__io_pmp_addr_4 = frontend__tlb__io_ptw_pmp_addr_4;
assign frontend__tlb__pmp__io_pmp_addr_5 = frontend__tlb__io_ptw_pmp_addr_5;
assign frontend__tlb__pmp__io_pmp_addr_6 = frontend__tlb__io_ptw_pmp_addr_6;
assign frontend__tlb__pmp__io_pmp_addr_7 = frontend__tlb__io_ptw_pmp_addr_7;
assign frontend__tlb__pmp__io_pmp_mask_0 = frontend__tlb__io_ptw_pmp_mask_0;
assign frontend__tlb__pmp__io_pmp_mask_1 = frontend__tlb__io_ptw_pmp_mask_1;
assign frontend__tlb__pmp__io_pmp_mask_2 = frontend__tlb__io_ptw_pmp_mask_2;
assign frontend__tlb__pmp__io_pmp_mask_3 = frontend__tlb__io_ptw_pmp_mask_3;
assign frontend__tlb__pmp__io_pmp_mask_4 = frontend__tlb__io_ptw_pmp_mask_4;
assign frontend__tlb__pmp__io_pmp_mask_5 = frontend__tlb__io_ptw_pmp_mask_5;
assign frontend__tlb__pmp__io_pmp_mask_6 = frontend__tlb__io_ptw_pmp_mask_6;
assign frontend__tlb__pmp__io_pmp_mask_7 = frontend__tlb__io_ptw_pmp_mask_7;
assign frontend__tlb__pmp__io_addr = frontend__tlb__io_req_bits_vaddr[31:0];
assign frontend__tlb___pmp_io_x = frontend__tlb__pmp__io_x;
  
  
wire  frontend__tlb__entries_barrier__io_x_u;
wire  frontend__tlb__entries_barrier__io_x_ae_ptw;
wire  frontend__tlb__entries_barrier__io_x_ae_final;
wire  frontend__tlb__entries_barrier__io_x_pf;
wire  frontend__tlb__entries_barrier__io_x_gf;
wire  frontend__tlb__entries_barrier__io_x_sw;
wire  frontend__tlb__entries_barrier__io_x_sx;
wire  frontend__tlb__entries_barrier__io_x_sr;
wire  frontend__tlb__entries_barrier__io_x_pw;
wire  frontend__tlb__entries_barrier__io_x_px;
wire  frontend__tlb__entries_barrier__io_x_pr;
wire  frontend__tlb__entries_barrier__io_x_ppp;
wire  frontend__tlb__entries_barrier__io_x_pal;
wire  frontend__tlb__entries_barrier__io_x_paa;
wire  frontend__tlb__entries_barrier__io_x_eff;
wire  frontend__tlb__entries_barrier__io_x_c;
wire  frontend__tlb__entries_barrier__io_y_u;
wire  frontend__tlb__entries_barrier__io_y_ae_ptw;
wire  frontend__tlb__entries_barrier__io_y_ae_final;
wire  frontend__tlb__entries_barrier__io_y_pf;
wire  frontend__tlb__entries_barrier__io_y_gf;
wire  frontend__tlb__entries_barrier__io_y_sw;
wire  frontend__tlb__entries_barrier__io_y_sx;
wire  frontend__tlb__entries_barrier__io_y_sr;
wire  frontend__tlb__entries_barrier__io_y_pw;
wire  frontend__tlb__entries_barrier__io_y_px;
wire  frontend__tlb__entries_barrier__io_y_pr;
wire  frontend__tlb__entries_barrier__io_y_ppp;
wire  frontend__tlb__entries_barrier__io_y_pal;
wire  frontend__tlb__entries_barrier__io_y_paa;
wire  frontend__tlb__entries_barrier__io_y_eff;
wire  frontend__tlb__entries_barrier__io_y_c;
wire  frontend__tlb__entries_barrier_1__io_x_u;
wire  frontend__tlb__entries_barrier_1__io_x_ae_ptw;
wire  frontend__tlb__entries_barrier_1__io_x_ae_final;
wire  frontend__tlb__entries_barrier_1__io_x_pf;
wire  frontend__tlb__entries_barrier_1__io_x_gf;
wire  frontend__tlb__entries_barrier_1__io_x_sw;
wire  frontend__tlb__entries_barrier_1__io_x_sx;
wire  frontend__tlb__entries_barrier_1__io_x_sr;
wire  frontend__tlb__entries_barrier_1__io_x_pw;
wire  frontend__tlb__entries_barrier_1__io_x_px;
wire  frontend__tlb__entries_barrier_1__io_x_pr;
wire  frontend__tlb__entries_barrier_1__io_x_ppp;
wire  frontend__tlb__entries_barrier_1__io_x_pal;
wire  frontend__tlb__entries_barrier_1__io_x_paa;
wire  frontend__tlb__entries_barrier_1__io_x_eff;
wire  frontend__tlb__entries_barrier_1__io_x_c;
wire  frontend__tlb__entries_barrier_1__io_y_u;
wire  frontend__tlb__entries_barrier_1__io_y_ae_ptw;
wire  frontend__tlb__entries_barrier_1__io_y_ae_final;
wire  frontend__tlb__entries_barrier_1__io_y_pf;
wire  frontend__tlb__entries_barrier_1__io_y_gf;
wire  frontend__tlb__entries_barrier_1__io_y_sw;
wire  frontend__tlb__entries_barrier_1__io_y_sx;
wire  frontend__tlb__entries_barrier_1__io_y_sr;
wire  frontend__tlb__entries_barrier_1__io_y_pw;
wire  frontend__tlb__entries_barrier_1__io_y_px;
wire  frontend__tlb__entries_barrier_1__io_y_pr;
wire  frontend__tlb__entries_barrier_1__io_y_ppp;
wire  frontend__tlb__entries_barrier_1__io_y_pal;
wire  frontend__tlb__entries_barrier_1__io_y_paa;
wire  frontend__tlb__entries_barrier_1__io_y_eff;
wire  frontend__tlb__entries_barrier_1__io_y_c;
wire  frontend__tlb__entries_barrier_2__io_x_u;
wire  frontend__tlb__entries_barrier_2__io_x_ae_ptw;
wire  frontend__tlb__entries_barrier_2__io_x_ae_final;
wire  frontend__tlb__entries_barrier_2__io_x_pf;
wire  frontend__tlb__entries_barrier_2__io_x_gf;
wire  frontend__tlb__entries_barrier_2__io_x_sw;
wire  frontend__tlb__entries_barrier_2__io_x_sx;
wire  frontend__tlb__entries_barrier_2__io_x_sr;
wire  frontend__tlb__entries_barrier_2__io_x_pw;
wire  frontend__tlb__entries_barrier_2__io_x_px;
wire  frontend__tlb__entries_barrier_2__io_x_pr;
wire  frontend__tlb__entries_barrier_2__io_x_ppp;
wire  frontend__tlb__entries_barrier_2__io_x_pal;
wire  frontend__tlb__entries_barrier_2__io_x_paa;
wire  frontend__tlb__entries_barrier_2__io_x_eff;
wire  frontend__tlb__entries_barrier_2__io_x_c;
wire  frontend__tlb__entries_barrier_2__io_y_u;
wire  frontend__tlb__entries_barrier_2__io_y_ae_ptw;
wire  frontend__tlb__entries_barrier_2__io_y_ae_final;
wire  frontend__tlb__entries_barrier_2__io_y_pf;
wire  frontend__tlb__entries_barrier_2__io_y_gf;
wire  frontend__tlb__entries_barrier_2__io_y_sw;
wire  frontend__tlb__entries_barrier_2__io_y_sx;
wire  frontend__tlb__entries_barrier_2__io_y_sr;
wire  frontend__tlb__entries_barrier_2__io_y_pw;
wire  frontend__tlb__entries_barrier_2__io_y_px;
wire  frontend__tlb__entries_barrier_2__io_y_pr;
wire  frontend__tlb__entries_barrier_2__io_y_ppp;
wire  frontend__tlb__entries_barrier_2__io_y_pal;
wire  frontend__tlb__entries_barrier_2__io_y_paa;
wire  frontend__tlb__entries_barrier_2__io_y_eff;
wire  frontend__tlb__entries_barrier_2__io_y_c;
wire  frontend__tlb__entries_barrier_3__io_x_u;
wire  frontend__tlb__entries_barrier_3__io_x_ae_ptw;
wire  frontend__tlb__entries_barrier_3__io_x_ae_final;
wire  frontend__tlb__entries_barrier_3__io_x_pf;
wire  frontend__tlb__entries_barrier_3__io_x_gf;
wire  frontend__tlb__entries_barrier_3__io_x_sw;
wire  frontend__tlb__entries_barrier_3__io_x_sx;
wire  frontend__tlb__entries_barrier_3__io_x_sr;
wire  frontend__tlb__entries_barrier_3__io_x_pw;
wire  frontend__tlb__entries_barrier_3__io_x_px;
wire  frontend__tlb__entries_barrier_3__io_x_pr;
wire  frontend__tlb__entries_barrier_3__io_x_ppp;
wire  frontend__tlb__entries_barrier_3__io_x_pal;
wire  frontend__tlb__entries_barrier_3__io_x_paa;
wire  frontend__tlb__entries_barrier_3__io_x_eff;
wire  frontend__tlb__entries_barrier_3__io_x_c;
wire  frontend__tlb__entries_barrier_3__io_y_u;
wire  frontend__tlb__entries_barrier_3__io_y_ae_ptw;
wire  frontend__tlb__entries_barrier_3__io_y_ae_final;
wire  frontend__tlb__entries_barrier_3__io_y_pf;
wire  frontend__tlb__entries_barrier_3__io_y_gf;
wire  frontend__tlb__entries_barrier_3__io_y_sw;
wire  frontend__tlb__entries_barrier_3__io_y_sx;
wire  frontend__tlb__entries_barrier_3__io_y_sr;
wire  frontend__tlb__entries_barrier_3__io_y_pw;
wire  frontend__tlb__entries_barrier_3__io_y_px;
wire  frontend__tlb__entries_barrier_3__io_y_pr;
wire  frontend__tlb__entries_barrier_3__io_y_ppp;
wire  frontend__tlb__entries_barrier_3__io_y_pal;
wire  frontend__tlb__entries_barrier_3__io_y_paa;
wire  frontend__tlb__entries_barrier_3__io_y_eff;
wire  frontend__tlb__entries_barrier_3__io_y_c;
wire  frontend__tlb__entries_barrier_4__io_x_u;
wire  frontend__tlb__entries_barrier_4__io_x_ae_ptw;
wire  frontend__tlb__entries_barrier_4__io_x_ae_final;
wire  frontend__tlb__entries_barrier_4__io_x_pf;
wire  frontend__tlb__entries_barrier_4__io_x_gf;
wire  frontend__tlb__entries_barrier_4__io_x_sw;
wire  frontend__tlb__entries_barrier_4__io_x_sx;
wire  frontend__tlb__entries_barrier_4__io_x_sr;
wire  frontend__tlb__entries_barrier_4__io_x_pw;
wire  frontend__tlb__entries_barrier_4__io_x_px;
wire  frontend__tlb__entries_barrier_4__io_x_pr;
wire  frontend__tlb__entries_barrier_4__io_x_ppp;
wire  frontend__tlb__entries_barrier_4__io_x_pal;
wire  frontend__tlb__entries_barrier_4__io_x_paa;
wire  frontend__tlb__entries_barrier_4__io_x_eff;
wire  frontend__tlb__entries_barrier_4__io_x_c;
wire  frontend__tlb__entries_barrier_4__io_y_u;
wire  frontend__tlb__entries_barrier_4__io_y_ae_ptw;
wire  frontend__tlb__entries_barrier_4__io_y_ae_final;
wire  frontend__tlb__entries_barrier_4__io_y_pf;
wire  frontend__tlb__entries_barrier_4__io_y_gf;
wire  frontend__tlb__entries_barrier_4__io_y_sw;
wire  frontend__tlb__entries_barrier_4__io_y_sx;
wire  frontend__tlb__entries_barrier_4__io_y_sr;
wire  frontend__tlb__entries_barrier_4__io_y_pw;
wire  frontend__tlb__entries_barrier_4__io_y_px;
wire  frontend__tlb__entries_barrier_4__io_y_pr;
wire  frontend__tlb__entries_barrier_4__io_y_ppp;
wire  frontend__tlb__entries_barrier_4__io_y_pal;
wire  frontend__tlb__entries_barrier_4__io_y_paa;
wire  frontend__tlb__entries_barrier_4__io_y_eff;
wire  frontend__tlb__entries_barrier_4__io_y_c;
wire  frontend__tlb__entries_barrier_5__io_x_u;
wire  frontend__tlb__entries_barrier_5__io_x_ae_ptw;
wire  frontend__tlb__entries_barrier_5__io_x_ae_final;
wire  frontend__tlb__entries_barrier_5__io_x_pf;
wire  frontend__tlb__entries_barrier_5__io_x_gf;
wire  frontend__tlb__entries_barrier_5__io_x_sw;
wire  frontend__tlb__entries_barrier_5__io_x_sx;
wire  frontend__tlb__entries_barrier_5__io_x_sr;
wire  frontend__tlb__entries_barrier_5__io_x_pw;
wire  frontend__tlb__entries_barrier_5__io_x_px;
wire  frontend__tlb__entries_barrier_5__io_x_pr;
wire  frontend__tlb__entries_barrier_5__io_x_ppp;
wire  frontend__tlb__entries_barrier_5__io_x_pal;
wire  frontend__tlb__entries_barrier_5__io_x_paa;
wire  frontend__tlb__entries_barrier_5__io_x_eff;
wire  frontend__tlb__entries_barrier_5__io_x_c;
wire  frontend__tlb__entries_barrier_5__io_y_u;
wire  frontend__tlb__entries_barrier_5__io_y_ae_ptw;
wire  frontend__tlb__entries_barrier_5__io_y_ae_final;
wire  frontend__tlb__entries_barrier_5__io_y_pf;
wire  frontend__tlb__entries_barrier_5__io_y_gf;
wire  frontend__tlb__entries_barrier_5__io_y_sw;
wire  frontend__tlb__entries_barrier_5__io_y_sx;
wire  frontend__tlb__entries_barrier_5__io_y_sr;
wire  frontend__tlb__entries_barrier_5__io_y_pw;
wire  frontend__tlb__entries_barrier_5__io_y_px;
wire  frontend__tlb__entries_barrier_5__io_y_pr;
wire  frontend__tlb__entries_barrier_5__io_y_ppp;
wire  frontend__tlb__entries_barrier_5__io_y_pal;
wire  frontend__tlb__entries_barrier_5__io_y_paa;
wire  frontend__tlb__entries_barrier_5__io_y_eff;
wire  frontend__tlb__entries_barrier_5__io_y_c;
 
  assign   frontend__tlb__entries_barrier__io_y_u  =  frontend__tlb__entries_barrier__io_x_u  ; 
  assign   frontend__tlb__entries_barrier__io_y_ae_ptw  =  frontend__tlb__entries_barrier__io_x_ae_ptw  ; 
  assign   frontend__tlb__entries_barrier__io_y_ae_final  =  frontend__tlb__entries_barrier__io_x_ae_final  ; 
  assign   frontend__tlb__entries_barrier__io_y_pf  =  frontend__tlb__entries_barrier__io_x_pf  ; 
  assign   frontend__tlb__entries_barrier__io_y_gf  =  frontend__tlb__entries_barrier__io_x_gf  ; 
  assign   frontend__tlb__entries_barrier__io_y_sw  =  frontend__tlb__entries_barrier__io_x_sw  ; 
  assign   frontend__tlb__entries_barrier__io_y_sx  =  frontend__tlb__entries_barrier__io_x_sx  ; 
  assign   frontend__tlb__entries_barrier__io_y_sr  =  frontend__tlb__entries_barrier__io_x_sr  ; 
  assign   frontend__tlb__entries_barrier__io_y_pw  =  frontend__tlb__entries_barrier__io_x_pw  ; 
  assign   frontend__tlb__entries_barrier__io_y_px  =  frontend__tlb__entries_barrier__io_x_px  ; 
  assign   frontend__tlb__entries_barrier__io_y_pr  =  frontend__tlb__entries_barrier__io_x_pr  ; 
  assign   frontend__tlb__entries_barrier__io_y_ppp  =  frontend__tlb__entries_barrier__io_x_ppp  ; 
  assign   frontend__tlb__entries_barrier__io_y_pal  =  frontend__tlb__entries_barrier__io_x_pal  ; 
  assign   frontend__tlb__entries_barrier__io_y_paa  =  frontend__tlb__entries_barrier__io_x_paa  ; 
  assign   frontend__tlb__entries_barrier__io_y_eff  =  frontend__tlb__entries_barrier__io_x_eff  ; 
  assign   frontend__tlb__entries_barrier__io_y_c  =  frontend__tlb__entries_barrier__io_x_c  ;
  
  
 
  assign   frontend__tlb__entries_barrier_1__io_y_u  =  frontend__tlb__entries_barrier_1__io_x_u  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_ae_ptw  =  frontend__tlb__entries_barrier_1__io_x_ae_ptw  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_ae_final  =  frontend__tlb__entries_barrier_1__io_x_ae_final  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_pf  =  frontend__tlb__entries_barrier_1__io_x_pf  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_gf  =  frontend__tlb__entries_barrier_1__io_x_gf  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_sw  =  frontend__tlb__entries_barrier_1__io_x_sw  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_sx  =  frontend__tlb__entries_barrier_1__io_x_sx  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_sr  =  frontend__tlb__entries_barrier_1__io_x_sr  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_pw  =  frontend__tlb__entries_barrier_1__io_x_pw  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_px  =  frontend__tlb__entries_barrier_1__io_x_px  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_pr  =  frontend__tlb__entries_barrier_1__io_x_pr  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_ppp  =  frontend__tlb__entries_barrier_1__io_x_ppp  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_pal  =  frontend__tlb__entries_barrier_1__io_x_pal  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_paa  =  frontend__tlb__entries_barrier_1__io_x_paa  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_eff  =  frontend__tlb__entries_barrier_1__io_x_eff  ; 
  assign   frontend__tlb__entries_barrier_1__io_y_c  =  frontend__tlb__entries_barrier_1__io_x_c  ;
  
  
 
  assign   frontend__tlb__entries_barrier_2__io_y_u  =  frontend__tlb__entries_barrier_2__io_x_u  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_ae_ptw  =  frontend__tlb__entries_barrier_2__io_x_ae_ptw  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_ae_final  =  frontend__tlb__entries_barrier_2__io_x_ae_final  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_pf  =  frontend__tlb__entries_barrier_2__io_x_pf  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_gf  =  frontend__tlb__entries_barrier_2__io_x_gf  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_sw  =  frontend__tlb__entries_barrier_2__io_x_sw  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_sx  =  frontend__tlb__entries_barrier_2__io_x_sx  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_sr  =  frontend__tlb__entries_barrier_2__io_x_sr  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_pw  =  frontend__tlb__entries_barrier_2__io_x_pw  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_px  =  frontend__tlb__entries_barrier_2__io_x_px  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_pr  =  frontend__tlb__entries_barrier_2__io_x_pr  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_ppp  =  frontend__tlb__entries_barrier_2__io_x_ppp  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_pal  =  frontend__tlb__entries_barrier_2__io_x_pal  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_paa  =  frontend__tlb__entries_barrier_2__io_x_paa  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_eff  =  frontend__tlb__entries_barrier_2__io_x_eff  ; 
  assign   frontend__tlb__entries_barrier_2__io_y_c  =  frontend__tlb__entries_barrier_2__io_x_c  ;
  
  
 
  assign   frontend__tlb__entries_barrier_3__io_y_u  =  frontend__tlb__entries_barrier_3__io_x_u  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_ae_ptw  =  frontend__tlb__entries_barrier_3__io_x_ae_ptw  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_ae_final  =  frontend__tlb__entries_barrier_3__io_x_ae_final  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_pf  =  frontend__tlb__entries_barrier_3__io_x_pf  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_gf  =  frontend__tlb__entries_barrier_3__io_x_gf  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_sw  =  frontend__tlb__entries_barrier_3__io_x_sw  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_sx  =  frontend__tlb__entries_barrier_3__io_x_sx  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_sr  =  frontend__tlb__entries_barrier_3__io_x_sr  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_pw  =  frontend__tlb__entries_barrier_3__io_x_pw  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_px  =  frontend__tlb__entries_barrier_3__io_x_px  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_pr  =  frontend__tlb__entries_barrier_3__io_x_pr  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_ppp  =  frontend__tlb__entries_barrier_3__io_x_ppp  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_pal  =  frontend__tlb__entries_barrier_3__io_x_pal  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_paa  =  frontend__tlb__entries_barrier_3__io_x_paa  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_eff  =  frontend__tlb__entries_barrier_3__io_x_eff  ; 
  assign   frontend__tlb__entries_barrier_3__io_y_c  =  frontend__tlb__entries_barrier_3__io_x_c  ;
  
  
 
  assign   frontend__tlb__entries_barrier_4__io_y_u  =  frontend__tlb__entries_barrier_4__io_x_u  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_ae_ptw  =  frontend__tlb__entries_barrier_4__io_x_ae_ptw  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_ae_final  =  frontend__tlb__entries_barrier_4__io_x_ae_final  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_pf  =  frontend__tlb__entries_barrier_4__io_x_pf  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_gf  =  frontend__tlb__entries_barrier_4__io_x_gf  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_sw  =  frontend__tlb__entries_barrier_4__io_x_sw  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_sx  =  frontend__tlb__entries_barrier_4__io_x_sx  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_sr  =  frontend__tlb__entries_barrier_4__io_x_sr  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_pw  =  frontend__tlb__entries_barrier_4__io_x_pw  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_px  =  frontend__tlb__entries_barrier_4__io_x_px  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_pr  =  frontend__tlb__entries_barrier_4__io_x_pr  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_ppp  =  frontend__tlb__entries_barrier_4__io_x_ppp  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_pal  =  frontend__tlb__entries_barrier_4__io_x_pal  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_paa  =  frontend__tlb__entries_barrier_4__io_x_paa  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_eff  =  frontend__tlb__entries_barrier_4__io_x_eff  ; 
  assign   frontend__tlb__entries_barrier_4__io_y_c  =  frontend__tlb__entries_barrier_4__io_x_c  ;
  
  
 
  assign   frontend__tlb__entries_barrier_5__io_y_u  =  frontend__tlb__entries_barrier_5__io_x_u  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_ae_ptw  =  frontend__tlb__entries_barrier_5__io_x_ae_ptw  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_ae_final  =  frontend__tlb__entries_barrier_5__io_x_ae_final  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_pf  =  frontend__tlb__entries_barrier_5__io_x_pf  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_gf  =  frontend__tlb__entries_barrier_5__io_x_gf  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_sw  =  frontend__tlb__entries_barrier_5__io_x_sw  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_sx  =  frontend__tlb__entries_barrier_5__io_x_sx  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_sr  =  frontend__tlb__entries_barrier_5__io_x_sr  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_pw  =  frontend__tlb__entries_barrier_5__io_x_pw  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_px  =  frontend__tlb__entries_barrier_5__io_x_px  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_pr  =  frontend__tlb__entries_barrier_5__io_x_pr  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_ppp  =  frontend__tlb__entries_barrier_5__io_x_ppp  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_pal  =  frontend__tlb__entries_barrier_5__io_x_pal  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_paa  =  frontend__tlb__entries_barrier_5__io_x_paa  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_eff  =  frontend__tlb__entries_barrier_5__io_x_eff  ; 
  assign   frontend__tlb__entries_barrier_5__io_y_c  =  frontend__tlb__entries_barrier_5__io_x_c  ;
assign frontend__tlb__entries_barrier__io_x_u = 1'h0;
assign frontend__tlb__entries_barrier__io_x_ae_ptw = 1'h0;
assign frontend__tlb__entries_barrier__io_x_ae_final = 1'h0;
assign frontend__tlb__entries_barrier__io_x_pf = 1'h0;
assign frontend__tlb__entries_barrier__io_x_gf = 1'h0;
assign frontend__tlb__entries_barrier__io_x_sw = 1'h0;
assign frontend__tlb__entries_barrier__io_x_sx = 1'h0;
assign frontend__tlb__entries_barrier__io_x_sr = 1'h0;
assign frontend__tlb__entries_barrier__io_x_pw = 1'h0;
assign frontend__tlb__entries_barrier__io_x_px = 1'h0;
assign frontend__tlb__entries_barrier__io_x_pr = 1'h0;
assign frontend__tlb__entries_barrier__io_x_ppp = 1'h0;
assign frontend__tlb__entries_barrier__io_x_pal = 1'h0;
assign frontend__tlb__entries_barrier__io_x_paa = 1'h0;
assign frontend__tlb__entries_barrier__io_x_eff = 1'h0;
assign frontend__tlb__entries_barrier__io_x_c = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_u = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_ae_ptw = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_ae_final = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_pf = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_gf = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_sw = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_sx = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_sr = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_pw = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_px = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_pr = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_ppp = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_pal = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_paa = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_eff = 1'h0;
assign frontend__tlb__entries_barrier_1__io_x_c = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_u = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_ae_ptw = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_ae_final = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_pf = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_gf = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_sw = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_sx = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_sr = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_pw = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_px = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_pr = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_ppp = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_pal = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_paa = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_eff = 1'h0;
assign frontend__tlb__entries_barrier_2__io_x_c = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_u = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_ae_ptw = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_ae_final = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_pf = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_gf = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_sw = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_sx = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_sr = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_pw = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_px = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_pr = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_ppp = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_pal = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_paa = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_eff = 1'h0;
assign frontend__tlb__entries_barrier_3__io_x_c = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_u = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_ae_ptw = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_ae_final = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_pf = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_gf = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_sw = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_sx = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_sr = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_pw = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_px = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_pr = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_ppp = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_pal = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_paa = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_eff = 1'h0;
assign frontend__tlb__entries_barrier_4__io_x_c = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_u = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_ae_ptw = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_ae_final = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_pf = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_gf = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_sw = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_sx = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_sr = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_pw = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_px = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_pr = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_ppp = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_pal = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_paa = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_eff = 1'h0;
assign frontend__tlb__entries_barrier_5__io_x_c = 1'h0;
 
  assign   frontend__tlb__io_resp_paddr  =  frontend__tlb__io_req_bits_vaddr  [31:0]; 
  assign   frontend__tlb__io_resp_pf_inst  =1'h0; 
  assign   frontend__tlb__io_resp_ae_inst  =~(  frontend__tlb__legal_address  &({  frontend__tlb__io_req_bits_vaddr  [31:30],  frontend__tlb__io_req_bits_vaddr  [27],  frontend__tlb__io_req_bits_vaddr  [25]}==4'h0|{  frontend__tlb__io_req_bits_vaddr  [31],~(  frontend__tlb__io_req_bits_vaddr  [30])}==2'h0|  frontend__tlb___GEN  [3:2]==2'h0)&~(~  frontend__tlb__io_ptw_status_debug  &~(|(  frontend__tlb__io_req_bits_vaddr  [33:12])))&  frontend__tlb___pmp_io_x  ); 
  assign   frontend__tlb__io_resp_cacheable  =  frontend__tlb__legal_address  &~(  frontend__tlb___GEN  [3]); 
  assign   frontend__tlb__io_ptw_req_bits_bits_need_gpa  =1'h0; 
  assign   frontend__tlb__io_ptw_req_bits_bits_stage2  =1'h0;
assign frontend__tlb__io_req_bits_vaddr = frontend__s1_pc;
assign frontend___tlb_io_resp_paddr = frontend__tlb__io_resp_paddr;
assign frontend___tlb_io_resp_pf_inst = frontend__tlb__io_resp_pf_inst;
assign frontend___tlb_io_resp_ae_inst = frontend__tlb__io_resp_ae_inst;
assign frontend___tlb_io_resp_cacheable = frontend__tlb__io_resp_cacheable;
assign frontend__io_ptw_req_bits_bits_need_gpa = frontend__tlb__io_ptw_req_bits_bits_need_gpa;
assign frontend__io_ptw_req_bits_bits_stage2 = frontend__tlb__io_ptw_req_bits_bits_stage2;
assign frontend__tlb__io_ptw_status_debug = frontend__io_ptw_status_debug;
assign frontend__tlb__io_ptw_pmp_cfg_l_0 = frontend__io_ptw_pmp_cfg_l_0;
assign frontend__tlb__io_ptw_pmp_cfg_l_1 = frontend__io_ptw_pmp_cfg_l_1;
assign frontend__tlb__io_ptw_pmp_cfg_l_2 = frontend__io_ptw_pmp_cfg_l_2;
assign frontend__tlb__io_ptw_pmp_cfg_l_3 = frontend__io_ptw_pmp_cfg_l_3;
assign frontend__tlb__io_ptw_pmp_cfg_l_4 = frontend__io_ptw_pmp_cfg_l_4;
assign frontend__tlb__io_ptw_pmp_cfg_l_5 = frontend__io_ptw_pmp_cfg_l_5;
assign frontend__tlb__io_ptw_pmp_cfg_l_6 = frontend__io_ptw_pmp_cfg_l_6;
assign frontend__tlb__io_ptw_pmp_cfg_l_7 = frontend__io_ptw_pmp_cfg_l_7;
assign frontend__tlb__io_ptw_pmp_cfg_a_0 = frontend__io_ptw_pmp_cfg_a_0;
assign frontend__tlb__io_ptw_pmp_cfg_a_1 = frontend__io_ptw_pmp_cfg_a_1;
assign frontend__tlb__io_ptw_pmp_cfg_a_2 = frontend__io_ptw_pmp_cfg_a_2;
assign frontend__tlb__io_ptw_pmp_cfg_a_3 = frontend__io_ptw_pmp_cfg_a_3;
assign frontend__tlb__io_ptw_pmp_cfg_a_4 = frontend__io_ptw_pmp_cfg_a_4;
assign frontend__tlb__io_ptw_pmp_cfg_a_5 = frontend__io_ptw_pmp_cfg_a_5;
assign frontend__tlb__io_ptw_pmp_cfg_a_6 = frontend__io_ptw_pmp_cfg_a_6;
assign frontend__tlb__io_ptw_pmp_cfg_a_7 = frontend__io_ptw_pmp_cfg_a_7;
assign frontend__tlb__io_ptw_pmp_cfg_x_0 = frontend__io_ptw_pmp_cfg_x_0;
assign frontend__tlb__io_ptw_pmp_cfg_x_1 = frontend__io_ptw_pmp_cfg_x_1;
assign frontend__tlb__io_ptw_pmp_cfg_x_2 = frontend__io_ptw_pmp_cfg_x_2;
assign frontend__tlb__io_ptw_pmp_cfg_x_3 = frontend__io_ptw_pmp_cfg_x_3;
assign frontend__tlb__io_ptw_pmp_cfg_x_4 = frontend__io_ptw_pmp_cfg_x_4;
assign frontend__tlb__io_ptw_pmp_cfg_x_5 = frontend__io_ptw_pmp_cfg_x_5;
assign frontend__tlb__io_ptw_pmp_cfg_x_6 = frontend__io_ptw_pmp_cfg_x_6;
assign frontend__tlb__io_ptw_pmp_cfg_x_7 = frontend__io_ptw_pmp_cfg_x_7;
assign frontend__tlb__io_ptw_pmp_addr_0 = frontend__io_ptw_pmp_addr_0;
assign frontend__tlb__io_ptw_pmp_addr_1 = frontend__io_ptw_pmp_addr_1;
assign frontend__tlb__io_ptw_pmp_addr_2 = frontend__io_ptw_pmp_addr_2;
assign frontend__tlb__io_ptw_pmp_addr_3 = frontend__io_ptw_pmp_addr_3;
assign frontend__tlb__io_ptw_pmp_addr_4 = frontend__io_ptw_pmp_addr_4;
assign frontend__tlb__io_ptw_pmp_addr_5 = frontend__io_ptw_pmp_addr_5;
assign frontend__tlb__io_ptw_pmp_addr_6 = frontend__io_ptw_pmp_addr_6;
assign frontend__tlb__io_ptw_pmp_addr_7 = frontend__io_ptw_pmp_addr_7;
assign frontend__tlb__io_ptw_pmp_mask_0 = frontend__io_ptw_pmp_mask_0;
assign frontend__tlb__io_ptw_pmp_mask_1 = frontend__io_ptw_pmp_mask_1;
assign frontend__tlb__io_ptw_pmp_mask_2 = frontend__io_ptw_pmp_mask_2;
assign frontend__tlb__io_ptw_pmp_mask_3 = frontend__io_ptw_pmp_mask_3;
assign frontend__tlb__io_ptw_pmp_mask_4 = frontend__io_ptw_pmp_mask_4;
assign frontend__tlb__io_ptw_pmp_mask_5 = frontend__io_ptw_pmp_mask_5;
assign frontend__tlb__io_ptw_pmp_mask_6 = frontend__io_ptw_pmp_mask_6;
assign frontend__tlb__io_ptw_pmp_mask_7 = frontend__io_ptw_pmp_mask_7;

assign frontend__clock = clock;
assign frontend__reset = reset;
assign frontend__auto_icache_master_out_a_ready = _tlMasterXbar_auto_in_1_a_ready;
assign _frontend_auto_icache_master_out_a_valid = frontend__auto_icache_master_out_a_valid;
assign _frontend_auto_icache_master_out_a_bits_address = frontend__auto_icache_master_out_a_bits_address;
assign frontend__auto_icache_master_out_d_valid = _tlMasterXbar_auto_in_1_d_valid;
assign frontend__auto_icache_master_out_d_bits_opcode = _tlMasterXbar_auto_in_1_d_bits_opcode;
assign frontend__auto_icache_master_out_d_bits_size = _tlMasterXbar_auto_in_1_d_bits_size;
assign frontend__auto_icache_master_out_d_bits_data = _tlMasterXbar_auto_in_1_d_bits_data;
assign frontend__auto_icache_master_out_d_bits_corrupt = _tlMasterXbar_auto_in_1_d_bits_corrupt;
assign frontend__io_cpu_might_request = _core_io_imem_might_request;
assign frontend__io_cpu_req_valid = _core_io_imem_req_valid;
assign frontend__io_cpu_req_bits_pc = _core_io_imem_req_bits_pc;
assign frontend__io_cpu_req_bits_speculative = _core_io_imem_req_bits_speculative;
assign frontend__io_cpu_resp_ready = _core_io_imem_resp_ready;
assign _frontend_io_cpu_resp_valid = frontend__io_cpu_resp_valid;
assign _frontend_io_cpu_resp_bits_pc = frontend__io_cpu_resp_bits_pc;
assign _frontend_io_cpu_resp_bits_data = frontend__io_cpu_resp_bits_data;
assign _frontend_io_cpu_resp_bits_xcpt_pf_inst = frontend__io_cpu_resp_bits_xcpt_pf_inst;
assign _frontend_io_cpu_resp_bits_xcpt_gf_inst = frontend__io_cpu_resp_bits_xcpt_gf_inst;
assign _frontend_io_cpu_resp_bits_xcpt_ae_inst = frontend__io_cpu_resp_bits_xcpt_ae_inst;
assign _frontend_io_cpu_resp_bits_replay = frontend__io_cpu_resp_bits_replay;
assign frontend__io_cpu_btb_update_valid = _core_io_imem_btb_update_valid;
assign frontend__io_cpu_bht_update_valid = _core_io_imem_bht_update_valid;
assign frontend__io_cpu_flush_icache = _core_io_imem_flush_icache;
assign _frontend_io_ptw_req_bits_bits_need_gpa = frontend__io_ptw_req_bits_bits_need_gpa;
assign _frontend_io_ptw_req_bits_bits_stage2 = frontend__io_ptw_req_bits_bits_stage2;
assign frontend__io_ptw_status_debug = _ptw_io_requestor_1_status_debug;
assign frontend__io_ptw_pmp_cfg_l_0 = _ptw_io_requestor_1_pmp_cfg_l_0;
assign frontend__io_ptw_pmp_cfg_l_1 = _ptw_io_requestor_1_pmp_cfg_l_1;
assign frontend__io_ptw_pmp_cfg_l_2 = _ptw_io_requestor_1_pmp_cfg_l_2;
assign frontend__io_ptw_pmp_cfg_l_3 = _ptw_io_requestor_1_pmp_cfg_l_3;
assign frontend__io_ptw_pmp_cfg_l_4 = _ptw_io_requestor_1_pmp_cfg_l_4;
assign frontend__io_ptw_pmp_cfg_l_5 = _ptw_io_requestor_1_pmp_cfg_l_5;
assign frontend__io_ptw_pmp_cfg_l_6 = _ptw_io_requestor_1_pmp_cfg_l_6;
assign frontend__io_ptw_pmp_cfg_l_7 = _ptw_io_requestor_1_pmp_cfg_l_7;
assign frontend__io_ptw_pmp_cfg_a_0 = _ptw_io_requestor_1_pmp_cfg_a_0;
assign frontend__io_ptw_pmp_cfg_a_1 = _ptw_io_requestor_1_pmp_cfg_a_1;
assign frontend__io_ptw_pmp_cfg_a_2 = _ptw_io_requestor_1_pmp_cfg_a_2;
assign frontend__io_ptw_pmp_cfg_a_3 = _ptw_io_requestor_1_pmp_cfg_a_3;
assign frontend__io_ptw_pmp_cfg_a_4 = _ptw_io_requestor_1_pmp_cfg_a_4;
assign frontend__io_ptw_pmp_cfg_a_5 = _ptw_io_requestor_1_pmp_cfg_a_5;
assign frontend__io_ptw_pmp_cfg_a_6 = _ptw_io_requestor_1_pmp_cfg_a_6;
assign frontend__io_ptw_pmp_cfg_a_7 = _ptw_io_requestor_1_pmp_cfg_a_7;
assign frontend__io_ptw_pmp_cfg_x_0 = _ptw_io_requestor_1_pmp_cfg_x_0;
assign frontend__io_ptw_pmp_cfg_x_1 = _ptw_io_requestor_1_pmp_cfg_x_1;
assign frontend__io_ptw_pmp_cfg_x_2 = _ptw_io_requestor_1_pmp_cfg_x_2;
assign frontend__io_ptw_pmp_cfg_x_3 = _ptw_io_requestor_1_pmp_cfg_x_3;
assign frontend__io_ptw_pmp_cfg_x_4 = _ptw_io_requestor_1_pmp_cfg_x_4;
assign frontend__io_ptw_pmp_cfg_x_5 = _ptw_io_requestor_1_pmp_cfg_x_5;
assign frontend__io_ptw_pmp_cfg_x_6 = _ptw_io_requestor_1_pmp_cfg_x_6;
assign frontend__io_ptw_pmp_cfg_x_7 = _ptw_io_requestor_1_pmp_cfg_x_7;
assign frontend__io_ptw_pmp_addr_0 = _ptw_io_requestor_1_pmp_addr_0;
assign frontend__io_ptw_pmp_addr_1 = _ptw_io_requestor_1_pmp_addr_1;
assign frontend__io_ptw_pmp_addr_2 = _ptw_io_requestor_1_pmp_addr_2;
assign frontend__io_ptw_pmp_addr_3 = _ptw_io_requestor_1_pmp_addr_3;
assign frontend__io_ptw_pmp_addr_4 = _ptw_io_requestor_1_pmp_addr_4;
assign frontend__io_ptw_pmp_addr_5 = _ptw_io_requestor_1_pmp_addr_5;
assign frontend__io_ptw_pmp_addr_6 = _ptw_io_requestor_1_pmp_addr_6;
assign frontend__io_ptw_pmp_addr_7 = _ptw_io_requestor_1_pmp_addr_7;
assign frontend__io_ptw_pmp_mask_0 = _ptw_io_requestor_1_pmp_mask_0;
assign frontend__io_ptw_pmp_mask_1 = _ptw_io_requestor_1_pmp_mask_1;
assign frontend__io_ptw_pmp_mask_2 = _ptw_io_requestor_1_pmp_mask_2;
assign frontend__io_ptw_pmp_mask_3 = _ptw_io_requestor_1_pmp_mask_3;
assign frontend__io_ptw_pmp_mask_4 = _ptw_io_requestor_1_pmp_mask_4;
assign frontend__io_ptw_pmp_mask_5 = _ptw_io_requestor_1_pmp_mask_5;
assign frontend__io_ptw_pmp_mask_6 = _ptw_io_requestor_1_pmp_mask_6;
assign frontend__io_ptw_pmp_mask_7 = _ptw_io_requestor_1_pmp_mask_7;
assign frontend__io_ptw_customCSRs_csrs_0_value = _ptw_io_requestor_1_customCSRs_csrs_0_value;
 
  
wire  dcacheArb__io_requestor_0_req_ready;
wire  dcacheArb__io_requestor_0_req_valid;
wire [33:0] dcacheArb__io_requestor_0_req_bits_addr;
wire [5:0] dcacheArb__io_requestor_0_req_bits_tag;
wire [4:0] dcacheArb__io_requestor_0_req_bits_cmd;
wire [1:0] dcacheArb__io_requestor_0_req_bits_size;
wire  dcacheArb__io_requestor_0_req_bits_signed;
wire  dcacheArb__io_requestor_0_req_bits_dv;
wire  dcacheArb__io_requestor_0_s1_kill;
wire [63:0] dcacheArb__io_requestor_0_s1_data_data;
wire  dcacheArb__io_requestor_0_s2_nack;
wire  dcacheArb__io_requestor_0_resp_valid;
wire [5:0] dcacheArb__io_requestor_0_resp_bits_tag;
wire [63:0] dcacheArb__io_requestor_0_resp_bits_data;
wire  dcacheArb__io_requestor_0_resp_bits_replay;
wire  dcacheArb__io_requestor_0_resp_bits_has_data;
wire [63:0] dcacheArb__io_requestor_0_resp_bits_data_word_bypass;
wire  dcacheArb__io_requestor_0_replay_next;
wire  dcacheArb__io_requestor_0_s2_xcpt_ma_ld;
wire  dcacheArb__io_requestor_0_s2_xcpt_ma_st;
wire  dcacheArb__io_requestor_0_s2_xcpt_pf_ld;
wire  dcacheArb__io_requestor_0_s2_xcpt_pf_st;
wire  dcacheArb__io_requestor_0_s2_xcpt_ae_ld;
wire  dcacheArb__io_requestor_0_s2_xcpt_ae_st;
wire  dcacheArb__io_requestor_0_ordered;
wire  dcacheArb__io_requestor_0_perf_release;
wire  dcacheArb__io_requestor_0_perf_grant;
wire  dcacheArb__io_mem_req_ready;
wire  dcacheArb__io_mem_req_valid;
wire [33:0] dcacheArb__io_mem_req_bits_addr;
wire [5:0] dcacheArb__io_mem_req_bits_tag;
wire [4:0] dcacheArb__io_mem_req_bits_cmd;
wire [1:0] dcacheArb__io_mem_req_bits_size;
wire  dcacheArb__io_mem_req_bits_signed;
wire  dcacheArb__io_mem_req_bits_dv;
wire  dcacheArb__io_mem_s1_kill;
wire [63:0] dcacheArb__io_mem_s1_data_data;
wire  dcacheArb__io_mem_s2_nack;
wire  dcacheArb__io_mem_resp_valid;
wire [5:0] dcacheArb__io_mem_resp_bits_tag;
wire [63:0] dcacheArb__io_mem_resp_bits_data;
wire  dcacheArb__io_mem_resp_bits_replay;
wire  dcacheArb__io_mem_resp_bits_has_data;
wire [63:0] dcacheArb__io_mem_resp_bits_data_word_bypass;
wire  dcacheArb__io_mem_replay_next;
wire  dcacheArb__io_mem_s2_xcpt_ma_ld;
wire  dcacheArb__io_mem_s2_xcpt_ma_st;
wire  dcacheArb__io_mem_s2_xcpt_pf_ld;
wire  dcacheArb__io_mem_s2_xcpt_pf_st;
wire  dcacheArb__io_mem_s2_xcpt_ae_ld;
wire  dcacheArb__io_mem_s2_xcpt_ae_st;
wire  dcacheArb__io_mem_ordered;
wire  dcacheArb__io_mem_perf_release;
wire  dcacheArb__io_mem_perf_grant;
 
  assign   dcacheArb__io_requestor_0_req_ready  =  dcacheArb__io_mem_req_ready  ; 
  assign   dcacheArb__io_requestor_0_s2_nack  =  dcacheArb__io_mem_s2_nack  ; 
  assign   dcacheArb__io_requestor_0_resp_valid  =  dcacheArb__io_mem_resp_valid  ; 
  assign   dcacheArb__io_requestor_0_resp_bits_tag  =  dcacheArb__io_mem_resp_bits_tag  ; 
  assign   dcacheArb__io_requestor_0_resp_bits_data  =  dcacheArb__io_mem_resp_bits_data  ; 
  assign   dcacheArb__io_requestor_0_resp_bits_replay  =  dcacheArb__io_mem_resp_bits_replay  ; 
  assign   dcacheArb__io_requestor_0_resp_bits_has_data  =  dcacheArb__io_mem_resp_bits_has_data  ; 
  assign   dcacheArb__io_requestor_0_resp_bits_data_word_bypass  =  dcacheArb__io_mem_resp_bits_data_word_bypass  ; 
  assign   dcacheArb__io_requestor_0_replay_next  =  dcacheArb__io_mem_replay_next  ; 
  assign   dcacheArb__io_requestor_0_s2_xcpt_ma_ld  =  dcacheArb__io_mem_s2_xcpt_ma_ld  ; 
  assign   dcacheArb__io_requestor_0_s2_xcpt_ma_st  =  dcacheArb__io_mem_s2_xcpt_ma_st  ; 
  assign   dcacheArb__io_requestor_0_s2_xcpt_pf_ld  =  dcacheArb__io_mem_s2_xcpt_pf_ld  ; 
  assign   dcacheArb__io_requestor_0_s2_xcpt_pf_st  =  dcacheArb__io_mem_s2_xcpt_pf_st  ; 
  assign   dcacheArb__io_requestor_0_s2_xcpt_ae_ld  =  dcacheArb__io_mem_s2_xcpt_ae_ld  ; 
  assign   dcacheArb__io_requestor_0_s2_xcpt_ae_st  =  dcacheArb__io_mem_s2_xcpt_ae_st  ; 
  assign   dcacheArb__io_requestor_0_ordered  =  dcacheArb__io_mem_ordered  ; 
  assign   dcacheArb__io_requestor_0_perf_release  =  dcacheArb__io_mem_perf_release  ; 
  assign   dcacheArb__io_requestor_0_perf_grant  =  dcacheArb__io_mem_perf_grant  ; 
  assign   dcacheArb__io_mem_req_valid  =  dcacheArb__io_requestor_0_req_valid  ; 
  assign   dcacheArb__io_mem_req_bits_addr  =  dcacheArb__io_requestor_0_req_bits_addr  ; 
  assign   dcacheArb__io_mem_req_bits_tag  =  dcacheArb__io_requestor_0_req_bits_tag  ; 
  assign   dcacheArb__io_mem_req_bits_cmd  =  dcacheArb__io_requestor_0_req_bits_cmd  ; 
  assign   dcacheArb__io_mem_req_bits_size  =  dcacheArb__io_requestor_0_req_bits_size  ; 
  assign   dcacheArb__io_mem_req_bits_signed  =  dcacheArb__io_requestor_0_req_bits_signed  ; 
  assign   dcacheArb__io_mem_req_bits_dv  =  dcacheArb__io_requestor_0_req_bits_dv  ; 
  assign   dcacheArb__io_mem_s1_kill  =  dcacheArb__io_requestor_0_s1_kill  ; 
  assign   dcacheArb__io_mem_s1_data_data  =  dcacheArb__io_requestor_0_s1_data_data  ;
assign _dcacheArb_io_requestor_0_req_ready = dcacheArb__io_requestor_0_req_ready;
assign dcacheArb__io_requestor_0_req_valid = _core_io_dmem_req_valid;
assign dcacheArb__io_requestor_0_req_bits_addr = _core_io_dmem_req_bits_addr;
assign dcacheArb__io_requestor_0_req_bits_tag = _core_io_dmem_req_bits_tag;
assign dcacheArb__io_requestor_0_req_bits_cmd = _core_io_dmem_req_bits_cmd;
assign dcacheArb__io_requestor_0_req_bits_size = _core_io_dmem_req_bits_size;
assign dcacheArb__io_requestor_0_req_bits_signed = _core_io_dmem_req_bits_signed;
assign dcacheArb__io_requestor_0_req_bits_dv = _core_io_dmem_req_bits_dv;
assign dcacheArb__io_requestor_0_s1_kill = _core_io_dmem_s1_kill;
assign dcacheArb__io_requestor_0_s1_data_data = _core_io_dmem_s1_data_data;
assign _dcacheArb_io_requestor_0_s2_nack = dcacheArb__io_requestor_0_s2_nack;
assign _dcacheArb_io_requestor_0_resp_valid = dcacheArb__io_requestor_0_resp_valid;
assign _dcacheArb_io_requestor_0_resp_bits_tag = dcacheArb__io_requestor_0_resp_bits_tag;
assign _dcacheArb_io_requestor_0_resp_bits_data = dcacheArb__io_requestor_0_resp_bits_data;
assign _dcacheArb_io_requestor_0_resp_bits_replay = dcacheArb__io_requestor_0_resp_bits_replay;
assign _dcacheArb_io_requestor_0_resp_bits_has_data = dcacheArb__io_requestor_0_resp_bits_has_data;
assign _dcacheArb_io_requestor_0_resp_bits_data_word_bypass = dcacheArb__io_requestor_0_resp_bits_data_word_bypass;
assign _dcacheArb_io_requestor_0_replay_next = dcacheArb__io_requestor_0_replay_next;
assign _dcacheArb_io_requestor_0_s2_xcpt_ma_ld = dcacheArb__io_requestor_0_s2_xcpt_ma_ld;
assign _dcacheArb_io_requestor_0_s2_xcpt_ma_st = dcacheArb__io_requestor_0_s2_xcpt_ma_st;
assign _dcacheArb_io_requestor_0_s2_xcpt_pf_ld = dcacheArb__io_requestor_0_s2_xcpt_pf_ld;
assign _dcacheArb_io_requestor_0_s2_xcpt_pf_st = dcacheArb__io_requestor_0_s2_xcpt_pf_st;
assign _dcacheArb_io_requestor_0_s2_xcpt_ae_ld = dcacheArb__io_requestor_0_s2_xcpt_ae_ld;
assign _dcacheArb_io_requestor_0_s2_xcpt_ae_st = dcacheArb__io_requestor_0_s2_xcpt_ae_st;
assign _dcacheArb_io_requestor_0_ordered = dcacheArb__io_requestor_0_ordered;
assign _dcacheArb_io_requestor_0_perf_release = dcacheArb__io_requestor_0_perf_release;
assign _dcacheArb_io_requestor_0_perf_grant = dcacheArb__io_requestor_0_perf_grant;
assign dcacheArb__io_mem_req_ready = _dcache_io_cpu_req_ready;
assign _dcacheArb_io_mem_req_valid = dcacheArb__io_mem_req_valid;
assign _dcacheArb_io_mem_req_bits_addr = dcacheArb__io_mem_req_bits_addr;
assign _dcacheArb_io_mem_req_bits_tag = dcacheArb__io_mem_req_bits_tag;
assign _dcacheArb_io_mem_req_bits_cmd = dcacheArb__io_mem_req_bits_cmd;
assign _dcacheArb_io_mem_req_bits_size = dcacheArb__io_mem_req_bits_size;
assign _dcacheArb_io_mem_req_bits_signed = dcacheArb__io_mem_req_bits_signed;
assign _dcacheArb_io_mem_req_bits_dv = dcacheArb__io_mem_req_bits_dv;
assign _dcacheArb_io_mem_s1_kill = dcacheArb__io_mem_s1_kill;
assign _dcacheArb_io_mem_s1_data_data = dcacheArb__io_mem_s1_data_data;
assign dcacheArb__io_mem_s2_nack = _dcache_io_cpu_s2_nack;
assign dcacheArb__io_mem_resp_valid = _dcache_io_cpu_resp_valid;
assign dcacheArb__io_mem_resp_bits_tag = _dcache_io_cpu_resp_bits_tag;
assign dcacheArb__io_mem_resp_bits_data = _dcache_io_cpu_resp_bits_data;
assign dcacheArb__io_mem_resp_bits_replay = _dcache_io_cpu_resp_bits_replay;
assign dcacheArb__io_mem_resp_bits_has_data = _dcache_io_cpu_resp_bits_has_data;
assign dcacheArb__io_mem_resp_bits_data_word_bypass = _dcache_io_cpu_resp_bits_data_word_bypass;
assign dcacheArb__io_mem_replay_next = _dcache_io_cpu_replay_next;
assign dcacheArb__io_mem_s2_xcpt_ma_ld = _dcache_io_cpu_s2_xcpt_ma_ld;
assign dcacheArb__io_mem_s2_xcpt_ma_st = _dcache_io_cpu_s2_xcpt_ma_st;
assign dcacheArb__io_mem_s2_xcpt_pf_ld = _dcache_io_cpu_s2_xcpt_pf_ld;
assign dcacheArb__io_mem_s2_xcpt_pf_st = _dcache_io_cpu_s2_xcpt_pf_st;
assign dcacheArb__io_mem_s2_xcpt_ae_ld = _dcache_io_cpu_s2_xcpt_ae_ld;
assign dcacheArb__io_mem_s2_xcpt_ae_st = _dcache_io_cpu_s2_xcpt_ae_st;
assign dcacheArb__io_mem_ordered = _dcache_io_cpu_ordered;
assign dcacheArb__io_mem_perf_release = _dcache_io_cpu_perf_release;
assign dcacheArb__io_mem_perf_grant = _dcache_io_cpu_perf_grant;
 
  
wire  ptw__clock;
wire  ptw__io_requestor_0_req_bits_bits_need_gpa;
wire  ptw__io_requestor_0_req_bits_bits_stage2;
wire  ptw__io_requestor_0_status_debug;
wire  ptw__io_requestor_0_pmp_cfg_l_0;
wire  ptw__io_requestor_0_pmp_cfg_l_1;
wire  ptw__io_requestor_0_pmp_cfg_l_2;
wire  ptw__io_requestor_0_pmp_cfg_l_3;
wire  ptw__io_requestor_0_pmp_cfg_l_4;
wire  ptw__io_requestor_0_pmp_cfg_l_5;
wire  ptw__io_requestor_0_pmp_cfg_l_6;
wire  ptw__io_requestor_0_pmp_cfg_l_7;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_0;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_1;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_2;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_3;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_4;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_5;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_6;
wire [1:0] ptw__io_requestor_0_pmp_cfg_a_7;
wire  ptw__io_requestor_0_pmp_cfg_w_0;
wire  ptw__io_requestor_0_pmp_cfg_w_1;
wire  ptw__io_requestor_0_pmp_cfg_w_2;
wire  ptw__io_requestor_0_pmp_cfg_w_3;
wire  ptw__io_requestor_0_pmp_cfg_w_4;
wire  ptw__io_requestor_0_pmp_cfg_w_5;
wire  ptw__io_requestor_0_pmp_cfg_w_6;
wire  ptw__io_requestor_0_pmp_cfg_w_7;
wire  ptw__io_requestor_0_pmp_cfg_r_0;
wire  ptw__io_requestor_0_pmp_cfg_r_1;
wire  ptw__io_requestor_0_pmp_cfg_r_2;
wire  ptw__io_requestor_0_pmp_cfg_r_3;
wire  ptw__io_requestor_0_pmp_cfg_r_4;
wire  ptw__io_requestor_0_pmp_cfg_r_5;
wire  ptw__io_requestor_0_pmp_cfg_r_6;
wire  ptw__io_requestor_0_pmp_cfg_r_7;
wire [29:0] ptw__io_requestor_0_pmp_addr_0;
wire [29:0] ptw__io_requestor_0_pmp_addr_1;
wire [29:0] ptw__io_requestor_0_pmp_addr_2;
wire [29:0] ptw__io_requestor_0_pmp_addr_3;
wire [29:0] ptw__io_requestor_0_pmp_addr_4;
wire [29:0] ptw__io_requestor_0_pmp_addr_5;
wire [29:0] ptw__io_requestor_0_pmp_addr_6;
wire [29:0] ptw__io_requestor_0_pmp_addr_7;
wire [31:0] ptw__io_requestor_0_pmp_mask_0;
wire [31:0] ptw__io_requestor_0_pmp_mask_1;
wire [31:0] ptw__io_requestor_0_pmp_mask_2;
wire [31:0] ptw__io_requestor_0_pmp_mask_3;
wire [31:0] ptw__io_requestor_0_pmp_mask_4;
wire [31:0] ptw__io_requestor_0_pmp_mask_5;
wire [31:0] ptw__io_requestor_0_pmp_mask_6;
wire [31:0] ptw__io_requestor_0_pmp_mask_7;
wire  ptw__io_requestor_1_req_bits_bits_need_gpa;
wire  ptw__io_requestor_1_req_bits_bits_stage2;
wire  ptw__io_requestor_1_status_debug;
wire  ptw__io_requestor_1_pmp_cfg_l_0;
wire  ptw__io_requestor_1_pmp_cfg_l_1;
wire  ptw__io_requestor_1_pmp_cfg_l_2;
wire  ptw__io_requestor_1_pmp_cfg_l_3;
wire  ptw__io_requestor_1_pmp_cfg_l_4;
wire  ptw__io_requestor_1_pmp_cfg_l_5;
wire  ptw__io_requestor_1_pmp_cfg_l_6;
wire  ptw__io_requestor_1_pmp_cfg_l_7;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_0;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_1;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_2;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_3;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_4;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_5;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_6;
wire [1:0] ptw__io_requestor_1_pmp_cfg_a_7;
wire  ptw__io_requestor_1_pmp_cfg_x_0;
wire  ptw__io_requestor_1_pmp_cfg_x_1;
wire  ptw__io_requestor_1_pmp_cfg_x_2;
wire  ptw__io_requestor_1_pmp_cfg_x_3;
wire  ptw__io_requestor_1_pmp_cfg_x_4;
wire  ptw__io_requestor_1_pmp_cfg_x_5;
wire  ptw__io_requestor_1_pmp_cfg_x_6;
wire  ptw__io_requestor_1_pmp_cfg_x_7;
wire [29:0] ptw__io_requestor_1_pmp_addr_0;
wire [29:0] ptw__io_requestor_1_pmp_addr_1;
wire [29:0] ptw__io_requestor_1_pmp_addr_2;
wire [29:0] ptw__io_requestor_1_pmp_addr_3;
wire [29:0] ptw__io_requestor_1_pmp_addr_4;
wire [29:0] ptw__io_requestor_1_pmp_addr_5;
wire [29:0] ptw__io_requestor_1_pmp_addr_6;
wire [29:0] ptw__io_requestor_1_pmp_addr_7;
wire [31:0] ptw__io_requestor_1_pmp_mask_0;
wire [31:0] ptw__io_requestor_1_pmp_mask_1;
wire [31:0] ptw__io_requestor_1_pmp_mask_2;
wire [31:0] ptw__io_requestor_1_pmp_mask_3;
wire [31:0] ptw__io_requestor_1_pmp_mask_4;
wire [31:0] ptw__io_requestor_1_pmp_mask_5;
wire [31:0] ptw__io_requestor_1_pmp_mask_6;
wire [31:0] ptw__io_requestor_1_pmp_mask_7;
wire [63:0] ptw__io_requestor_1_customCSRs_csrs_0_value;
wire  ptw__io_dpath_status_debug;
wire  ptw__io_dpath_pmp_cfg_l_0;
wire  ptw__io_dpath_pmp_cfg_l_1;
wire  ptw__io_dpath_pmp_cfg_l_2;
wire  ptw__io_dpath_pmp_cfg_l_3;
wire  ptw__io_dpath_pmp_cfg_l_4;
wire  ptw__io_dpath_pmp_cfg_l_5;
wire  ptw__io_dpath_pmp_cfg_l_6;
wire  ptw__io_dpath_pmp_cfg_l_7;
wire [1:0] ptw__io_dpath_pmp_cfg_a_0;
wire [1:0] ptw__io_dpath_pmp_cfg_a_1;
wire [1:0] ptw__io_dpath_pmp_cfg_a_2;
wire [1:0] ptw__io_dpath_pmp_cfg_a_3;
wire [1:0] ptw__io_dpath_pmp_cfg_a_4;
wire [1:0] ptw__io_dpath_pmp_cfg_a_5;
wire [1:0] ptw__io_dpath_pmp_cfg_a_6;
wire [1:0] ptw__io_dpath_pmp_cfg_a_7;
wire  ptw__io_dpath_pmp_cfg_x_0;
wire  ptw__io_dpath_pmp_cfg_x_1;
wire  ptw__io_dpath_pmp_cfg_x_2;
wire  ptw__io_dpath_pmp_cfg_x_3;
wire  ptw__io_dpath_pmp_cfg_x_4;
wire  ptw__io_dpath_pmp_cfg_x_5;
wire  ptw__io_dpath_pmp_cfg_x_6;
wire  ptw__io_dpath_pmp_cfg_x_7;
wire  ptw__io_dpath_pmp_cfg_w_0;
wire  ptw__io_dpath_pmp_cfg_w_1;
wire  ptw__io_dpath_pmp_cfg_w_2;
wire  ptw__io_dpath_pmp_cfg_w_3;
wire  ptw__io_dpath_pmp_cfg_w_4;
wire  ptw__io_dpath_pmp_cfg_w_5;
wire  ptw__io_dpath_pmp_cfg_w_6;
wire  ptw__io_dpath_pmp_cfg_w_7;
wire  ptw__io_dpath_pmp_cfg_r_0;
wire  ptw__io_dpath_pmp_cfg_r_1;
wire  ptw__io_dpath_pmp_cfg_r_2;
wire  ptw__io_dpath_pmp_cfg_r_3;
wire  ptw__io_dpath_pmp_cfg_r_4;
wire  ptw__io_dpath_pmp_cfg_r_5;
wire  ptw__io_dpath_pmp_cfg_r_6;
wire  ptw__io_dpath_pmp_cfg_r_7;
wire [29:0] ptw__io_dpath_pmp_addr_0;
wire [29:0] ptw__io_dpath_pmp_addr_1;
wire [29:0] ptw__io_dpath_pmp_addr_2;
wire [29:0] ptw__io_dpath_pmp_addr_3;
wire [29:0] ptw__io_dpath_pmp_addr_4;
wire [29:0] ptw__io_dpath_pmp_addr_5;
wire [29:0] ptw__io_dpath_pmp_addr_6;
wire [29:0] ptw__io_dpath_pmp_addr_7;
wire [31:0] ptw__io_dpath_pmp_mask_0;
wire [31:0] ptw__io_dpath_pmp_mask_1;
wire [31:0] ptw__io_dpath_pmp_mask_2;
wire [31:0] ptw__io_dpath_pmp_mask_3;
wire [31:0] ptw__io_dpath_pmp_mask_4;
wire [31:0] ptw__io_dpath_pmp_mask_5;
wire [31:0] ptw__io_dpath_pmp_mask_6;
wire [31:0] ptw__io_dpath_pmp_mask_7;
wire [63:0] ptw__io_dpath_customCSRs_csrs_0_value;
  
  
wire  ptw__arb__io_in_0_bits_bits_need_gpa;
wire  ptw__arb__io_in_0_bits_bits_stage2;
wire  ptw__arb__io_in_1_bits_bits_need_gpa;
wire  ptw__arb__io_in_1_bits_bits_stage2;
wire  ptw__arb__io_out_bits_bits_need_gpa;
wire  ptw__arb__io_out_bits_bits_stage2;
 
  assign   ptw__arb__io_out_bits_bits_need_gpa  =  ptw__arb__io_in_1_bits_bits_need_gpa  ; 
  assign   ptw__arb__io_out_bits_bits_stage2  =  ptw__arb__io_in_1_bits_bits_stage2  ;
assign ptw__arb__io_in_0_bits_bits_need_gpa = ptw__io_requestor_0_req_bits_bits_need_gpa;
assign ptw__arb__io_in_0_bits_bits_stage2 = ptw__io_requestor_0_req_bits_bits_stage2;
assign ptw__arb__io_in_1_bits_bits_need_gpa = ptw__io_requestor_1_req_bits_bits_need_gpa;
assign ptw__arb__io_in_1_bits_bits_stage2 = ptw__io_requestor_1_req_bits_bits_stage2;
 
  assign   ptw__io_requestor_0_status_debug  =  ptw__io_dpath_status_debug  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_0  =  ptw__io_dpath_pmp_cfg_l_0  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_1  =  ptw__io_dpath_pmp_cfg_l_1  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_2  =  ptw__io_dpath_pmp_cfg_l_2  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_3  =  ptw__io_dpath_pmp_cfg_l_3  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_4  =  ptw__io_dpath_pmp_cfg_l_4  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_5  =  ptw__io_dpath_pmp_cfg_l_5  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_6  =  ptw__io_dpath_pmp_cfg_l_6  ; 
  assign   ptw__io_requestor_0_pmp_cfg_l_7  =  ptw__io_dpath_pmp_cfg_l_7  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_0  =  ptw__io_dpath_pmp_cfg_a_0  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_1  =  ptw__io_dpath_pmp_cfg_a_1  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_2  =  ptw__io_dpath_pmp_cfg_a_2  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_3  =  ptw__io_dpath_pmp_cfg_a_3  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_4  =  ptw__io_dpath_pmp_cfg_a_4  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_5  =  ptw__io_dpath_pmp_cfg_a_5  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_6  =  ptw__io_dpath_pmp_cfg_a_6  ; 
  assign   ptw__io_requestor_0_pmp_cfg_a_7  =  ptw__io_dpath_pmp_cfg_a_7  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_0  =  ptw__io_dpath_pmp_cfg_w_0  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_1  =  ptw__io_dpath_pmp_cfg_w_1  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_2  =  ptw__io_dpath_pmp_cfg_w_2  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_3  =  ptw__io_dpath_pmp_cfg_w_3  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_4  =  ptw__io_dpath_pmp_cfg_w_4  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_5  =  ptw__io_dpath_pmp_cfg_w_5  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_6  =  ptw__io_dpath_pmp_cfg_w_6  ; 
  assign   ptw__io_requestor_0_pmp_cfg_w_7  =  ptw__io_dpath_pmp_cfg_w_7  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_0  =  ptw__io_dpath_pmp_cfg_r_0  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_1  =  ptw__io_dpath_pmp_cfg_r_1  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_2  =  ptw__io_dpath_pmp_cfg_r_2  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_3  =  ptw__io_dpath_pmp_cfg_r_3  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_4  =  ptw__io_dpath_pmp_cfg_r_4  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_5  =  ptw__io_dpath_pmp_cfg_r_5  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_6  =  ptw__io_dpath_pmp_cfg_r_6  ; 
  assign   ptw__io_requestor_0_pmp_cfg_r_7  =  ptw__io_dpath_pmp_cfg_r_7  ; 
  assign   ptw__io_requestor_0_pmp_addr_0  =  ptw__io_dpath_pmp_addr_0  ; 
  assign   ptw__io_requestor_0_pmp_addr_1  =  ptw__io_dpath_pmp_addr_1  ; 
  assign   ptw__io_requestor_0_pmp_addr_2  =  ptw__io_dpath_pmp_addr_2  ; 
  assign   ptw__io_requestor_0_pmp_addr_3  =  ptw__io_dpath_pmp_addr_3  ; 
  assign   ptw__io_requestor_0_pmp_addr_4  =  ptw__io_dpath_pmp_addr_4  ; 
  assign   ptw__io_requestor_0_pmp_addr_5  =  ptw__io_dpath_pmp_addr_5  ; 
  assign   ptw__io_requestor_0_pmp_addr_6  =  ptw__io_dpath_pmp_addr_6  ; 
  assign   ptw__io_requestor_0_pmp_addr_7  =  ptw__io_dpath_pmp_addr_7  ; 
  assign   ptw__io_requestor_0_pmp_mask_0  =  ptw__io_dpath_pmp_mask_0  ; 
  assign   ptw__io_requestor_0_pmp_mask_1  =  ptw__io_dpath_pmp_mask_1  ; 
  assign   ptw__io_requestor_0_pmp_mask_2  =  ptw__io_dpath_pmp_mask_2  ; 
  assign   ptw__io_requestor_0_pmp_mask_3  =  ptw__io_dpath_pmp_mask_3  ; 
  assign   ptw__io_requestor_0_pmp_mask_4  =  ptw__io_dpath_pmp_mask_4  ; 
  assign   ptw__io_requestor_0_pmp_mask_5  =  ptw__io_dpath_pmp_mask_5  ; 
  assign   ptw__io_requestor_0_pmp_mask_6  =  ptw__io_dpath_pmp_mask_6  ; 
  assign   ptw__io_requestor_0_pmp_mask_7  =  ptw__io_dpath_pmp_mask_7  ; 
  assign   ptw__io_requestor_1_status_debug  =  ptw__io_dpath_status_debug  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_0  =  ptw__io_dpath_pmp_cfg_l_0  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_1  =  ptw__io_dpath_pmp_cfg_l_1  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_2  =  ptw__io_dpath_pmp_cfg_l_2  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_3  =  ptw__io_dpath_pmp_cfg_l_3  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_4  =  ptw__io_dpath_pmp_cfg_l_4  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_5  =  ptw__io_dpath_pmp_cfg_l_5  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_6  =  ptw__io_dpath_pmp_cfg_l_6  ; 
  assign   ptw__io_requestor_1_pmp_cfg_l_7  =  ptw__io_dpath_pmp_cfg_l_7  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_0  =  ptw__io_dpath_pmp_cfg_a_0  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_1  =  ptw__io_dpath_pmp_cfg_a_1  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_2  =  ptw__io_dpath_pmp_cfg_a_2  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_3  =  ptw__io_dpath_pmp_cfg_a_3  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_4  =  ptw__io_dpath_pmp_cfg_a_4  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_5  =  ptw__io_dpath_pmp_cfg_a_5  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_6  =  ptw__io_dpath_pmp_cfg_a_6  ; 
  assign   ptw__io_requestor_1_pmp_cfg_a_7  =  ptw__io_dpath_pmp_cfg_a_7  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_0  =  ptw__io_dpath_pmp_cfg_x_0  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_1  =  ptw__io_dpath_pmp_cfg_x_1  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_2  =  ptw__io_dpath_pmp_cfg_x_2  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_3  =  ptw__io_dpath_pmp_cfg_x_3  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_4  =  ptw__io_dpath_pmp_cfg_x_4  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_5  =  ptw__io_dpath_pmp_cfg_x_5  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_6  =  ptw__io_dpath_pmp_cfg_x_6  ; 
  assign   ptw__io_requestor_1_pmp_cfg_x_7  =  ptw__io_dpath_pmp_cfg_x_7  ; 
  assign   ptw__io_requestor_1_pmp_addr_0  =  ptw__io_dpath_pmp_addr_0  ; 
  assign   ptw__io_requestor_1_pmp_addr_1  =  ptw__io_dpath_pmp_addr_1  ; 
  assign   ptw__io_requestor_1_pmp_addr_2  =  ptw__io_dpath_pmp_addr_2  ; 
  assign   ptw__io_requestor_1_pmp_addr_3  =  ptw__io_dpath_pmp_addr_3  ; 
  assign   ptw__io_requestor_1_pmp_addr_4  =  ptw__io_dpath_pmp_addr_4  ; 
  assign   ptw__io_requestor_1_pmp_addr_5  =  ptw__io_dpath_pmp_addr_5  ; 
  assign   ptw__io_requestor_1_pmp_addr_6  =  ptw__io_dpath_pmp_addr_6  ; 
  assign   ptw__io_requestor_1_pmp_addr_7  =  ptw__io_dpath_pmp_addr_7  ; 
  assign   ptw__io_requestor_1_pmp_mask_0  =  ptw__io_dpath_pmp_mask_0  ; 
  assign   ptw__io_requestor_1_pmp_mask_1  =  ptw__io_dpath_pmp_mask_1  ; 
  assign   ptw__io_requestor_1_pmp_mask_2  =  ptw__io_dpath_pmp_mask_2  ; 
  assign   ptw__io_requestor_1_pmp_mask_3  =  ptw__io_dpath_pmp_mask_3  ; 
  assign   ptw__io_requestor_1_pmp_mask_4  =  ptw__io_dpath_pmp_mask_4  ; 
  assign   ptw__io_requestor_1_pmp_mask_5  =  ptw__io_dpath_pmp_mask_5  ; 
  assign   ptw__io_requestor_1_pmp_mask_6  =  ptw__io_dpath_pmp_mask_6  ; 
  assign   ptw__io_requestor_1_pmp_mask_7  =  ptw__io_dpath_pmp_mask_7  ; 
  assign   ptw__io_requestor_1_customCSRs_csrs_0_value  =  ptw__io_dpath_customCSRs_csrs_0_value  ;
assign ptw__clock = clock;
assign ptw__io_requestor_0_req_bits_bits_need_gpa = _dcache_io_ptw_req_bits_bits_need_gpa;
assign ptw__io_requestor_0_req_bits_bits_stage2 = _dcache_io_ptw_req_bits_bits_stage2;
assign _ptw_io_requestor_0_status_debug = ptw__io_requestor_0_status_debug;
assign _ptw_io_requestor_0_pmp_cfg_l_0 = ptw__io_requestor_0_pmp_cfg_l_0;
assign _ptw_io_requestor_0_pmp_cfg_l_1 = ptw__io_requestor_0_pmp_cfg_l_1;
assign _ptw_io_requestor_0_pmp_cfg_l_2 = ptw__io_requestor_0_pmp_cfg_l_2;
assign _ptw_io_requestor_0_pmp_cfg_l_3 = ptw__io_requestor_0_pmp_cfg_l_3;
assign _ptw_io_requestor_0_pmp_cfg_l_4 = ptw__io_requestor_0_pmp_cfg_l_4;
assign _ptw_io_requestor_0_pmp_cfg_l_5 = ptw__io_requestor_0_pmp_cfg_l_5;
assign _ptw_io_requestor_0_pmp_cfg_l_6 = ptw__io_requestor_0_pmp_cfg_l_6;
assign _ptw_io_requestor_0_pmp_cfg_l_7 = ptw__io_requestor_0_pmp_cfg_l_7;
assign _ptw_io_requestor_0_pmp_cfg_a_0 = ptw__io_requestor_0_pmp_cfg_a_0;
assign _ptw_io_requestor_0_pmp_cfg_a_1 = ptw__io_requestor_0_pmp_cfg_a_1;
assign _ptw_io_requestor_0_pmp_cfg_a_2 = ptw__io_requestor_0_pmp_cfg_a_2;
assign _ptw_io_requestor_0_pmp_cfg_a_3 = ptw__io_requestor_0_pmp_cfg_a_3;
assign _ptw_io_requestor_0_pmp_cfg_a_4 = ptw__io_requestor_0_pmp_cfg_a_4;
assign _ptw_io_requestor_0_pmp_cfg_a_5 = ptw__io_requestor_0_pmp_cfg_a_5;
assign _ptw_io_requestor_0_pmp_cfg_a_6 = ptw__io_requestor_0_pmp_cfg_a_6;
assign _ptw_io_requestor_0_pmp_cfg_a_7 = ptw__io_requestor_0_pmp_cfg_a_7;
assign _ptw_io_requestor_0_pmp_cfg_w_0 = ptw__io_requestor_0_pmp_cfg_w_0;
assign _ptw_io_requestor_0_pmp_cfg_w_1 = ptw__io_requestor_0_pmp_cfg_w_1;
assign _ptw_io_requestor_0_pmp_cfg_w_2 = ptw__io_requestor_0_pmp_cfg_w_2;
assign _ptw_io_requestor_0_pmp_cfg_w_3 = ptw__io_requestor_0_pmp_cfg_w_3;
assign _ptw_io_requestor_0_pmp_cfg_w_4 = ptw__io_requestor_0_pmp_cfg_w_4;
assign _ptw_io_requestor_0_pmp_cfg_w_5 = ptw__io_requestor_0_pmp_cfg_w_5;
assign _ptw_io_requestor_0_pmp_cfg_w_6 = ptw__io_requestor_0_pmp_cfg_w_6;
assign _ptw_io_requestor_0_pmp_cfg_w_7 = ptw__io_requestor_0_pmp_cfg_w_7;
assign _ptw_io_requestor_0_pmp_cfg_r_0 = ptw__io_requestor_0_pmp_cfg_r_0;
assign _ptw_io_requestor_0_pmp_cfg_r_1 = ptw__io_requestor_0_pmp_cfg_r_1;
assign _ptw_io_requestor_0_pmp_cfg_r_2 = ptw__io_requestor_0_pmp_cfg_r_2;
assign _ptw_io_requestor_0_pmp_cfg_r_3 = ptw__io_requestor_0_pmp_cfg_r_3;
assign _ptw_io_requestor_0_pmp_cfg_r_4 = ptw__io_requestor_0_pmp_cfg_r_4;
assign _ptw_io_requestor_0_pmp_cfg_r_5 = ptw__io_requestor_0_pmp_cfg_r_5;
assign _ptw_io_requestor_0_pmp_cfg_r_6 = ptw__io_requestor_0_pmp_cfg_r_6;
assign _ptw_io_requestor_0_pmp_cfg_r_7 = ptw__io_requestor_0_pmp_cfg_r_7;
assign _ptw_io_requestor_0_pmp_addr_0 = ptw__io_requestor_0_pmp_addr_0;
assign _ptw_io_requestor_0_pmp_addr_1 = ptw__io_requestor_0_pmp_addr_1;
assign _ptw_io_requestor_0_pmp_addr_2 = ptw__io_requestor_0_pmp_addr_2;
assign _ptw_io_requestor_0_pmp_addr_3 = ptw__io_requestor_0_pmp_addr_3;
assign _ptw_io_requestor_0_pmp_addr_4 = ptw__io_requestor_0_pmp_addr_4;
assign _ptw_io_requestor_0_pmp_addr_5 = ptw__io_requestor_0_pmp_addr_5;
assign _ptw_io_requestor_0_pmp_addr_6 = ptw__io_requestor_0_pmp_addr_6;
assign _ptw_io_requestor_0_pmp_addr_7 = ptw__io_requestor_0_pmp_addr_7;
assign _ptw_io_requestor_0_pmp_mask_0 = ptw__io_requestor_0_pmp_mask_0;
assign _ptw_io_requestor_0_pmp_mask_1 = ptw__io_requestor_0_pmp_mask_1;
assign _ptw_io_requestor_0_pmp_mask_2 = ptw__io_requestor_0_pmp_mask_2;
assign _ptw_io_requestor_0_pmp_mask_3 = ptw__io_requestor_0_pmp_mask_3;
assign _ptw_io_requestor_0_pmp_mask_4 = ptw__io_requestor_0_pmp_mask_4;
assign _ptw_io_requestor_0_pmp_mask_5 = ptw__io_requestor_0_pmp_mask_5;
assign _ptw_io_requestor_0_pmp_mask_6 = ptw__io_requestor_0_pmp_mask_6;
assign _ptw_io_requestor_0_pmp_mask_7 = ptw__io_requestor_0_pmp_mask_7;
assign ptw__io_requestor_1_req_bits_bits_need_gpa = _frontend_io_ptw_req_bits_bits_need_gpa;
assign ptw__io_requestor_1_req_bits_bits_stage2 = _frontend_io_ptw_req_bits_bits_stage2;
assign _ptw_io_requestor_1_status_debug = ptw__io_requestor_1_status_debug;
assign _ptw_io_requestor_1_pmp_cfg_l_0 = ptw__io_requestor_1_pmp_cfg_l_0;
assign _ptw_io_requestor_1_pmp_cfg_l_1 = ptw__io_requestor_1_pmp_cfg_l_1;
assign _ptw_io_requestor_1_pmp_cfg_l_2 = ptw__io_requestor_1_pmp_cfg_l_2;
assign _ptw_io_requestor_1_pmp_cfg_l_3 = ptw__io_requestor_1_pmp_cfg_l_3;
assign _ptw_io_requestor_1_pmp_cfg_l_4 = ptw__io_requestor_1_pmp_cfg_l_4;
assign _ptw_io_requestor_1_pmp_cfg_l_5 = ptw__io_requestor_1_pmp_cfg_l_5;
assign _ptw_io_requestor_1_pmp_cfg_l_6 = ptw__io_requestor_1_pmp_cfg_l_6;
assign _ptw_io_requestor_1_pmp_cfg_l_7 = ptw__io_requestor_1_pmp_cfg_l_7;
assign _ptw_io_requestor_1_pmp_cfg_a_0 = ptw__io_requestor_1_pmp_cfg_a_0;
assign _ptw_io_requestor_1_pmp_cfg_a_1 = ptw__io_requestor_1_pmp_cfg_a_1;
assign _ptw_io_requestor_1_pmp_cfg_a_2 = ptw__io_requestor_1_pmp_cfg_a_2;
assign _ptw_io_requestor_1_pmp_cfg_a_3 = ptw__io_requestor_1_pmp_cfg_a_3;
assign _ptw_io_requestor_1_pmp_cfg_a_4 = ptw__io_requestor_1_pmp_cfg_a_4;
assign _ptw_io_requestor_1_pmp_cfg_a_5 = ptw__io_requestor_1_pmp_cfg_a_5;
assign _ptw_io_requestor_1_pmp_cfg_a_6 = ptw__io_requestor_1_pmp_cfg_a_6;
assign _ptw_io_requestor_1_pmp_cfg_a_7 = ptw__io_requestor_1_pmp_cfg_a_7;
assign _ptw_io_requestor_1_pmp_cfg_x_0 = ptw__io_requestor_1_pmp_cfg_x_0;
assign _ptw_io_requestor_1_pmp_cfg_x_1 = ptw__io_requestor_1_pmp_cfg_x_1;
assign _ptw_io_requestor_1_pmp_cfg_x_2 = ptw__io_requestor_1_pmp_cfg_x_2;
assign _ptw_io_requestor_1_pmp_cfg_x_3 = ptw__io_requestor_1_pmp_cfg_x_3;
assign _ptw_io_requestor_1_pmp_cfg_x_4 = ptw__io_requestor_1_pmp_cfg_x_4;
assign _ptw_io_requestor_1_pmp_cfg_x_5 = ptw__io_requestor_1_pmp_cfg_x_5;
assign _ptw_io_requestor_1_pmp_cfg_x_6 = ptw__io_requestor_1_pmp_cfg_x_6;
assign _ptw_io_requestor_1_pmp_cfg_x_7 = ptw__io_requestor_1_pmp_cfg_x_7;
assign _ptw_io_requestor_1_pmp_addr_0 = ptw__io_requestor_1_pmp_addr_0;
assign _ptw_io_requestor_1_pmp_addr_1 = ptw__io_requestor_1_pmp_addr_1;
assign _ptw_io_requestor_1_pmp_addr_2 = ptw__io_requestor_1_pmp_addr_2;
assign _ptw_io_requestor_1_pmp_addr_3 = ptw__io_requestor_1_pmp_addr_3;
assign _ptw_io_requestor_1_pmp_addr_4 = ptw__io_requestor_1_pmp_addr_4;
assign _ptw_io_requestor_1_pmp_addr_5 = ptw__io_requestor_1_pmp_addr_5;
assign _ptw_io_requestor_1_pmp_addr_6 = ptw__io_requestor_1_pmp_addr_6;
assign _ptw_io_requestor_1_pmp_addr_7 = ptw__io_requestor_1_pmp_addr_7;
assign _ptw_io_requestor_1_pmp_mask_0 = ptw__io_requestor_1_pmp_mask_0;
assign _ptw_io_requestor_1_pmp_mask_1 = ptw__io_requestor_1_pmp_mask_1;
assign _ptw_io_requestor_1_pmp_mask_2 = ptw__io_requestor_1_pmp_mask_2;
assign _ptw_io_requestor_1_pmp_mask_3 = ptw__io_requestor_1_pmp_mask_3;
assign _ptw_io_requestor_1_pmp_mask_4 = ptw__io_requestor_1_pmp_mask_4;
assign _ptw_io_requestor_1_pmp_mask_5 = ptw__io_requestor_1_pmp_mask_5;
assign _ptw_io_requestor_1_pmp_mask_6 = ptw__io_requestor_1_pmp_mask_6;
assign _ptw_io_requestor_1_pmp_mask_7 = ptw__io_requestor_1_pmp_mask_7;
assign _ptw_io_requestor_1_customCSRs_csrs_0_value = ptw__io_requestor_1_customCSRs_csrs_0_value;
assign ptw__io_dpath_status_debug = _core_io_ptw_status_debug;
assign ptw__io_dpath_pmp_cfg_l_0 = _core_io_ptw_pmp_cfg_l_0;
assign ptw__io_dpath_pmp_cfg_l_1 = _core_io_ptw_pmp_cfg_l_1;
assign ptw__io_dpath_pmp_cfg_l_2 = _core_io_ptw_pmp_cfg_l_2;
assign ptw__io_dpath_pmp_cfg_l_3 = _core_io_ptw_pmp_cfg_l_3;
assign ptw__io_dpath_pmp_cfg_l_4 = _core_io_ptw_pmp_cfg_l_4;
assign ptw__io_dpath_pmp_cfg_l_5 = _core_io_ptw_pmp_cfg_l_5;
assign ptw__io_dpath_pmp_cfg_l_6 = _core_io_ptw_pmp_cfg_l_6;
assign ptw__io_dpath_pmp_cfg_l_7 = _core_io_ptw_pmp_cfg_l_7;
assign ptw__io_dpath_pmp_cfg_a_0 = _core_io_ptw_pmp_cfg_a_0;
assign ptw__io_dpath_pmp_cfg_a_1 = _core_io_ptw_pmp_cfg_a_1;
assign ptw__io_dpath_pmp_cfg_a_2 = _core_io_ptw_pmp_cfg_a_2;
assign ptw__io_dpath_pmp_cfg_a_3 = _core_io_ptw_pmp_cfg_a_3;
assign ptw__io_dpath_pmp_cfg_a_4 = _core_io_ptw_pmp_cfg_a_4;
assign ptw__io_dpath_pmp_cfg_a_5 = _core_io_ptw_pmp_cfg_a_5;
assign ptw__io_dpath_pmp_cfg_a_6 = _core_io_ptw_pmp_cfg_a_6;
assign ptw__io_dpath_pmp_cfg_a_7 = _core_io_ptw_pmp_cfg_a_7;
assign ptw__io_dpath_pmp_cfg_x_0 = _core_io_ptw_pmp_cfg_x_0;
assign ptw__io_dpath_pmp_cfg_x_1 = _core_io_ptw_pmp_cfg_x_1;
assign ptw__io_dpath_pmp_cfg_x_2 = _core_io_ptw_pmp_cfg_x_2;
assign ptw__io_dpath_pmp_cfg_x_3 = _core_io_ptw_pmp_cfg_x_3;
assign ptw__io_dpath_pmp_cfg_x_4 = _core_io_ptw_pmp_cfg_x_4;
assign ptw__io_dpath_pmp_cfg_x_5 = _core_io_ptw_pmp_cfg_x_5;
assign ptw__io_dpath_pmp_cfg_x_6 = _core_io_ptw_pmp_cfg_x_6;
assign ptw__io_dpath_pmp_cfg_x_7 = _core_io_ptw_pmp_cfg_x_7;
assign ptw__io_dpath_pmp_cfg_w_0 = _core_io_ptw_pmp_cfg_w_0;
assign ptw__io_dpath_pmp_cfg_w_1 = _core_io_ptw_pmp_cfg_w_1;
assign ptw__io_dpath_pmp_cfg_w_2 = _core_io_ptw_pmp_cfg_w_2;
assign ptw__io_dpath_pmp_cfg_w_3 = _core_io_ptw_pmp_cfg_w_3;
assign ptw__io_dpath_pmp_cfg_w_4 = _core_io_ptw_pmp_cfg_w_4;
assign ptw__io_dpath_pmp_cfg_w_5 = _core_io_ptw_pmp_cfg_w_5;
assign ptw__io_dpath_pmp_cfg_w_6 = _core_io_ptw_pmp_cfg_w_6;
assign ptw__io_dpath_pmp_cfg_w_7 = _core_io_ptw_pmp_cfg_w_7;
assign ptw__io_dpath_pmp_cfg_r_0 = _core_io_ptw_pmp_cfg_r_0;
assign ptw__io_dpath_pmp_cfg_r_1 = _core_io_ptw_pmp_cfg_r_1;
assign ptw__io_dpath_pmp_cfg_r_2 = _core_io_ptw_pmp_cfg_r_2;
assign ptw__io_dpath_pmp_cfg_r_3 = _core_io_ptw_pmp_cfg_r_3;
assign ptw__io_dpath_pmp_cfg_r_4 = _core_io_ptw_pmp_cfg_r_4;
assign ptw__io_dpath_pmp_cfg_r_5 = _core_io_ptw_pmp_cfg_r_5;
assign ptw__io_dpath_pmp_cfg_r_6 = _core_io_ptw_pmp_cfg_r_6;
assign ptw__io_dpath_pmp_cfg_r_7 = _core_io_ptw_pmp_cfg_r_7;
assign ptw__io_dpath_pmp_addr_0 = _core_io_ptw_pmp_addr_0;
assign ptw__io_dpath_pmp_addr_1 = _core_io_ptw_pmp_addr_1;
assign ptw__io_dpath_pmp_addr_2 = _core_io_ptw_pmp_addr_2;
assign ptw__io_dpath_pmp_addr_3 = _core_io_ptw_pmp_addr_3;
assign ptw__io_dpath_pmp_addr_4 = _core_io_ptw_pmp_addr_4;
assign ptw__io_dpath_pmp_addr_5 = _core_io_ptw_pmp_addr_5;
assign ptw__io_dpath_pmp_addr_6 = _core_io_ptw_pmp_addr_6;
assign ptw__io_dpath_pmp_addr_7 = _core_io_ptw_pmp_addr_7;
assign ptw__io_dpath_pmp_mask_0 = _core_io_ptw_pmp_mask_0;
assign ptw__io_dpath_pmp_mask_1 = _core_io_ptw_pmp_mask_1;
assign ptw__io_dpath_pmp_mask_2 = _core_io_ptw_pmp_mask_2;
assign ptw__io_dpath_pmp_mask_3 = _core_io_ptw_pmp_mask_3;
assign ptw__io_dpath_pmp_mask_4 = _core_io_ptw_pmp_mask_4;
assign ptw__io_dpath_pmp_mask_5 = _core_io_ptw_pmp_mask_5;
assign ptw__io_dpath_pmp_mask_6 = _core_io_ptw_pmp_mask_6;
assign ptw__io_dpath_pmp_mask_7 = _core_io_ptw_pmp_mask_7;
assign ptw__io_dpath_customCSRs_csrs_0_value = _core_io_ptw_customCSRs_csrs_0_value;
 
  
wire  core__clock;
wire  core__reset;
wire  core__io_hartid;
wire  core__io_interrupts_debug;
wire  core__io_interrupts_mtip;
wire  core__io_interrupts_msip;
wire  core__io_interrupts_meip;
wire  core__io_imem_might_request;
wire  core__io_imem_req_valid;
wire [33:0] core__io_imem_req_bits_pc;
wire  core__io_imem_req_bits_speculative;
wire  core__io_imem_resp_ready;
wire  core__io_imem_resp_valid;
wire [33:0] core__io_imem_resp_bits_pc;
wire [31:0] core__io_imem_resp_bits_data;
wire  core__io_imem_resp_bits_xcpt_pf_inst;
wire  core__io_imem_resp_bits_xcpt_gf_inst;
wire  core__io_imem_resp_bits_xcpt_ae_inst;
wire  core__io_imem_resp_bits_replay;
wire  core__io_imem_btb_update_valid;
wire  core__io_imem_bht_update_valid;
wire  core__io_imem_flush_icache;
wire  core__io_dmem_req_ready;
wire  core__io_dmem_req_valid;
wire [33:0] core__io_dmem_req_bits_addr;
wire [5:0] core__io_dmem_req_bits_tag;
wire [4:0] core__io_dmem_req_bits_cmd;
wire [1:0] core__io_dmem_req_bits_size;
wire  core__io_dmem_req_bits_signed;
wire  core__io_dmem_req_bits_dv;
wire  core__io_dmem_s1_kill;
wire [63:0] core__io_dmem_s1_data_data;
wire  core__io_dmem_s2_nack;
wire  core__io_dmem_resp_valid;
wire [5:0] core__io_dmem_resp_bits_tag;
wire [63:0] core__io_dmem_resp_bits_data;
wire  core__io_dmem_resp_bits_replay;
wire  core__io_dmem_resp_bits_has_data;
wire [63:0] core__io_dmem_resp_bits_data_word_bypass;
wire  core__io_dmem_replay_next;
wire  core__io_dmem_s2_xcpt_ma_ld;
wire  core__io_dmem_s2_xcpt_ma_st;
wire  core__io_dmem_s2_xcpt_pf_ld;
wire  core__io_dmem_s2_xcpt_pf_st;
wire  core__io_dmem_s2_xcpt_ae_ld;
wire  core__io_dmem_s2_xcpt_ae_st;
wire  core__io_dmem_ordered;
wire  core__io_dmem_perf_release;
wire  core__io_dmem_perf_grant;
wire  core__io_ptw_status_debug;
wire  core__io_ptw_pmp_cfg_l_0;
wire  core__io_ptw_pmp_cfg_l_1;
wire  core__io_ptw_pmp_cfg_l_2;
wire  core__io_ptw_pmp_cfg_l_3;
wire  core__io_ptw_pmp_cfg_l_4;
wire  core__io_ptw_pmp_cfg_l_5;
wire  core__io_ptw_pmp_cfg_l_6;
wire  core__io_ptw_pmp_cfg_l_7;
wire [1:0] core__io_ptw_pmp_cfg_a_0;
wire [1:0] core__io_ptw_pmp_cfg_a_1;
wire [1:0] core__io_ptw_pmp_cfg_a_2;
wire [1:0] core__io_ptw_pmp_cfg_a_3;
wire [1:0] core__io_ptw_pmp_cfg_a_4;
wire [1:0] core__io_ptw_pmp_cfg_a_5;
wire [1:0] core__io_ptw_pmp_cfg_a_6;
wire [1:0] core__io_ptw_pmp_cfg_a_7;
wire  core__io_ptw_pmp_cfg_x_0;
wire  core__io_ptw_pmp_cfg_x_1;
wire  core__io_ptw_pmp_cfg_x_2;
wire  core__io_ptw_pmp_cfg_x_3;
wire  core__io_ptw_pmp_cfg_x_4;
wire  core__io_ptw_pmp_cfg_x_5;
wire  core__io_ptw_pmp_cfg_x_6;
wire  core__io_ptw_pmp_cfg_x_7;
wire  core__io_ptw_pmp_cfg_w_0;
wire  core__io_ptw_pmp_cfg_w_1;
wire  core__io_ptw_pmp_cfg_w_2;
wire  core__io_ptw_pmp_cfg_w_3;
wire  core__io_ptw_pmp_cfg_w_4;
wire  core__io_ptw_pmp_cfg_w_5;
wire  core__io_ptw_pmp_cfg_w_6;
wire  core__io_ptw_pmp_cfg_w_7;
wire  core__io_ptw_pmp_cfg_r_0;
wire  core__io_ptw_pmp_cfg_r_1;
wire  core__io_ptw_pmp_cfg_r_2;
wire  core__io_ptw_pmp_cfg_r_3;
wire  core__io_ptw_pmp_cfg_r_4;
wire  core__io_ptw_pmp_cfg_r_5;
wire  core__io_ptw_pmp_cfg_r_6;
wire  core__io_ptw_pmp_cfg_r_7;
wire [29:0] core__io_ptw_pmp_addr_0;
wire [29:0] core__io_ptw_pmp_addr_1;
wire [29:0] core__io_ptw_pmp_addr_2;
wire [29:0] core__io_ptw_pmp_addr_3;
wire [29:0] core__io_ptw_pmp_addr_4;
wire [29:0] core__io_ptw_pmp_addr_5;
wire [29:0] core__io_ptw_pmp_addr_6;
wire [29:0] core__io_ptw_pmp_addr_7;
wire [31:0] core__io_ptw_pmp_mask_0;
wire [31:0] core__io_ptw_pmp_mask_1;
wire [31:0] core__io_ptw_pmp_mask_2;
wire [31:0] core__io_ptw_pmp_mask_3;
wire [31:0] core__io_ptw_pmp_mask_4;
wire [31:0] core__io_ptw_pmp_mask_5;
wire [31:0] core__io_ptw_pmp_mask_6;
wire [31:0] core__io_ptw_pmp_mask_7;
wire [63:0] core__io_ptw_customCSRs_csrs_0_value;
wire  core__io_wfi;
 
   wire  core__io_dmem_req_valid_0  ; 
   wire  core__div_io_resp_ready  ; 
   wire  core__take_pc_wb  ; 
   wire  core__take_pc_mem  ; 
   wire  core___div_io_req_ready  ; 
   wire  core___div_io_resp_valid  ; 
   wire[63:0]  core___div_io_resp_bits_data  ; 
   wire[4:0]  core___div_io_resp_bits_tag  ; 
   wire[63:0]  core___alu_io_out  ; 
   wire[63:0]  core___alu_io_adder_out  ; 
   wire  core___alu_io_cmp_out  ; 
   wire  core___bpu_io_xcpt_if  ; 
   wire  core___bpu_io_xcpt_ld  ; 
   wire  core___bpu_io_xcpt_st  ; 
   wire  core___bpu_io_debug_if  ; 
   wire  core___bpu_io_debug_ld  ; 
   wire  core___bpu_io_debug_st  ; 
   wire[63:0]  core___csr_io_rw_rdata  ; 
   wire  core___csr_io_decode_0_read_illegal  ; 
   wire  core___csr_io_decode_0_write_illegal  ; 
   wire  core___csr_io_decode_0_write_flush  ; 
   wire  core___csr_io_decode_0_system_illegal  ; 
   wire  core___csr_io_decode_0_virtual_access_illegal  ; 
   wire  core___csr_io_decode_0_virtual_system_illegal  ; 
   wire  core___csr_io_csr_stall  ; 
   wire  core___csr_io_eret  ; 
   wire  core___csr_io_singleStep  ; 
   wire  core___csr_io_status_debug  ; 
   wire[31:0]  core___csr_io_status_isa  ; 
   wire  core___csr_io_status_dv  ; 
   wire  core___csr_io_status_v  ; 
   wire[33:0]  core___csr_io_evec  ; 
   wire[63:0]  core___csr_io_time  ; 
   wire  core___csr_io_interrupt  ; 
   wire[63:0]  core___csr_io_interrupt_cause  ; 
   wire  core___csr_io_bp_0_control_action  ; 
   wire[1:0]  core___csr_io_bp_0_control_tmatch  ; 
   wire  core___csr_io_bp_0_control_x  ; 
   wire  core___csr_io_bp_0_control_w  ; 
   wire  core___csr_io_bp_0_control_r  ; 
   wire[32:0]  core___csr_io_bp_0_address  ; 
   wire  core___csr_io_inhibit_cycle  ; 
   wire  core___csr_io_trace_valid_0  ; 
   wire[33:0]  core___csr_io_trace_iaddr_0  ; 
   wire[31:0]  core___csr_io_trace_insn_0  ; 
   wire  core___csr_io_trace_exception_0  ; 
   wire[63:0]  core___csr_io_customCSRs_0_value  ; 
   wire[63:0]  core___rf_ext_R0_data  ; 
   wire[63:0]  core___rf_ext_R1_data  ; 
   wire[33:0]  core___ibuf_io_pc  ; 
   wire  core___ibuf_io_inst_0_valid  ; 
   wire  core___ibuf_io_inst_0_bits_xcpt0_pf_inst  ; 
   wire  core___ibuf_io_inst_0_bits_xcpt0_gf_inst  ; 
   wire  core___ibuf_io_inst_0_bits_xcpt0_ae_inst  ; 
   wire  core___ibuf_io_inst_0_bits_xcpt1_pf_inst  ; 
   wire  core___ibuf_io_inst_0_bits_xcpt1_gf_inst  ; 
   wire  core___ibuf_io_inst_0_bits_xcpt1_ae_inst  ; 
   wire  core___ibuf_io_inst_0_bits_replay  ; 
   wire  core___ibuf_io_inst_0_bits_rvc  ; 
   wire[31:0]  core___ibuf_io_inst_0_bits_inst_bits  ; 
   wire[4:0]  core___ibuf_io_inst_0_bits_inst_rd  ; 
   wire[4:0]  core___ibuf_io_inst_0_bits_inst_rs1  ; 
   wire[4:0]  core___ibuf_io_inst_0_bits_inst_rs2  ; 
   wire[31:0]  core___ibuf_io_inst_0_bits_raw  ; 
   reg  core__id_reg_pause  ; 
   reg  core__imem_might_request_reg  ; 
   reg  core__ex_ctrl_fp  ; 
   reg  core__ex_ctrl_rocc  ; 
   reg  core__ex_ctrl_branch  ; 
   reg  core__ex_ctrl_jal  ; 
   reg  core__ex_ctrl_jalr  ; 
   reg  core__ex_ctrl_rxs2  ; 
   reg  core__ex_ctrl_rxs1  ; 
   reg[1:0]  core__ex_ctrl_sel_alu2  ; 
   reg[1:0]  core__ex_ctrl_sel_alu1  ; 
   reg[2:0]  core__ex_ctrl_sel_imm  ; 
   reg  core__ex_ctrl_alu_dw  ; 
   reg[3:0]  core__ex_ctrl_alu_fn  ; 
   reg  core__ex_ctrl_mem  ; 
   reg[4:0]  core__ex_ctrl_mem_cmd  ; 
   reg  core__ex_ctrl_rfs1  ; 
   reg  core__ex_ctrl_rfs2  ; 
   reg  core__ex_ctrl_wfd  ; 
   reg  core__ex_ctrl_mul  ; 
   reg  core__ex_ctrl_div  ; 
   reg  core__ex_ctrl_wxd  ; 
   reg[2:0]  core__ex_ctrl_csr  ; 
   reg  core__ex_ctrl_fence_i  ; 
   reg  core__mem_ctrl_fp  ; 
   reg  core__mem_ctrl_rocc  ; 
   reg  core__mem_ctrl_branch  ; 
   reg  core__mem_ctrl_jal  ; 
   reg  core__mem_ctrl_jalr  ; 
   reg  core__mem_ctrl_rxs2  ; 
   reg  core__mem_ctrl_rxs1  ; 
   reg  core__mem_ctrl_mem  ; 
   reg  core__mem_ctrl_rfs1  ; 
   reg  core__mem_ctrl_rfs2  ; 
   reg  core__mem_ctrl_wfd  ; 
   reg  core__mem_ctrl_mul  ; 
   reg  core__mem_ctrl_div  ; 
   reg  core__mem_ctrl_wxd  ; 
   reg[2:0]  core__mem_ctrl_csr  ; 
   reg  core__mem_ctrl_fence_i  ; 
   reg  core__wb_ctrl_rocc  ; 
   reg  core__wb_ctrl_rxs2  ; 
   reg  core__wb_ctrl_rxs1  ; 
   reg  core__wb_ctrl_mem  ; 
   reg  core__wb_ctrl_rfs1  ; 
   reg  core__wb_ctrl_rfs2  ; 
   reg  core__wb_ctrl_wfd  ; 
   reg  core__wb_ctrl_div  ; 
   reg  core__wb_ctrl_wxd  ; 
   reg[2:0]  core__wb_ctrl_csr  ; 
   reg  core__wb_ctrl_fence_i  ; 
   reg  core__ex_reg_xcpt_interrupt  ; 
   reg  core__ex_reg_valid  ; 
   reg  core__ex_reg_rvc  ; 
   reg  core__ex_reg_xcpt  ; 
   reg  core__ex_reg_flush_pipe  ; 
   reg  core__ex_reg_load_use  ; 
   reg[63:0]  core__ex_reg_cause  ; 
   reg  core__ex_reg_replay  ; 
   reg[33:0]  core__ex_reg_pc  ; 
   reg[1:0]  core__ex_reg_mem_size  ; 
   reg[31:0]  core__ex_reg_inst  ; 
   reg[31:0]  core__ex_reg_raw_inst  ; 
   reg  core__mem_reg_xcpt_interrupt  ; 
   reg  core__mem_reg_valid  ; 
   reg  core__mem_reg_rvc  ; 
   reg  core__mem_reg_xcpt  ; 
   reg  core__mem_reg_replay  ; 
   reg  core__mem_reg_flush_pipe  ; 
   reg[63:0]  core__mem_reg_cause  ; 
   reg  core__mem_mem_cmd_bh  ; 
   reg  core__mem_reg_load  ; 
   reg  core__mem_reg_store  ; 
   reg[33:0]  core__mem_reg_pc  ; 
   reg[31:0]  core__mem_reg_inst  ; 
   reg  core__mem_reg_hls_or_dv  ; 
   reg[31:0]  core__mem_reg_raw_inst  ; 
   reg[63:0]  core__mem_reg_wdata  ; 
   reg[63:0]  core__mem_reg_rs2  ; 
   reg  core__mem_br_taken  ; 
   reg  core__wb_reg_valid  ; 
   reg  core__wb_reg_xcpt  ; 
   reg  core__wb_reg_replay  ; 
   reg  core__wb_reg_flush_pipe  ; 
   reg[63:0]  core__wb_reg_cause  ; 
   reg[33:0]  core__wb_reg_pc  ; 
   reg  core__wb_reg_hls_or_dv  ; 
   reg[31:0]  core__wb_reg_inst  ; 
   reg[31:0]  core__wb_reg_raw_inst  ; 
   reg[63:0]  core__wb_reg_wdata  ; 
   wire  core__ibuf_io_kill  =  core__take_pc_wb  |  core__take_pc_mem  ; 
   wire[29:0]  core__id_ctrl_decoder_decoded_invInputs  =~(  core___ibuf_io_inst_0_bits_inst_bits  [31:2]); 
   wire[6:0]  core___id_ctrl_decoder_decoded_T  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_4  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [11]}; 
   wire[6:0]  core___id_ctrl_decoder_decoded_T_6  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_8  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[8:0]  core___id_ctrl_decoder_decoded_T_12  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[5:0]  core___id_ctrl_decoder_decoded_T_14  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [4]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_18  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[14:0]  core___id_ctrl_decoder_decoded_T_22  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[12:0]  core___id_ctrl_decoder_decoded_T_26  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[14:0]  core___id_ctrl_decoder_decoded_T_28  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[8:0]  core___id_ctrl_decoder_decoded_T_36  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[9:0]  core___id_ctrl_decoder_decoded_T_38  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[6:0]  core___id_ctrl_decoder_decoded_T_40  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6]}; 
   wire[9:0]  core___id_ctrl_decoder_decoded_T_46  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[13:0]  core___id_ctrl_decoder_decoded_T_48  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[14:0]  core___id_ctrl_decoder_decoded_T_52  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[8:0]  core___id_ctrl_decoder_decoded_T_60  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_62  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [12]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_64  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13]}; 
   wire[10:0]  core___id_ctrl_decoder_decoded_T_68  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_74  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [13]}; 
   wire[8:0]  core___id_ctrl_decoder_decoded_T_76  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_86  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [14]}; 
   wire[14:0]  core___id_ctrl_decoder_decoded_T_88  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[14:0]  core___id_ctrl_decoder_decoded_T_92  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[14:0]  core___id_ctrl_decoder_decoded_T_98  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[13:0]  core___id_ctrl_decoder_decoded_T_130  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[12:0]  core___id_ctrl_decoder_decoded_T_136  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core___ibuf_io_inst_0_bits_inst_bits  [27],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[16:0]  core___id_ctrl_decoder_decoded_T_138  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [18],  core__id_ctrl_decoder_decoded_invInputs  [19],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [25],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[18:0]  core___id_ctrl_decoder_decoded_T_140  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [18],  core__id_ctrl_decoder_decoded_invInputs  [19],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [25],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[2:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T  ={&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_138  }; 
   wire[21:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_8  ={&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_8  ,&  core___id_ctrl_decoder_decoded_T_12  ,&  core___id_ctrl_decoder_decoded_T_14  ,&  core___id_ctrl_decoder_decoded_T_22  ,&  core___id_ctrl_decoder_decoded_T_26  ,&  core___id_ctrl_decoder_decoded_T_28  ,&  core___id_ctrl_decoder_decoded_T_38  ,&  core___id_ctrl_decoder_decoded_T_40  ,&  core___id_ctrl_decoder_decoded_T_48  ,&  core___id_ctrl_decoder_decoded_T_52  ,&  core___id_ctrl_decoder_decoded_T_62  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_74  ,&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_92  ,&  core___id_ctrl_decoder_decoded_T_98  ,&  core___id_ctrl_decoder_decoded_T_130  ,&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_138  }; 
   wire[2:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_10  ={&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_130  }; 
   wire[5:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_19  ={&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10]},&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_6  ,&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_140  }; 
   wire[20:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_45  ={&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_6  ,&  core___id_ctrl_decoder_decoded_T_12  ,&  core___id_ctrl_decoder_decoded_T_22  ,&  core___id_ctrl_decoder_decoded_T_26  ,&  core___id_ctrl_decoder_decoded_T_28  ,&  core___id_ctrl_decoder_decoded_T_36  ,&  core___id_ctrl_decoder_decoded_T_48  ,&  core___id_ctrl_decoder_decoded_T_52  ,&  core___id_ctrl_decoder_decoded_T_60  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_76  ,&  core___id_ctrl_decoder_decoded_T_86  ,&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_92  ,&  core___id_ctrl_decoder_decoded_T_98  ,&  core___id_ctrl_decoder_decoded_T_130  ,&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_138  }; 
   wire[11:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_47  ={&  core___id_ctrl_decoder_decoded_T_18  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]},&  core___id_ctrl_decoder_decoded_T_22  ,&  core___id_ctrl_decoder_decoded_T_26  ,&  core___id_ctrl_decoder_decoded_T_28  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_86  ,&  core___id_ctrl_decoder_decoded_T_98  ,&  core___id_ctrl_decoder_decoded_T_130  ,&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_138  }; 
   reg  core__id_reg_fence  ; 
   wire  core__id_mem_busy  =~  core__io_dmem_ordered  |  core__io_dmem_req_valid_0  ; 
   wire  core___io_rocc_cmd_valid_T  =  core__wb_reg_valid  &  core__wb_ctrl_rocc  ; 
   wire  core___dcache_kill_mem_T  =  core__mem_reg_valid  &  core__mem_ctrl_wxd  ; 
   wire  core___fp_data_hazard_ex_T_1  =  core__ex_reg_inst  [11:7]==  core___ibuf_io_inst_0_bits_inst_rs1  ; 
   wire  core___fp_data_hazard_mem_T_1  =  core__mem_reg_inst  [11:7]==  core___ibuf_io_inst_0_bits_inst_rs1  ; 
   wire  core___fp_data_hazard_ex_T_3  =  core__ex_reg_inst  [11:7]==  core___ibuf_io_inst_0_bits_inst_rs2  ; 
   wire  core___fp_data_hazard_mem_T_3  =  core__mem_reg_inst  [11:7]==  core___ibuf_io_inst_0_bits_inst_rs2  ; 
   reg  core__ex_reg_rs_bypass_0  ; 
   reg  core__ex_reg_rs_bypass_1  ; 
   reg[1:0]  core__ex_reg_rs_lsb_0  ; 
   reg[1:0]  core__ex_reg_rs_lsb_1  ; 
   reg[61:0]  core__ex_reg_rs_msb_0  ; 
   reg[61:0]  core__ex_reg_rs_msb_1  ; 
   reg[63:0]  core__casez_tmp  ; 
  always @(*)
       begin 
         casez (  core__ex_reg_rs_lsb_0  )
          2 'b00: 
              core__casez_tmp   =64'h0;
          2 'b01: 
              core__casez_tmp   =  core__mem_reg_wdata  ;
          2 'b10: 
              core__casez_tmp   =  core__wb_reg_wdata  ;
          default : 
              core__casez_tmp   =  core__io_dmem_resp_bits_data_word_bypass  ;
         endcase 
       end
  
   wire[63:0]  core__ex_rs_0  =  core__ex_reg_rs_bypass_0   ?   core__casez_tmp  :{  core__ex_reg_rs_msb_0  ,  core__ex_reg_rs_lsb_0  }; 
   reg[63:0]  core__casez_tmp_0  ; 
  always @(*)
       begin 
         casez (  core__ex_reg_rs_lsb_1  )
          2 'b00: 
              core__casez_tmp_0   =64'h0;
          2 'b01: 
              core__casez_tmp_0   =  core__mem_reg_wdata  ;
          2 'b10: 
              core__casez_tmp_0   =  core__wb_reg_wdata  ;
          default : 
              core__casez_tmp_0   =  core__io_dmem_resp_bits_data_word_bypass  ;
         endcase 
       end
  
   wire[63:0]  core__ex_rs_1  =  core__ex_reg_rs_bypass_1   ?   core__casez_tmp_0  :{  core__ex_reg_rs_msb_1  ,  core__ex_reg_rs_lsb_1  }; 
   reg[63:0]  core__casez_tmp_1  ; 
   wire[3:0]  core___ex_op2_T_1  =  core__ex_reg_rvc   ? 4'h2:4'h4; 
   wire  core___ex_imm_b0_T_4  =  core__ex_ctrl_sel_imm  ==3'h5; 
   wire  core__ex_imm_sign  =~  core___ex_imm_b0_T_4  &  core__ex_reg_inst  [31]; 
   wire  core___ex_imm_b4_1_T  =  core__ex_ctrl_sel_imm  ==3'h2; 
   wire  core___ex_imm_b4_1_T_2  =  core__ex_ctrl_sel_imm  ==3'h1; 
   wire  core___ex_imm_b0_T  =  core__ex_ctrl_sel_imm  ==3'h0; 
  always @(*)
       begin 
         casez (  core__ex_ctrl_sel_alu2  )
          2 'b00: 
              core__casez_tmp_1   =64'h0;
          2 'b01: 
              core__casez_tmp_1   ={{60{  core___ex_op2_T_1  [3]}},  core___ex_op2_T_1  };
          2 'b10: 
              core__casez_tmp_1   =  core__ex_rs_1  ;
          default : 
              core__casez_tmp_1   ={{33{  core__ex_imm_sign  }},  core___ex_imm_b4_1_T   ?   core__ex_reg_inst  [30:20]:{11{  core__ex_imm_sign  }},  core__ex_ctrl_sel_imm  !=3'h2&  core__ex_ctrl_sel_imm  !=3'h3 ? {8{  core__ex_imm_sign  }}:  core__ex_reg_inst  [19:12],~(  core___ex_imm_b4_1_T  |  core___ex_imm_b0_T_4  )&(  core__ex_ctrl_sel_imm  ==3'h3 ?   core__ex_reg_inst  [20]:  core___ex_imm_b4_1_T_2   ?   core__ex_reg_inst  [7]:  core__ex_imm_sign  ),  core___ex_imm_b4_1_T  |  core___ex_imm_b0_T_4   ? 6'h0:  core__ex_reg_inst  [30:25],  core___ex_imm_b4_1_T   ? 4'h0:  core___ex_imm_b0_T  |  core___ex_imm_b4_1_T_2   ?   core__ex_reg_inst  [11:8]:  core___ex_imm_b0_T_4   ?   core__ex_reg_inst  [19:16]:  core__ex_reg_inst  [24:21],  core___ex_imm_b0_T   ?   core__ex_reg_inst  [7]:  core__ex_ctrl_sel_imm  ==3'h4 ?   core__ex_reg_inst  [20]:  core___ex_imm_b0_T_4  &  core__ex_reg_inst  [15]};
         endcase 
       end
  
   wire  core__div_io_req_valid  =  core__ex_reg_valid  &  core__ex_ctrl_div  ; 
   wire  core__ex_pc_valid  =  core__ex_reg_valid  |  core__ex_reg_replay  |  core__ex_reg_xcpt_interrupt  ; 
   wire  core__wb_dcache_miss  =  core__wb_ctrl_mem  &~  core__io_dmem_resp_valid  ; 
   wire  core___mem_cfi_taken_T  =  core__mem_ctrl_branch  &  core__mem_br_taken  ; 
   wire[3:0]  core___mem_br_target_T_6  =  core__mem_reg_rvc   ? 4'h2:4'h4; 
   wire[31:0]  core___mem_br_target_T_8  =  core___mem_cfi_taken_T   ? {{20{  core__mem_reg_inst  [31]}},  core__mem_reg_inst  [7],  core__mem_reg_inst  [30:25],  core__mem_reg_inst  [11:8],1'h0}:  core__mem_ctrl_jal   ? {{12{  core__mem_reg_inst  [31]}},  core__mem_reg_inst  [19:12],  core__mem_reg_inst  [20],  core__mem_reg_inst  [30:21],1'h0}:{{28{  core___mem_br_target_T_6  [3]}},  core___mem_br_target_T_6  }; 
   wire[33:0]  core___mem_br_target_T_9  =  core__mem_reg_pc  +{{2{  core___mem_br_target_T_8  [31]}},  core___mem_br_target_T_8  }; 
   wire[33:0]  core___mem_npc_T_4  =  core__mem_ctrl_jalr   ? {  core__mem_reg_wdata  [63:33]==31'h0|(&(  core__mem_reg_wdata  [63:33])) ?   core__mem_reg_wdata  [33]:~(  core__mem_reg_wdata  [32]),  core__mem_reg_wdata  [32:0]}:  core___mem_br_target_T_9  ; 
   wire[33:0]  core__mem_npc  =  core___mem_npc_T_4  &34'h3FFFFFFFE; 
   wire  core__mem_cfi_taken  =  core___mem_cfi_taken_T  |  core__mem_ctrl_jalr  |  core__mem_ctrl_jal  ; 
  assign   core__take_pc_mem  =  core__mem_reg_valid  &~  core__mem_reg_xcpt  &  core__mem_cfi_taken  ; 
   reg[63:0]  core__casez_tmp_2  ; 
  always @(*)
       begin 
         casez (  core__ex_ctrl_rocc   ? 2'h3:  core__ex_reg_mem_size  )
          2 'b00: 
              core__casez_tmp_2   ={2{{2{{2{  core__ex_rs_1  [7:0]}}}}}};
          2 'b01: 
              core__casez_tmp_2   ={2{{2{  core__ex_rs_1  [15:0]}}}};
          2 'b10: 
              core__casez_tmp_2   ={2{  core__ex_rs_1  [31:0]}};
          default : 
              core__casez_tmp_2   =  core__ex_rs_1  ;
         endcase 
       end
  
   wire  core__mem_debug_breakpoint  =  core__mem_reg_load  &  core___bpu_io_debug_ld  |  core__mem_reg_store  &  core___bpu_io_debug_st  ; 
   wire  core__mem_ldst_xcpt  =  core__mem_debug_breakpoint  |  core__mem_reg_load  &  core___bpu_io_xcpt_ld  |  core__mem_reg_store  &  core___bpu_io_xcpt_st  ; 
   wire  core__dcache_kill_mem  =  core___dcache_kill_mem_T  &  core__io_dmem_replay_next  ; 
   wire  core__killm_common  =  core__dcache_kill_mem  |  core__take_pc_wb  |  core__mem_reg_xcpt  |~  core__mem_reg_valid  ; 
   reg  core__div_io_kill_REG  ; 
   wire  core___GEN  =  core__wb_reg_valid  &  core__wb_ctrl_mem  ; 
   wire  core___GEN_0  =  core___GEN  &  core__io_dmem_s2_xcpt_pf_st  ; 
   wire  core___GEN_1  =  core___GEN  &  core__io_dmem_s2_xcpt_pf_ld  ; 
   wire  core___GEN_2  =  core___GEN  &  core__io_dmem_s2_xcpt_ae_st  ; 
   wire  core___GEN_3  =  core___GEN  &  core__io_dmem_s2_xcpt_ae_ld  ; 
   wire  core___GEN_4  =  core___GEN  &  core__io_dmem_s2_xcpt_ma_st  ; 
   wire  core__wb_xcpt  =  core__wb_reg_xcpt  |  core___GEN_0  |  core___GEN_1  |  core___GEN_2  |  core___GEN_3  |  core___GEN_4  |  core___GEN  &  core__io_dmem_s2_xcpt_ma_ld  ; 
   wire  core__wb_wxd  =  core__wb_reg_valid  &  core__wb_ctrl_wxd  ; 
   wire  core__wb_set_sboard  =  core__wb_ctrl_div  |  core__wb_dcache_miss  |  core__wb_ctrl_rocc  ; 
   wire  core__replay_wb_common  =  core__io_dmem_s2_nack  |  core__wb_reg_replay  ; 
   wire  core___replay_wb_T  =  core__replay_wb_common  |  core___io_rocc_cmd_valid_T  ; 
  assign   core__take_pc_wb  =  core___replay_wb_T  |  core__wb_xcpt  |  core___csr_io_eret  |  core__wb_reg_flush_pipe  ; 
   wire  core__dmem_resp_valid  =  core__io_dmem_resp_valid  &  core__io_dmem_resp_bits_has_data  ; 
   wire  core___GEN_5  =  core__dmem_resp_valid  &  core__io_dmem_resp_bits_replay  &~(  core__io_dmem_resp_bits_tag  [0]); 
  assign   core__div_io_resp_ready  =~  core___GEN_5  &~  core__wb_wxd  ; 
   wire[4:0]  core__ll_waddr  =  core___GEN_5   ?   core__io_dmem_resp_bits_tag  [5:1]:  core___div_io_resp_bits_tag  ; 
   wire  core__ll_wen  =  core___GEN_5  |  core__div_io_resp_ready  &  core___div_io_resp_valid  ; 
   wire  core__wb_valid  =  core__wb_reg_valid  &~  core___replay_wb_T  &~  core__wb_xcpt  ; 
   wire  core__wb_wen  =  core__wb_valid  &  core__wb_ctrl_wxd  ; 
   wire  core__rf_wen  =  core__wb_wen  |  core__ll_wen  ; 
   wire[4:0]  core__rf_waddr  =  core__ll_wen   ?   core__ll_waddr  :  core__wb_reg_inst  [11:7]; 
   wire[63:0]  core__rf_wdata  =  core__dmem_resp_valid  &~(  core__io_dmem_resp_bits_tag  [0]) ?   core__io_dmem_resp_bits_data  :  core__ll_wen   ?   core___div_io_resp_bits_data  :(|  core__wb_ctrl_csr  ) ?   core___csr_io_rw_rdata  :  core__wb_reg_wdata  ; 
   wire[63:0]  core__id_rs_0  =  core__rf_wen  &(|  core__rf_waddr  )&  core__rf_waddr  ==  core___ibuf_io_inst_0_bits_inst_rs1   ?   core__rf_wdata  :  core___rf_ext_R1_data  ; 
   wire[63:0]  core__id_rs_1  =  core__rf_wen  &(|  core__rf_waddr  )&  core__rf_waddr  ==  core___ibuf_io_inst_0_bits_inst_rs2   ?   core__rf_wdata  :  core___rf_ext_R0_data  ; 
   wire  core___csr_io_htval_htval_valid_imem_T  =  core__wb_reg_cause  ==64'h14; 
   wire  core__tval_any_addr  =~  core__wb_reg_xcpt  |  core__wb_reg_cause  ==64'h3|  core__wb_reg_cause  ==64'h1|  core__wb_reg_cause  ==64'hC|  core___csr_io_htval_htval_valid_imem_T  ; 
   wire  core___GEN_6  =(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_45  )&(|  core___ibuf_io_inst_0_bits_inst_rs1  ); 
   wire  core___GEN_7  =(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_47  )&(|  core___ibuf_io_inst_0_bits_inst_rs2  ); 
   wire  core___GEN_8  =(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_8  )&(|  core___ibuf_io_inst_0_bits_inst_rd  ); 
   reg[31:0]  core___r  ; 
   wire[31:0]  core__r  ={  core___r  [31:1],1'h0}; 
   wire[31:0]  core___id_sboard_hazard_T  =  core__r  >>  core___ibuf_io_inst_0_bits_inst_rs1  ; 
   wire[31:0]  core___id_sboard_hazard_T_7  =  core__r  >>  core___ibuf_io_inst_0_bits_inst_rs2  ; 
   wire[31:0]  core___id_sboard_hazard_T_14  =  core__r  >>  core___ibuf_io_inst_0_bits_inst_rd  ; 
   wire  core__data_hazard_mem  =  core__mem_ctrl_wxd  &(  core___GEN_6  &  core___fp_data_hazard_mem_T_1  |  core___GEN_7  &  core___fp_data_hazard_mem_T_3  |  core___GEN_8  &  core___ibuf_io_inst_0_bits_inst_rd  ==  core__mem_reg_inst  [11:7]); 
   reg  core__dcache_blocked_blocked  ; 
   reg  core__rocc_blocked  ; 
   wire  core___ctrl_stalld_T_28  =  core__ex_reg_valid  &  core__ex_ctrl_wxd  &(  core___GEN_6  &  core___fp_data_hazard_ex_T_1  |  core___GEN_7  &  core___fp_data_hazard_ex_T_3  |  core___GEN_8  &  core___ibuf_io_inst_0_bits_inst_rd  ==  core__ex_reg_inst  [11:7])&((|  core__ex_ctrl_csr  )|  core__ex_ctrl_jalr  |  core__ex_ctrl_mem  |  core__ex_ctrl_mul  |  core__ex_ctrl_div  |  core__ex_ctrl_fp  |  core__ex_ctrl_rocc  )|  core__mem_reg_valid  &  core__data_hazard_mem  &((|  core__mem_ctrl_csr  )|  core__mem_ctrl_mem  &  core__mem_mem_cmd_bh  |  core__mem_ctrl_mul  |  core__mem_ctrl_div  |  core__mem_ctrl_fp  |  core__mem_ctrl_rocc  )|  core__wb_reg_valid  &  core__wb_ctrl_wxd  &(  core___GEN_6  &  core___ibuf_io_inst_0_bits_inst_rs1  ==  core__wb_reg_inst  [11:7]|  core___GEN_7  &  core___ibuf_io_inst_0_bits_inst_rs2  ==  core__wb_reg_inst  [11:7]|  core___GEN_8  &  core___ibuf_io_inst_0_bits_inst_rd  ==  core__wb_reg_inst  [11:7])&  core__wb_set_sboard  |  core___GEN_6  &  core___id_sboard_hazard_T  [0]&~(  core__ll_wen  &  core__ll_waddr  ==  core___ibuf_io_inst_0_bits_inst_rs1  )|  core___GEN_7  &  core___id_sboard_hazard_T_7  [0]&~(  core__ll_wen  &  core__ll_waddr  ==  core___ibuf_io_inst_0_bits_inst_rs2  )|  core___GEN_8  &  core___id_sboard_hazard_T_14  [0]&~(  core__ll_wen  &  core__ll_waddr  ==  core___ibuf_io_inst_0_bits_inst_rd  )|  core___csr_io_singleStep  &(  core__ex_reg_valid  |  core__mem_reg_valid  |  core__wb_reg_valid  )|(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_19  )&  core__dcache_blocked_blocked  &~  core__io_dmem_perf_grant  |(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_10  )&(~(  core___div_io_req_ready  |  core___div_io_resp_valid  &~  core__wb_wxd  )|  core__div_io_req_valid  )|  core__id_mem_busy  &((|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T  )&  core___ibuf_io_inst_0_bits_inst_bits  [25]|(&  core___id_ctrl_decoder_decoded_T_46  )|  core__id_reg_fence  &(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_19  ))|  core___csr_io_csr_stall  |  core__id_reg_pause  ; 
   wire  core__ctrl_killd  =~  core___ibuf_io_inst_0_valid  |  core___ibuf_io_inst_0_bits_replay  |  core__ibuf_io_kill  |  core___ctrl_stalld_T_28  |  core___csr_io_interrupt  ; 
  assign   core__io_dmem_req_valid_0  =  core__ex_reg_valid  &  core__ex_ctrl_mem  ; 
   reg[63:0]  core__coreMonitorBundle_rd0val_REG  ; 
   reg[63:0]  core__coreMonitorBundle_rd0val_REG_1  ; 
   reg[63:0]  core__coreMonitorBundle_rd1val_REG  ; 
   reg[63:0]  core__coreMonitorBundle_rd1val_REG_1  ; 
   wire  core__coreMonitorBundle_wrenx  =  core__wb_wen  &~  core__wb_set_sboard  ; 
   wire  core___GEN_9  =  core__wb_ctrl_rxs1  |  core__wb_ctrl_rfs1  ; 
   wire  core___GEN_10  =  core__wb_ctrl_rxs2  |  core__wb_ctrl_rfs2  ; 
  always @( posedge   core__clock  )
       begin 
         if (~  core__reset  &  core__wb_reg_xcpt  &  core___csr_io_htval_htval_valid_imem_T  )
            begin 
              if (1)$display("Assertion failed\n    at RocketCore.scala:718 assert(!htval_valid_imem || io.imem.gpa.valid)\n");
              if (1)$display("");
            end 
         if ((1)&  core___csr_io_trace_valid_0  &~  core__reset  )
            begin $fwrite(32'h80000001,"C%d: %d [%d] pc=[%x] W[r%d=%x][%d] R[r%d=%x] R[r%d=%x] inst=[%x] DASM(%x)\n",  core__io_hartid  ,  core___csr_io_time  [31:0],  core___csr_io_trace_valid_0  &~  core___csr_io_trace_exception_0  ,{{30{  core___csr_io_trace_iaddr_0  [33]}},  core___csr_io_trace_iaddr_0  },  core__wb_ctrl_wxd  |  core__wb_ctrl_wfd   ?   core__wb_reg_inst  [11:7]:5'h0,  core__coreMonitorBundle_wrenx   ?   core__rf_wdata  :64'h0,  core__coreMonitorBundle_wrenx  ,  core___GEN_9   ?   core__wb_reg_inst  [19:15]:5'h0,  core___GEN_9   ?   core__coreMonitorBundle_rd0val_REG_1  :64'h0,  core___GEN_10   ?   core__wb_reg_inst  [24:20]:5'h0,  core___GEN_10   ?   core__coreMonitorBundle_rd1val_REG_1  :64'h0,  core___csr_io_trace_insn_0  ,  core___csr_io_trace_insn_0  );
            end 
       end
  
   wire[7:0]  core___id_ctrl_decoder_decoded_T_32  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [11]}; 
   wire[14:0]  core___id_ctrl_decoder_decoded_T_50  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[15:0]  core___id_ctrl_decoder_decoded_T_54  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[15:0]  core___id_ctrl_decoder_decoded_T_94  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_104  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [14]}; 
   wire[8:0]  core___id_ctrl_decoder_decoded_T_108  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [14]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_114  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [14]}; 
   wire[8:0]  core___id_ctrl_decoder_decoded_T_118  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [14]}; 
   wire[13:0]  core___id_ctrl_decoder_decoded_T_146  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core___ibuf_io_inst_0_bits_inst_bits  [27],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[2:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_16  ={&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_138  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core___ibuf_io_inst_0_bits_inst_bits  [31]}}; 
   wire[2:0]  core___GEN_11  ={  core___ibuf_io_inst_0_bits_xcpt1_pf_inst  ,  core___ibuf_io_inst_0_bits_xcpt1_gf_inst  ,  core___ibuf_io_inst_0_bits_xcpt1_ae_inst  }; 
   wire  core___GEN_12  =  core___bpu_io_xcpt_if  |(|{  core___ibuf_io_inst_0_bits_xcpt0_pf_inst  ,  core___ibuf_io_inst_0_bits_xcpt0_gf_inst  ,  core___ibuf_io_inst_0_bits_xcpt0_ae_inst  }); 
   wire[31:0]  core__inst  =  core___ibuf_io_inst_0_bits_rvc   ? {16'h0,  core___ibuf_io_inst_0_bits_raw  [15:0]}:  core___ibuf_io_inst_0_bits_raw  ; 
   wire  core___mem_reg_store_T_3  =  core__ex_ctrl_mem_cmd  ==5'h7; 
   wire  core___mem_reg_store_T_5  =  core__ex_ctrl_mem_cmd  ==5'h4; 
   wire  core___mem_reg_store_T_6  =  core__ex_ctrl_mem_cmd  ==5'h9; 
   wire  core___mem_reg_store_T_7  =  core__ex_ctrl_mem_cmd  ==5'hA; 
   wire  core___mem_reg_store_T_8  =  core__ex_ctrl_mem_cmd  ==5'hB; 
   wire  core___mem_reg_store_T_12  =  core__ex_ctrl_mem_cmd  ==5'h8; 
   wire  core___mem_reg_store_T_13  =  core__ex_ctrl_mem_cmd  ==5'hC; 
   wire  core___mem_reg_store_T_14  =  core__ex_ctrl_mem_cmd  ==5'hD; 
   wire  core___mem_reg_store_T_15  =  core__ex_ctrl_mem_cmd  ==5'hE; 
   wire  core___mem_reg_store_T_16  =  core__ex_ctrl_mem_cmd  ==5'hF; 
   wire[31:0]  core___GEN_13  =  core__r  &~(  core__ll_wen   ? 32'h1<<  core__ll_waddr  :32'h0); 
   wire  core___GEN_14  =  core__wb_set_sboard  &  core__wb_wen  ; 
   wire[8:0]  core___id_ctrl_decoder_decoded_T_10  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]}; 
   wire[7:0]  core___id_ctrl_decoder_decoded_T_56  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11]}; 
   wire[27:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_53  ={&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_6  ,&  core___id_ctrl_decoder_decoded_T_10  ,&  core___id_ctrl_decoder_decoded_T_12  ,&  core___id_ctrl_decoder_decoded_T_14  ,&  core___id_ctrl_decoder_decoded_T_22  ,&  core___id_ctrl_decoder_decoded_T_26  ,&  core___id_ctrl_decoder_decoded_T_28  ,&  core___id_ctrl_decoder_decoded_T_36  ,&  core___id_ctrl_decoder_decoded_T_40  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core__id_ctrl_decoder_decoded_invInputs  [19],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_48  ,&  core___id_ctrl_decoder_decoded_T_52  ,&  core___id_ctrl_decoder_decoded_T_56  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_74  ,&  core___id_ctrl_decoder_decoded_T_86  ,&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_92  ,&  core___id_ctrl_decoder_decoded_T_98  ,&  core___id_ctrl_decoder_decoded_T_130  ,&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_140  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core___ibuf_io_inst_0_bits_inst_bits  [20],  core__id_ctrl_decoder_decoded_invInputs  [19],  core___ibuf_io_inst_0_bits_inst_bits  [22],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core__id_ctrl_decoder_decoded_invInputs  [18],  core___ibuf_io_inst_0_bits_inst_bits  [21],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core___ibuf_io_inst_0_bits_inst_bits  [29],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core__id_ctrl_decoder_decoded_invInputs  [18],  core___ibuf_io_inst_0_bits_inst_bits  [21],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core___ibuf_io_inst_0_bits_inst_bits  [24],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core___ibuf_io_inst_0_bits_inst_bits  [27],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core___ibuf_io_inst_0_bits_inst_bits  [29],  core___ibuf_io_inst_0_bits_inst_bits  [30],  core__id_ctrl_decoder_decoded_invInputs  [29]}}; 
   wire[2:0]  core__id_ctrl_csr  ={|{&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core__id_ctrl_decoder_decoded_invInputs  [19],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_62  ,&  core___id_ctrl_decoder_decoded_T_74  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core___ibuf_io_inst_0_bits_inst_bits  [20],  core__id_ctrl_decoder_decoded_invInputs  [19],  core___ibuf_io_inst_0_bits_inst_bits  [22],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core__id_ctrl_decoder_decoded_invInputs  [18],  core___ibuf_io_inst_0_bits_inst_bits  [21],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core__id_ctrl_decoder_decoded_invInputs  [22],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core___ibuf_io_inst_0_bits_inst_bits  [29],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [5],  core__id_ctrl_decoder_decoded_invInputs  [6],  core__id_ctrl_decoder_decoded_invInputs  [7],  core__id_ctrl_decoder_decoded_invInputs  [8],  core__id_ctrl_decoder_decoded_invInputs  [9],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [13],  core__id_ctrl_decoder_decoded_invInputs  [14],  core__id_ctrl_decoder_decoded_invInputs  [15],  core__id_ctrl_decoder_decoded_invInputs  [16],  core__id_ctrl_decoder_decoded_invInputs  [17],  core__id_ctrl_decoder_decoded_invInputs  [18],  core___ibuf_io_inst_0_bits_inst_bits  [21],  core__id_ctrl_decoder_decoded_invInputs  [20],  core__id_ctrl_decoder_decoded_invInputs  [21],  core___ibuf_io_inst_0_bits_inst_bits  [24],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core___ibuf_io_inst_0_bits_inst_bits  [27],  core___ibuf_io_inst_0_bits_inst_bits  [28],  core___ibuf_io_inst_0_bits_inst_bits  [29],  core___ibuf_io_inst_0_bits_inst_bits  [30],  core__id_ctrl_decoder_decoded_invInputs  [29]}},&  core___id_ctrl_decoder_decoded_T_74  ,&  core___id_ctrl_decoder_decoded_T_62  }; 
   wire  core___id_csr_ren_T  =  core__id_ctrl_csr  ==3'h6; 
   wire  core__id_csr_en  =  core___id_csr_ren_T  |(&  core__id_ctrl_csr  )|  core__id_ctrl_csr  ==3'h5; 
   wire  core__id_system_insn  =  core__id_ctrl_csr  ==3'h4; 
   wire  core__id_csr_ren  =(  core___id_csr_ren_T  |(&  core__id_ctrl_csr  ))&~(|  core___ibuf_io_inst_0_bits_inst_rs1  ); 
   wire  core__id_illegal_insn  =~(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_53  )|(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_10  )&~(  core___csr_io_status_isa  [12])|(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T  )&~(  core___csr_io_status_isa  [0])|  core___ibuf_io_inst_0_bits_rvc  &~(  core___csr_io_status_isa  [2])|  core__id_csr_en  &(  core___csr_io_decode_0_read_illegal  |~  core__id_csr_ren  &  core___csr_io_decode_0_write_illegal  )|~  core___ibuf_io_inst_0_bits_rvc  &  core__id_system_insn  &  core___csr_io_decode_0_system_illegal  ; 
   wire  core__id_virtual_insn  =(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_53  )&(  core__id_csr_en  &~(~  core__id_csr_ren  &  core___csr_io_decode_0_write_illegal  )&  core___csr_io_decode_0_virtual_access_illegal  |~  core___ibuf_io_inst_0_bits_rvc  &  core__id_system_insn  &  core___csr_io_decode_0_virtual_system_illegal  ); 
   wire  core__id_xcpt  =  core___csr_io_interrupt  |  core___bpu_io_debug_if  |  core___bpu_io_xcpt_if  |  core___ibuf_io_inst_0_bits_xcpt0_pf_inst  |  core___ibuf_io_inst_0_bits_xcpt0_gf_inst  |  core___ibuf_io_inst_0_bits_xcpt0_ae_inst  |  core___ibuf_io_inst_0_bits_xcpt1_pf_inst  |  core___ibuf_io_inst_0_bits_xcpt1_gf_inst  |  core___ibuf_io_inst_0_bits_xcpt1_ae_inst  |  core__id_virtual_insn  |  core__id_illegal_insn  ; 
   wire  core___GEN_15  =  core__ex_reg_valid  &  core__ex_ctrl_wxd  ; 
   wire  core___GEN_16  =  core___dcache_kill_mem_T  &~  core__mem_ctrl_mem  ; 
   wire  core__id_bypass_src_1_1  =  core___GEN_15  &  core___fp_data_hazard_ex_T_3  ; 
   wire  core__id_bypass_src_1_2  =  core___GEN_16  &  core___fp_data_hazard_mem_T_3  ; 
   wire  core__do_bypass_1  =~(|  core___ibuf_io_inst_0_bits_inst_rs2  )|  core__id_bypass_src_1_1  |  core__id_bypass_src_1_2  |  core___dcache_kill_mem_T  &  core___fp_data_hazard_mem_T_3  ; 
   wire  core___GEN_17  =(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_47  )&~  core__do_bypass_1  ; 
   wire  core__replay_ex  =  core__ex_reg_replay  |  core__ex_reg_valid  &(  core__ex_ctrl_mem  &~  core__io_dmem_req_ready  |  core__ex_ctrl_div  &~  core___div_io_req_ready  |  core__wb_dcache_miss  &  core__ex_reg_load_use  ); 
   wire  core__ctrl_killx  =  core__ibuf_io_kill  |  core__replay_ex  |~  core__ex_reg_valid  ; 
   wire  core__mem_pc_valid  =  core__mem_reg_valid  |  core__mem_reg_replay  |  core__mem_reg_xcpt_interrupt  ; 
   wire  core___mem_npc_misaligned_T_3  =~(  core___csr_io_status_isa  [2])&  core___mem_npc_T_4  [1]; 
   wire  core___GEN_18  =  core__mem_reg_valid  &  core__mem_reg_flush_pipe  ; 
   wire  core___GEN_19  =  core___GEN_18  |~  core__ex_pc_valid  ; 
   wire  core___GEN_20  =  core__ex_ctrl_jalr  &  core___csr_io_status_debug  ; 
   wire  core___GEN_21  =  core__mem_reg_xcpt_interrupt  |  core__mem_reg_xcpt  ; 
   wire  core___GEN_22  =  core__mem_reg_valid  &  core___mem_npc_misaligned_T_3  ; 
   wire  core__mem_xcpt  =  core___GEN_21  |  core___GEN_22  |  core__mem_reg_valid  &  core__mem_ldst_xcpt  ; 
   wire  core___ctrl_killm_T  =  core__killm_common  |  core__mem_xcpt  ; 
   wire[15:0]  core___id_ctrl_decoder_decoded_T_154  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core___ibuf_io_inst_0_bits_inst_bits  [30],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[15:0]  core___id_ctrl_decoder_decoded_T_158  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core___ibuf_io_inst_0_bits_inst_bits  [30],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[15:0]  core___id_ctrl_decoder_decoded_T_160  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core___ibuf_io_inst_0_bits_inst_bits  [30],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[15:0]  core___id_ctrl_decoder_decoded_T_162  ={  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core___ibuf_io_inst_0_bits_inst_bits  [30],  core__id_ctrl_decoder_decoded_invInputs  [29]}; 
   wire[2:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_12  ={&  core___id_ctrl_decoder_decoded_T_18  ,&  core___id_ctrl_decoder_decoded_T_146  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core___ibuf_io_inst_0_bits_inst_bits  [29]}}; 
   wire[2:0]  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_14  ={&  core___id_ctrl_decoder_decoded_T_138  ,&  core___id_ctrl_decoder_decoded_T_146  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core___ibuf_io_inst_0_bits_inst_bits  [30]}}; 
   wire  core__id_bypass_src_0_1  =  core___GEN_15  &  core___fp_data_hazard_ex_T_1  ; 
   wire  core__id_bypass_src_0_2  =  core___GEN_16  &  core___fp_data_hazard_mem_T_1  ; 
   wire  core__do_bypass  =~(|  core___ibuf_io_inst_0_bits_inst_rs1  )|  core__id_bypass_src_0_1  |  core__id_bypass_src_0_2  |  core___dcache_kill_mem_T  &  core___fp_data_hazard_mem_T_1  ; 
   wire  core___GEN_23  =(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_45  )&~  core__do_bypass  ; 
   wire  core___GEN_24  =  core__id_illegal_insn  |  core__id_virtual_insn  ; 
   wire[3:0]  core__id_ctrl_alu_fn  ={|{&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_86  ,&  core___id_ctrl_decoder_decoded_T_154  ,&  core___id_ctrl_decoder_decoded_T_158  ,&  core___id_ctrl_decoder_decoded_T_160  ,&  core___id_ctrl_decoder_decoded_T_162  },|{&  core___id_ctrl_decoder_decoded_T_64  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10],  core___ibuf_io_inst_0_bits_inst_bits  [14]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_86  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [3],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_130  },|{&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [13]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [14]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [14]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_154  ,&  core___id_ctrl_decoder_decoded_T_158  ,&  core___id_ctrl_decoder_decoded_T_160  ,&  core___id_ctrl_decoder_decoded_T_162  },|{&  core___id_ctrl_decoder_decoded_T_48  ,&  core___id_ctrl_decoder_decoded_T_52  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11]},&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_92  ,&  core___id_ctrl_decoder_decoded_T_98  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core__id_ctrl_decoder_decoded_invInputs  [2],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core___ibuf_io_inst_0_bits_inst_bits  [6],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [14]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [13],  core___ibuf_io_inst_0_bits_inst_bits  [14]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]},&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core___ibuf_io_inst_0_bits_inst_bits  [25],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [28],  core__id_ctrl_decoder_decoded_invInputs  [29]}}}; 
  always @( posedge   core__clock  )
       begin  
          core__id_reg_pause   <=~(  core___csr_io_time  [4:0]==5'h0|  core___csr_io_inhibit_cycle  |  core__io_dmem_perf_release  |  core__ibuf_io_kill  )&(~  core__ctrl_killd  &(&  core___id_ctrl_decoder_decoded_T_10  )&  core___ibuf_io_inst_0_bits_inst_bits  [23:20]==4'h0|  core__id_reg_pause  ); 
          core__imem_might_request_reg   <=  core__ex_pc_valid  |  core__mem_pc_valid  |  core___csr_io_customCSRs_0_value  [1]; 
          core__ex_ctrl_fp   <=  core__ctrl_killd  &  core__ex_ctrl_fp  ; 
          core__ex_ctrl_rocc   <=  core__ctrl_killd  &  core__ex_ctrl_rocc  ;
         if (~  core__ctrl_killd  )
            begin  
               core__ex_ctrl_branch   <=|{&  core___id_ctrl_decoder_decoded_T_32  ,&  core___id_ctrl_decoder_decoded_T_86  }; 
               core__ex_ctrl_jal   <=&  core___id_ctrl_decoder_decoded_T_40  ; 
               core__ex_ctrl_jalr   <=&  core___id_ctrl_decoder_decoded_T_38  ; 
               core__ex_ctrl_rxs2   <=|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_47  ; 
               core__ex_ctrl_rxs1   <=|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_45  ; 
               core__ex_ctrl_sel_alu2   <=  core__id_xcpt   ? (  core___GEN_12   ? 2'h0:{1'h0,|  core___GEN_11  }):{|{&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_6  ,&  core___id_ctrl_decoder_decoded_T_12  ,&  core___id_ctrl_decoder_decoded_T_14  ,&  core___id_ctrl_decoder_decoded_T_22  ,&  core___id_ctrl_decoder_decoded_T_26  ,&  core___id_ctrl_decoder_decoded_T_28  ,&  core___id_ctrl_decoder_decoded_T_32  ,&  core___id_ctrl_decoder_decoded_T_36  ,&  core___id_ctrl_decoder_decoded_T_48  ,&  core___id_ctrl_decoder_decoded_T_52  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_92  ,&  core___id_ctrl_decoder_decoded_T_98  ,&  core___id_ctrl_decoder_decoded_T_104  ,&  core___id_ctrl_decoder_decoded_T_114  ,&  core___id_ctrl_decoder_decoded_T_130  },|{&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_6  ,&  core___id_ctrl_decoder_decoded_T_12  ,&  core___id_ctrl_decoder_decoded_T_14  ,&  core___id_ctrl_decoder_decoded_T_38  ,&  core___id_ctrl_decoder_decoded_T_40  ,&  core___id_ctrl_decoder_decoded_T_50  ,&  core___id_ctrl_decoder_decoded_T_54  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_94  ,&  core___id_ctrl_decoder_decoded_T_108  ,&  core___id_ctrl_decoder_decoded_T_118  }}; 
               core__ex_ctrl_sel_alu1   <=  core__id_xcpt   ? (  core___GEN_12  |(|  core___GEN_11  ) ? 2'h2:2'h1):{|{&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core___ibuf_io_inst_0_bits_inst_bits  [2],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core__id_ctrl_decoder_decoded_invInputs  [3],  core__id_ctrl_decoder_decoded_invInputs  [4]},&  core___id_ctrl_decoder_decoded_T_40  },|{&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_6  ,&  core___id_ctrl_decoder_decoded_T_12  ,&  core___id_ctrl_decoder_decoded_T_22  ,&  core___id_ctrl_decoder_decoded_T_26  ,&  core___id_ctrl_decoder_decoded_T_28  ,&  core___id_ctrl_decoder_decoded_T_36  ,&  core___id_ctrl_decoder_decoded_T_48  ,&  core___id_ctrl_decoder_decoded_T_52  ,&  core___id_ctrl_decoder_decoded_T_60  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_76  ,&  core___id_ctrl_decoder_decoded_T_86  ,&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_92  ,&  core___id_ctrl_decoder_decoded_T_98  ,&  core___id_ctrl_decoder_decoded_T_130  ,&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_138  }}; 
               core__ex_ctrl_sel_imm   <={|{&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_8  ,&  core___id_ctrl_decoder_decoded_T_12  ,&  core___id_ctrl_decoder_decoded_T_38  ,&  core___id_ctrl_decoder_decoded_T_50  ,&  core___id_ctrl_decoder_decoded_T_54  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_88  ,&  core___id_ctrl_decoder_decoded_T_94  ,&  core___id_ctrl_decoder_decoded_T_108  ,&  core___id_ctrl_decoder_decoded_T_118  },|{&  core___id_ctrl_decoder_decoded_T_14  ,&  core___id_ctrl_decoder_decoded_T_40  },|{&  core___id_ctrl_decoder_decoded_T_32  ,&  core___id_ctrl_decoder_decoded_T_40  ,&  core___id_ctrl_decoder_decoded_T_104  ,&  core___id_ctrl_decoder_decoded_T_114  }}; 
               core__ex_ctrl_alu_dw   <=  core__id_xcpt  |(|{&  core___id_ctrl_decoder_decoded_T  ,&  core___id_ctrl_decoder_decoded_T_4  ,&  core___id_ctrl_decoder_decoded_T_6  ,&  core___id_ctrl_decoder_decoded_T_14  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core__id_ctrl_decoder_decoded_invInputs  [10],  core__id_ctrl_decoder_decoded_invInputs  [11],  core__id_ctrl_decoder_decoded_invInputs  [12],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_26  ,&  core___id_ctrl_decoder_decoded_T_36  ,&  core___id_ctrl_decoder_decoded_T_40  ,&  core___id_ctrl_decoder_decoded_T_48  ,&  core___id_ctrl_decoder_decoded_T_56  ,&  core___id_ctrl_decoder_decoded_T_64  ,&  core___id_ctrl_decoder_decoded_T_68  ,&  core___id_ctrl_decoder_decoded_T_74  ,&  core___id_ctrl_decoder_decoded_T_86  ,&  core___id_ctrl_decoder_decoded_T_88  ,&{  core___ibuf_io_inst_0_bits_inst_bits  [0],  core___ibuf_io_inst_0_bits_inst_bits  [1],  core__id_ctrl_decoder_decoded_invInputs  [0],  core__id_ctrl_decoder_decoded_invInputs  [1],  core___ibuf_io_inst_0_bits_inst_bits  [4],  core___ibuf_io_inst_0_bits_inst_bits  [5],  core__id_ctrl_decoder_decoded_invInputs  [4],  core___ibuf_io_inst_0_bits_inst_bits  [12],  core__id_ctrl_decoder_decoded_invInputs  [11],  core___ibuf_io_inst_0_bits_inst_bits  [14],  core__id_ctrl_decoder_decoded_invInputs  [23],  core__id_ctrl_decoder_decoded_invInputs  [24],  core__id_ctrl_decoder_decoded_invInputs  [25],  core__id_ctrl_decoder_decoded_invInputs  [26],  core__id_ctrl_decoder_decoded_invInputs  [27],  core__id_ctrl_decoder_decoded_invInputs  [29]},&  core___id_ctrl_decoder_decoded_T_136  ,&  core___id_ctrl_decoder_decoded_T_138  }); 
               core__ex_ctrl_alu_fn   <=  core__id_xcpt   ? 4'h0:  core__id_ctrl_alu_fn  ; 
               core__ex_ctrl_mem   <=|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_19  ; 
               core__ex_ctrl_mem_cmd   <={1'h0,&  core___id_ctrl_decoder_decoded_T_68  ,|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_16  ,|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_14  ,|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_12  }; 
               core__ex_ctrl_div   <=|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_10  ; 
               core__ex_ctrl_wxd   <=|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_8  ; 
               core__ex_ctrl_csr   <=  core__id_system_insn  &(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_19  ) ? 3'h0:  core__id_csr_ren   ? 3'h2:  core__id_ctrl_csr  ; 
               core__ex_ctrl_fence_i   <=&  core___id_ctrl_decoder_decoded_T_46  ; 
               core__ex_reg_rvc   <=  core__id_xcpt  &(|  core___GEN_11  )|  core___ibuf_io_inst_0_bits_rvc  ; 
               core__ex_reg_flush_pipe   <=(&  core___id_ctrl_decoder_decoded_T_46  )|  core__id_system_insn  |  core__id_csr_en  &~  core__id_csr_ren  &  core___csr_io_decode_0_write_flush  ; 
               core__ex_reg_load_use   <=  core__mem_reg_valid  &  core__data_hazard_mem  &  core__mem_ctrl_mem  ; 
               core__ex_reg_mem_size   <={&  core___id_ctrl_decoder_decoded_T_68  ,|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_16  ,|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_14  ,|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T_12  }==4'h5 ? {|  core___ibuf_io_inst_0_bits_inst_rs2  ,|  core___ibuf_io_inst_0_bits_inst_rs1  }:  core___ibuf_io_inst_0_bits_inst_bits  [13:12]; 
               core__ex_reg_rs_bypass_0   <=~  core___GEN_24  &  core__do_bypass  ; 
               core__ex_reg_rs_bypass_1   <=  core__do_bypass_1  ; 
               core__ex_reg_rs_lsb_0   <=  core___GEN_24   ?   core__inst  [1:0]:  core___GEN_23   ?   core__id_rs_0  [1:0]:(|  core___ibuf_io_inst_0_bits_inst_rs1  ) ? (  core__id_bypass_src_0_1   ? 2'h1:{1'h1,~  core__id_bypass_src_0_2  }):2'h0; 
               core__ex_reg_rs_lsb_1   <=  core___GEN_17   ?   core__id_rs_1  [1:0]:(|  core___ibuf_io_inst_0_bits_inst_rs2  ) ? (  core__id_bypass_src_1_1   ? 2'h1:{1'h1,~  core__id_bypass_src_1_2  }):2'h0;
              if (  core___GEN_24  ) 
                  core__ex_reg_rs_msb_0   <={32'h0,  core__inst  [31:2]};
               else 
                 if (  core___GEN_23  ) 
                     core__ex_reg_rs_msb_0   <=  core__id_rs_0  [63:2];
            end  
          core__ex_ctrl_rfs1   <=  core__ctrl_killd  &  core__ex_ctrl_rfs1  ; 
          core__ex_ctrl_rfs2   <=  core__ctrl_killd  &  core__ex_ctrl_rfs2  ; 
          core__ex_ctrl_wfd   <=  core__ctrl_killd  &  core__ex_ctrl_wfd  ; 
          core__ex_ctrl_mul   <=  core__ctrl_killd  &  core__ex_ctrl_mul  ;
         if (  core___GEN_19  )
            begin 
            end 
          else 
            begin  
               core__mem_ctrl_fp   <=  core__ex_ctrl_fp  ; 
               core__mem_ctrl_rocc   <=  core__ex_ctrl_rocc  ; 
               core__mem_ctrl_branch   <=  core__ex_ctrl_branch  ; 
               core__mem_ctrl_jal   <=  core__ex_ctrl_jal  ; 
               core__mem_ctrl_jalr   <=  core__ex_ctrl_jalr  ; 
               core__mem_ctrl_rxs2   <=  core__ex_ctrl_rxs2  ; 
               core__mem_ctrl_rxs1   <=  core__ex_ctrl_rxs1  ; 
               core__mem_ctrl_mem   <=  core__ex_ctrl_mem  ; 
               core__mem_ctrl_rfs1   <=  core__ex_ctrl_rfs1  ; 
               core__mem_ctrl_rfs2   <=  core__ex_ctrl_rfs2  ; 
               core__mem_ctrl_wfd   <=  core__ex_ctrl_wfd  ; 
               core__mem_ctrl_mul   <=  core__ex_ctrl_mul  ; 
               core__mem_ctrl_div   <=  core__ex_ctrl_div  ; 
               core__mem_ctrl_wxd   <=  core__ex_ctrl_wxd  ; 
               core__mem_ctrl_csr   <=  core__ex_ctrl_csr  ; 
               core__mem_ctrl_fence_i   <=  core___GEN_20  |  core__ex_ctrl_fence_i  ;
            end 
         if (  core__mem_pc_valid  )
            begin  
               core__wb_ctrl_rocc   <=  core__mem_ctrl_rocc  ; 
               core__wb_ctrl_rxs2   <=  core__mem_ctrl_rxs2  ; 
               core__wb_ctrl_rxs1   <=  core__mem_ctrl_rxs1  ; 
               core__wb_ctrl_mem   <=  core__mem_ctrl_mem  ; 
               core__wb_ctrl_rfs1   <=  core__mem_ctrl_rfs1  ; 
               core__wb_ctrl_rfs2   <=  core__mem_ctrl_rfs2  ; 
               core__wb_ctrl_wfd   <=  core__mem_ctrl_wfd  ; 
               core__wb_ctrl_div   <=  core__mem_ctrl_div  ; 
               core__wb_ctrl_wxd   <=  core__mem_ctrl_wxd  ; 
               core__wb_ctrl_csr   <=  core__mem_ctrl_csr  ; 
               core__wb_ctrl_fence_i   <=  core__mem_ctrl_fence_i  ; 
               core__wb_reg_cause   <=  core___GEN_21   ?   core__mem_reg_cause  :{60'h0,  core___GEN_22   ? 4'h0:  core__mem_debug_breakpoint   ? 4'hE:4'h3}; 
               core__wb_reg_pc   <=  core__mem_reg_pc  ; 
               core__wb_reg_hls_or_dv   <=  core__mem_reg_hls_or_dv  ; 
               core__wb_reg_inst   <=  core__mem_reg_inst  ; 
               core__wb_reg_raw_inst   <=  core__mem_reg_raw_inst  ; 
               core__wb_reg_wdata   <=~  core__mem_reg_xcpt  &  core__mem_ctrl_fp  &  core__mem_ctrl_wxd   ? 64'h0:~  core__mem_reg_xcpt  &(  core__mem_ctrl_jalr  ^  core___mem_npc_misaligned_T_3  ) ? {{30{  core___mem_br_target_T_9  [33]}},  core___mem_br_target_T_9  }:  core__mem_reg_wdata  ;
            end  
          core__ex_reg_xcpt_interrupt   <=~  core__ibuf_io_kill  &  core___ibuf_io_inst_0_valid  &  core___csr_io_interrupt  ; 
          core__ex_reg_valid   <=~  core__ctrl_killd  ; 
          core__ex_reg_xcpt   <=~  core__ctrl_killd  &  core__id_xcpt  ;
         if (~  core__ctrl_killd  |  core___csr_io_interrupt  |  core___ibuf_io_inst_0_bits_replay  )
            begin  
               core__ex_reg_cause   <=  core___csr_io_interrupt   ?   core___csr_io_interrupt_cause  :{59'h0,  core___bpu_io_debug_if   ? 5'hE:  core___bpu_io_xcpt_if   ? 5'h3:  core___ibuf_io_inst_0_bits_xcpt0_pf_inst   ? 5'hC:  core___ibuf_io_inst_0_bits_xcpt0_gf_inst   ? 5'h14:  core___ibuf_io_inst_0_bits_xcpt0_ae_inst   ? 5'h1:  core___ibuf_io_inst_0_bits_xcpt1_pf_inst   ? 5'hC:  core___ibuf_io_inst_0_bits_xcpt1_gf_inst   ? 5'h14:  core___ibuf_io_inst_0_bits_xcpt1_ae_inst   ? 5'h1:  core__id_virtual_insn   ? 5'h16:5'h2}; 
               core__ex_reg_pc   <=  core___ibuf_io_pc  ; 
               core__ex_reg_inst   <=  core___ibuf_io_inst_0_bits_inst_bits  ; 
               core__ex_reg_raw_inst   <=  core___ibuf_io_inst_0_bits_raw  ;
            end  
          core__ex_reg_replay   <=~  core__ibuf_io_kill  &  core___ibuf_io_inst_0_valid  &  core___ibuf_io_inst_0_bits_replay  ; 
          core__mem_reg_xcpt_interrupt   <=~  core__ibuf_io_kill  &  core__ex_reg_xcpt_interrupt  ; 
          core__mem_reg_valid   <=~  core__ctrl_killx  ;
         if (  core___GEN_19  )
            begin 
            end 
          else  
             core__mem_reg_rvc   <=  core__ex_reg_rvc  ; 
          core__mem_reg_xcpt   <=~  core__ctrl_killx  &(  core__ex_reg_xcpt_interrupt  |  core__ex_reg_xcpt  ); 
          core__mem_reg_replay   <=~  core__ibuf_io_kill  &  core__replay_ex  ;
         if (  core___GEN_19  )
            begin 
            end 
          else 
            begin  
               core__mem_reg_flush_pipe   <=  core___GEN_20  |  core__ex_reg_flush_pipe  ; 
               core__mem_reg_cause   <=  core__ex_reg_cause  ; 
               core__mem_mem_cmd_bh   <=  core___mem_reg_store_T_3  |~(  core__ex_reg_mem_size  [1]); 
               core__mem_reg_load   <=  core__ex_ctrl_mem  &(  core__ex_ctrl_mem_cmd  ==5'h0|  core__ex_ctrl_mem_cmd  ==5'h10|  core__ex_ctrl_mem_cmd  ==5'h6|  core___mem_reg_store_T_3  |  core___mem_reg_store_T_5  |  core___mem_reg_store_T_6  |  core___mem_reg_store_T_7  |  core___mem_reg_store_T_8  |  core___mem_reg_store_T_12  |  core___mem_reg_store_T_13  |  core___mem_reg_store_T_14  |  core___mem_reg_store_T_15  |  core___mem_reg_store_T_16  ); 
               core__mem_reg_store   <=  core__ex_ctrl_mem  &(  core__ex_ctrl_mem_cmd  ==5'h1|  core__ex_ctrl_mem_cmd  ==5'h11|  core___mem_reg_store_T_3  |  core___mem_reg_store_T_5  |  core___mem_reg_store_T_6  |  core___mem_reg_store_T_7  |  core___mem_reg_store_T_8  |  core___mem_reg_store_T_12  |  core___mem_reg_store_T_13  |  core___mem_reg_store_T_14  |  core___mem_reg_store_T_15  |  core___mem_reg_store_T_16  ); 
               core__mem_reg_pc   <=  core__ex_reg_pc  ; 
               core__mem_reg_inst   <=  core__ex_reg_inst  ; 
               core__mem_reg_hls_or_dv   <=  core___csr_io_status_dv  ; 
               core__mem_reg_raw_inst   <=  core__ex_reg_raw_inst  ; 
               core__mem_reg_wdata   <=  core___alu_io_out  ;
            end 
         if (  core___GEN_18  |~(  core__ex_pc_valid  &  core__ex_ctrl_rxs2  &(  core__ex_ctrl_mem  |  core__ex_ctrl_rocc  )))
            begin 
            end 
          else  
             core__mem_reg_rs2   <=  core__casez_tmp_2  ;
         if (  core___GEN_19  )
            begin 
            end 
          else  
             core__mem_br_taken   <=  core___alu_io_cmp_out  ; 
          core__wb_reg_valid   <=~  core___ctrl_killm_T  ; 
          core__wb_reg_xcpt   <=  core__mem_xcpt  &~  core__take_pc_wb  ; 
          core__wb_reg_replay   <=(  core__dcache_kill_mem  |  core__mem_reg_replay  )&~  core__take_pc_wb  ; 
          core__wb_reg_flush_pipe   <=~  core___ctrl_killm_T  &  core__mem_reg_flush_pipe  ;
         if (~  core__ctrl_killd  &  core___GEN_17  ) 
             core__ex_reg_rs_msb_1   <=  core__id_rs_1  [63:2]; 
          core__div_io_kill_REG   <=  core___div_io_req_ready  &  core__div_io_req_valid  ; 
          core__dcache_blocked_blocked   <=~  core__io_dmem_req_ready  &~  core__io_dmem_perf_grant  &(  core__dcache_blocked_blocked  |  core__io_dmem_req_valid_0  |  core__io_dmem_s2_nack  ); 
          core__rocc_blocked   <=~  core__wb_xcpt  &(  core___io_rocc_cmd_valid_T  &~  core__replay_wb_common  |  core__rocc_blocked  ); 
          core__coreMonitorBundle_rd0val_REG   <=  core__ex_rs_0  ; 
          core__coreMonitorBundle_rd0val_REG_1   <=  core__coreMonitorBundle_rd0val_REG  ; 
          core__coreMonitorBundle_rd1val_REG   <=  core__ex_rs_1  ; 
          core__coreMonitorBundle_rd1val_REG_1   <=  core__coreMonitorBundle_rd1val_REG  ;
         if (  core__reset  )
            begin  
               core__id_reg_fence   <=1'h0; 
               core___r   <=32'h0;
            end 
          else 
            begin  
               core__id_reg_fence   <=~  core__ctrl_killd  &((&  core___id_ctrl_decoder_decoded_T_10  )|(|  core___id_ctrl_decoder_decoded_orMatrixOutputs_T  )&  core___ibuf_io_inst_0_bits_inst_bits  [26])|  core__id_mem_busy  &  core__id_reg_fence  ;
              if (  core__ll_wen  |  core___GEN_14  ) 
                  core___r   <=  core___GEN_13  |(  core___GEN_14   ? 32'h1<<  core__wb_reg_inst  [11:7]:32'h0);
               else 
                 if (  core__ll_wen  ) 
                     core___r   <=  core___GEN_13  ;
            end 
       end
   
  
wire  core__ibuf__clock;
wire  core__ibuf__reset;
wire  core__ibuf__io_imem_ready;
wire  core__ibuf__io_imem_valid;
wire [33:0] core__ibuf__io_imem_bits_pc;
wire [31:0] core__ibuf__io_imem_bits_data;
wire  core__ibuf__io_imem_bits_xcpt_pf_inst;
wire  core__ibuf__io_imem_bits_xcpt_gf_inst;
wire  core__ibuf__io_imem_bits_xcpt_ae_inst;
wire  core__ibuf__io_imem_bits_replay;
wire  core__ibuf__io_kill;
wire [33:0] core__ibuf__io_pc;
wire  core__ibuf__io_inst_0_ready;
wire  core__ibuf__io_inst_0_valid;
wire  core__ibuf__io_inst_0_bits_xcpt0_pf_inst;
wire  core__ibuf__io_inst_0_bits_xcpt0_gf_inst;
wire  core__ibuf__io_inst_0_bits_xcpt0_ae_inst;
wire  core__ibuf__io_inst_0_bits_xcpt1_pf_inst;
wire  core__ibuf__io_inst_0_bits_xcpt1_gf_inst;
wire  core__ibuf__io_inst_0_bits_xcpt1_ae_inst;
wire  core__ibuf__io_inst_0_bits_replay;
wire  core__ibuf__io_inst_0_bits_rvc;
wire [31:0] core__ibuf__io_inst_0_bits_inst_bits;
wire [4:0] core__ibuf__io_inst_0_bits_inst_rd;
wire [4:0] core__ibuf__io_inst_0_bits_inst_rs1;
wire [4:0] core__ibuf__io_inst_0_bits_inst_rs2;
wire [31:0] core__ibuf__io_inst_0_bits_raw;
 
   wire[1:0]  core__ibuf__nReady  ; 
   wire  core__ibuf___exp_io_rvc  ; 
   reg  core__ibuf__nBufValid  ; 
   reg[33:0]  core__ibuf__buf_pc  ; 
   reg[31:0]  core__ibuf__buf_data  ; 
   reg  core__ibuf__buf_xcpt_pf_inst  ; 
   reg  core__ibuf__buf_xcpt_gf_inst  ; 
   reg  core__ibuf__buf_xcpt_ae_inst  ; 
   reg  core__ibuf__buf_replay  ; 
   wire[1:0]  core__ibuf___GEN  ={1'h0,  core__ibuf__io_imem_bits_pc  [1]}; 
   wire[1:0]  core__ibuf___nIC_T_2  =2'h2-  core__ibuf___GEN  ; 
   wire[1:0]  core__ibuf___GEN_0  ={1'h0,  core__ibuf__nBufValid  }; 
   wire[1:0]  core__ibuf___nICReady_T  =  core__ibuf__nReady  -  core__ibuf___GEN_0  ; 
   wire  core__ibuf___nBufValid_T  =  core__ibuf__nReady  >=  core__ibuf___GEN_0  ; 
   wire[1:0]  core__ibuf___nBufValid_T_6  =  core__ibuf___nIC_T_2  -  core__ibuf___nICReady_T  ; 
   wire[190:0]  core__ibuf___icData_T_4  ={63'h0,{2{{2{  core__ibuf__io_imem_bits_data  [31:16]}}}},  core__ibuf__io_imem_bits_data  ,{2{  core__ibuf__io_imem_bits_data  [15:0]}}}<<{185'h0,  core__ibuf___GEN_0  -2'h2-  core__ibuf___GEN  ,4'h0}; 
   wire[62:0]  core__ibuf___icMask_T_2  =63'hFFFFFFFF<<{58'h0,  core__ibuf__nBufValid  ,4'h0}; 
   wire[31:0]  core__ibuf__inst  =  core__ibuf___icData_T_4  [95:64]&  core__ibuf___icMask_T_2  [31:0]|  core__ibuf__buf_data  &~(  core__ibuf___icMask_T_2  [31:0]); 
   wire[3:0]  core__ibuf___valid_T  =4'h1<<(  core__ibuf__io_imem_valid   ?   core__ibuf___nIC_T_2  :2'h0)+  core__ibuf___GEN_0  ; 
   wire[1:0]  core__ibuf___valid_T_1  =  core__ibuf___valid_T  [1:0]-2'h1; 
   wire[1:0]  core__ibuf___bufMask_T_1  =(2'h1<<  core__ibuf___GEN_0  )-2'h1; 
   wire[1:0]  core__ibuf__buf_replay_0  =  core__ibuf__buf_replay   ?   core__ibuf___bufMask_T_1  :2'h0; 
   wire[1:0]  core__ibuf__ic_replay  =  core__ibuf__buf_replay_0  |(  core__ibuf__io_imem_bits_replay   ?   core__ibuf___valid_T_1  &~  core__ibuf___bufMask_T_1  :2'h0); 
   wire  core__ibuf__full_insn  =  core__ibuf___exp_io_rvc  |  core__ibuf___valid_T_1  [1]|  core__ibuf__buf_replay_0  [0]; 
   wire[2:0]  core__ibuf___io_inst_0_bits_xcpt1_T_5  =  core__ibuf___exp_io_rvc   ? 3'h0:{  core__ibuf___bufMask_T_1  [1] ?   core__ibuf__buf_xcpt_pf_inst  :  core__ibuf__io_imem_bits_xcpt_pf_inst  ,  core__ibuf___bufMask_T_1  [1] ?   core__ibuf__buf_xcpt_gf_inst  :  core__ibuf__io_imem_bits_xcpt_gf_inst  ,  core__ibuf___bufMask_T_1  [1] ?   core__ibuf__buf_xcpt_ae_inst  :  core__ibuf__io_imem_bits_xcpt_ae_inst  }; 
  assign   core__ibuf__nReady  =  core__ibuf__full_insn   ? (  core__ibuf___exp_io_rvc   ? 2'h1:2'h2):2'h0; 
   wire[63:0]  core__ibuf___buf_data_T_1  ={{2{  core__ibuf__io_imem_bits_data  [31:16]}},  core__ibuf__io_imem_bits_data  }>>{58'h0,  core__ibuf___GEN  +  core__ibuf___nICReady_T  ,4'h0}; 
   wire  core__ibuf___GEN_1  =  core__ibuf__io_imem_valid  &  core__ibuf___nBufValid_T  &  core__ibuf___nICReady_T  <  core__ibuf___nIC_T_2  &~(  core__ibuf___nBufValid_T_6  [1]); 
  always @( posedge   core__ibuf__clock  )
       begin 
         if (  core__ibuf__reset  ) 
             core__ibuf__nBufValid   <=1'h0;
          else  
             core__ibuf__nBufValid   <=~  core__ibuf__io_kill  &(  core__ibuf__io_inst_0_ready   ? (  core__ibuf___GEN_1   ?   core__ibuf___nBufValid_T_6  [0]:~(  core__ibuf___nBufValid_T  |~  core__ibuf__nBufValid  )&  core__ibuf__nBufValid  -  core__ibuf__nReady  [0]):  core__ibuf__nBufValid  );
         if (  core__ibuf__io_inst_0_ready  &  core__ibuf___GEN_1  )
            begin  
               core__ibuf__buf_pc   <=  core__ibuf__io_imem_bits_pc  &34'h3FFFFFFFC|  core__ibuf__io_imem_bits_pc  +{31'h0,  core__ibuf___nICReady_T  ,1'h0}&34'h3; 
               core__ibuf__buf_data   <={16'h0,  core__ibuf___buf_data_T_1  [15:0]}; 
               core__ibuf__buf_xcpt_pf_inst   <=  core__ibuf__io_imem_bits_xcpt_pf_inst  ; 
               core__ibuf__buf_xcpt_gf_inst   <=  core__ibuf__io_imem_bits_xcpt_gf_inst  ; 
               core__ibuf__buf_xcpt_ae_inst   <=  core__ibuf__io_imem_bits_xcpt_ae_inst  ; 
               core__ibuf__buf_replay   <=  core__ibuf__io_imem_bits_replay  ;
            end 
       end
   
  
wire [31:0] core__ibuf__exp__io_in;
wire [31:0] core__ibuf__exp__io_out_bits;
wire [4:0] core__ibuf__exp__io_out_rd;
wire [4:0] core__ibuf__exp__io_out_rs1;
wire [4:0] core__ibuf__exp__io_out_rs2;
wire  core__ibuf__exp__io_rvc;
 
   reg[2:0]  core__ibuf__exp__casez_tmp  ; 
   wire[2:0]  core__ibuf__exp___io_out_s_funct_T_2  ={  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:5]}; 
   wire[2:0]  core__ibuf__exp___io_out_s_funct_T_4  ={  core__ibuf__exp___io_out_s_funct_T_2  ==3'h1,2'h0}; 
  always @(*)
       begin 
         casez (  core__ibuf__exp___io_out_s_funct_T_2  )
          3 'b000: 
              core__ibuf__exp__casez_tmp   =  core__ibuf__exp___io_out_s_funct_T_4  ;
          3 'b001: 
              core__ibuf__exp__casez_tmp   =  core__ibuf__exp___io_out_s_funct_T_4  ;
          3 'b010: 
              core__ibuf__exp__casez_tmp   =3'h6;
          3 'b011: 
              core__ibuf__exp__casez_tmp   =3'h7;
          3 'b100: 
              core__ibuf__exp__casez_tmp   =3'h0;
          3 'b101: 
              core__ibuf__exp__casez_tmp   =3'h0;
          3 'b110: 
              core__ibuf__exp__casez_tmp   =3'h2;
          default : 
              core__ibuf__exp__casez_tmp   =3'h3;
         endcase 
       end
  
   wire[3:0]  core__ibuf__exp___GEN  ={4{  core__ibuf__exp__io_in  [12]}}; 
   wire[6:0]  core__ibuf__exp__io_out_s_load_opc  =(|(  core__ibuf__exp__io_in  [11:7])) ? 7'h3:7'h1F; 
   wire[4:0]  core__ibuf__exp___io_out_T_2  ={  core__ibuf__exp__io_in  [1:0],  core__ibuf__exp__io_in  [15:13]}; 
   wire  core__ibuf__exp___io_out_T_29  =  core__ibuf__exp___io_out_T_2  ==5'hE; 
   wire  core__ibuf__exp___io_out_T_31  =  core__ibuf__exp___io_out_T_2  ==5'hF; 
   wire  core__ibuf__exp___io_out_T_33  =  core__ibuf__exp___io_out_T_2  ==5'h10; 
   wire  core__ibuf__exp___io_out_T_35  =  core__ibuf__exp___io_out_T_2  ==5'h11; 
   wire  core__ibuf__exp___io_out_T_37  =  core__ibuf__exp___io_out_T_2  ==5'h12; 
   wire  core__ibuf__exp___io_out_T_39  =  core__ibuf__exp___io_out_T_2  ==5'h13; 
   wire  core__ibuf__exp___io_out_T_41  =  core__ibuf__exp___io_out_T_2  ==5'h14; 
   wire[31:0]  core__ibuf__exp___io_out_T_42_bits  =  core__ibuf__exp___io_out_T_41   ? {7'h0,  core__ibuf__exp__io_in  [12] ? ((|(  core__ibuf__exp__io_in  [6:2])) ? {  core__ibuf__exp__io_in  [6:2],  core__ibuf__exp__io_in  [11:7],3'h0,  core__ibuf__exp__io_in  [11:7],7'h33}:(|(  core__ibuf__exp__io_in  [11:7])) ? {  core__ibuf__exp__io_in  [6:2],  core__ibuf__exp__io_in  [11:7],15'hE7}:{  core__ibuf__exp__io_in  [6:3],1'h1,  core__ibuf__exp__io_in  [11:7],15'h73}):{  core__ibuf__exp__io_in  [6:2],(|(  core__ibuf__exp__io_in  [6:2])) ? {8'h0,  core__ibuf__exp__io_in  [11:7],7'h33}:{  core__ibuf__exp__io_in  [11:7],(|(  core__ibuf__exp__io_in  [11:7])) ? 15'h67:15'h1F}}}:  core__ibuf__exp___io_out_T_39   ? {3'h0,  core__ibuf__exp__io_in  [4:2],  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:5],11'h13,  core__ibuf__exp__io_in  [11:7],  core__ibuf__exp__io_out_s_load_opc  }:  core__ibuf__exp___io_out_T_37   ? {4'h0,  core__ibuf__exp__io_in  [3:2],  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:4],10'h12,  core__ibuf__exp__io_in  [11:7],  core__ibuf__exp__io_out_s_load_opc  }:  core__ibuf__exp___io_out_T_35   ? {3'h0,  core__ibuf__exp__io_in  [4:2],  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:5],11'h13,  core__ibuf__exp__io_in  [11:7],7'h7}:  core__ibuf__exp___io_out_T_33   ? {6'h0,  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:2],  core__ibuf__exp__io_in  [11:7],3'h1,  core__ibuf__exp__io_in  [11:7],7'h13}:  core__ibuf__exp___io_out_T_31   ? {  core__ibuf__exp___GEN  ,  core__ibuf__exp__io_in  [6:5],  core__ibuf__exp__io_in  [2],7'h1,  core__ibuf__exp__io_in  [9:7],3'h1,  core__ibuf__exp__io_in  [11:10],  core__ibuf__exp__io_in  [4:3],  core__ibuf__exp__io_in  [12],7'h63}:  core__ibuf__exp___io_out_T_29   ? {  core__ibuf__exp___GEN  ,  core__ibuf__exp__io_in  [6:5],  core__ibuf__exp__io_in  [2],7'h1,  core__ibuf__exp__io_in  [9:7],3'h0,  core__ibuf__exp__io_in  [11:10],  core__ibuf__exp__io_in  [4:3],  core__ibuf__exp__io_in  [12],7'h63}:  core__ibuf__exp___io_out_T_2  ==5'hD ? {  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [8],  core__ibuf__exp__io_in  [10:9],  core__ibuf__exp__io_in  [6],  core__ibuf__exp__io_in  [7],  core__ibuf__exp__io_in  [2],  core__ibuf__exp__io_in  [11],  core__ibuf__exp__io_in  [5:3],{9{  core__ibuf__exp__io_in  [12]}},12'h6F}:  core__ibuf__exp___io_out_T_2  ==5'hC ? ((&(  core__ibuf__exp__io_in  [11:10])) ? {1'h0,  core__ibuf__exp__io_in  [6:5]==2'h0,7'h1,  core__ibuf__exp__io_in  [4:2],2'h1,  core__ibuf__exp__io_in  [9:7],  core__ibuf__exp__casez_tmp  ,2'h1,  core__ibuf__exp__io_in  [9:7],3'h3,  core__ibuf__exp__io_in  [12],3'h3}:{  core__ibuf__exp__io_in  [11:10]==2'h2 ? {{7{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [6:2],2'h1,  core__ibuf__exp__io_in  [9:7],5'h1D}:{1'h0,  core__ibuf__exp__io_in  [11:10]==2'h1,4'h0,  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:2],2'h1,  core__ibuf__exp__io_in  [9:7],5'h15},  core__ibuf__exp__io_in  [9:7],7'h13}):  core__ibuf__exp___io_out_T_2  ==5'hB ? {{3{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [11:7]==5'h0|  core__ibuf__exp__io_in  [11:7]==5'h2 ? {  core__ibuf__exp__io_in  [4:3],  core__ibuf__exp__io_in  [5],  core__ibuf__exp__io_in  [2],  core__ibuf__exp__io_in  [6],4'h0,  core__ibuf__exp__io_in  [11:7],3'h0,  core__ibuf__exp__io_in  [11:7],(|{{7{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [6:2]}) ? 7'h13:7'h1F}:{{12{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [6:2],  core__ibuf__exp__io_in  [11:7],3'h3,{{7{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [6:2]}==12'h0,3'h7}}:  core__ibuf__exp___io_out_T_2  ==5'hA ? {{7{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [6:2],8'h0,  core__ibuf__exp__io_in  [11:7],7'h13}:  core__ibuf__exp___io_out_T_2  ==5'h9 ? {{7{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [6:2],  core__ibuf__exp__io_in  [11:7],3'h0,  core__ibuf__exp__io_in  [11:7],4'h3,  core__ibuf__exp__io_in  [11:7]==5'h0,2'h3}:  core__ibuf__exp___io_out_T_2  ==5'h8 ? {{7{  core__ibuf__exp__io_in  [12]}},  core__ibuf__exp__io_in  [6:2],  core__ibuf__exp__io_in  [11:7],3'h0,  core__ibuf__exp__io_in  [11:7],7'h13}:  core__ibuf__exp___io_out_T_2  ==5'h7 ? {4'h0,  core__ibuf__exp__io_in  [6:5],  core__ibuf__exp__io_in  [12],2'h1,  core__ibuf__exp__io_in  [4:2],2'h1,  core__ibuf__exp__io_in  [9:7],3'h3,  core__ibuf__exp__io_in  [11:10],10'h23}:  core__ibuf__exp___io_out_T_2  ==5'h6 ? {5'h0,  core__ibuf__exp__io_in  [5],  core__ibuf__exp__io_in  [12],2'h1,  core__ibuf__exp__io_in  [4:2],2'h1,  core__ibuf__exp__io_in  [9:7],3'h2,  core__ibuf__exp__io_in  [11:10],  core__ibuf__exp__io_in  [6],9'h23}:  core__ibuf__exp___io_out_T_2  ==5'h5 ? {4'h0,  core__ibuf__exp__io_in  [6:5],  core__ibuf__exp__io_in  [12],2'h1,  core__ibuf__exp__io_in  [4:2],2'h1,  core__ibuf__exp__io_in  [9:7],3'h3,  core__ibuf__exp__io_in  [11:10],10'h27}:  core__ibuf__exp___io_out_T_2  ==5'h4 ? {5'h0,  core__ibuf__exp__io_in  [5],  core__ibuf__exp__io_in  [12],2'h1,  core__ibuf__exp__io_in  [4:2],2'h1,  core__ibuf__exp__io_in  [9:7],3'h2,  core__ibuf__exp__io_in  [11:10],  core__ibuf__exp__io_in  [6],9'h3F}:  core__ibuf__exp___io_out_T_2  ==5'h3 ? {4'h0,  core__ibuf__exp__io_in  [6:5],  core__ibuf__exp__io_in  [12:10],5'h1,  core__ibuf__exp__io_in  [9:7],5'hD,  core__ibuf__exp__io_in  [4:2],7'h3}:  core__ibuf__exp___io_out_T_2  ==5'h2 ? {5'h0,  core__ibuf__exp__io_in  [5],  core__ibuf__exp__io_in  [12:10],  core__ibuf__exp__io_in  [6],4'h1,  core__ibuf__exp__io_in  [9:7],5'h9,  core__ibuf__exp__io_in  [4:2],7'h3}:  core__ibuf__exp___io_out_T_2  ==5'h1 ? {4'h0,  core__ibuf__exp__io_in  [6:5],  core__ibuf__exp__io_in  [12:10],5'h1,  core__ibuf__exp__io_in  [9:7],5'hD,  core__ibuf__exp__io_in  [4:2],7'h7}:{2'h0,  core__ibuf__exp__io_in  [10:7],  core__ibuf__exp__io_in  [12:11],  core__ibuf__exp__io_in  [5],  core__ibuf__exp__io_in  [6],12'h41,  core__ibuf__exp__io_in  [4:2],(|(  core__ibuf__exp__io_in  [12:5])) ? 7'h13:7'h1F}; 
   wire  core__ibuf__exp___io_out_T_43  =  core__ibuf__exp___io_out_T_2  ==5'h15; 
   wire  core__ibuf__exp___io_out_T_45  =  core__ibuf__exp___io_out_T_2  ==5'h16; 
   wire  core__ibuf__exp___io_out_T_47  =  core__ibuf__exp___io_out_T_2  ==5'h17; 
   wire  core__ibuf__exp___io_out_T_49  =  core__ibuf__exp___io_out_T_2  ==5'h18; 
   wire  core__ibuf__exp___io_out_T_51  =  core__ibuf__exp___io_out_T_2  ==5'h19; 
   wire  core__ibuf__exp___io_out_T_53  =  core__ibuf__exp___io_out_T_2  ==5'h1A; 
   wire  core__ibuf__exp___io_out_T_55  =  core__ibuf__exp___io_out_T_2  ==5'h1B; 
   wire  core__ibuf__exp___io_out_T_57  =  core__ibuf__exp___io_out_T_2  ==5'h1C; 
   wire  core__ibuf__exp___io_out_T_59  =  core__ibuf__exp___io_out_T_2  ==5'h1D; 
   wire  core__ibuf__exp___io_out_T_61  =  core__ibuf__exp___io_out_T_2  ==5'h1E; 
   reg[4:0]  core__ibuf__exp__casez_tmp_0  ; 
   wire[4:0]  core__ibuf__exp__io_out_s_7_rd  ={2'h1,  core__ibuf__exp__io_in  [4:2]}; 
  always @(*)
       begin 
         casez (  core__ibuf__exp___io_out_T_2  )
          5 'b00000: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b00001: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b00010: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b00011: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b00100: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b00101: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b00110: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b00111: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_out_s_7_rd  ;
          5 'b01000: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b01001: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b01010: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b01011: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b01100: 
              core__ibuf__exp__casez_tmp_0   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b01101: 
              core__ibuf__exp__casez_tmp_0   =5'h0;
          5 'b01110: 
              core__ibuf__exp__casez_tmp_0   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b01111: 
              core__ibuf__exp__casez_tmp_0   =5'h0;
          5 'b10000: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b10001: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b10010: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b10011: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b10100: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [12] ? ((|(  core__ibuf__exp__io_in  [6:2])) ?   core__ibuf__exp__io_in  [11:7]:5'h1):(|(  core__ibuf__exp__io_in  [6:2])) ?   core__ibuf__exp__io_in  [11:7]:5'h0;
          5 'b10101: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b10110: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b10111: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b11000: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b11001: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b11010: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b11011: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b11100: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b11101: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          5 'b11110: 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
          default : 
              core__ibuf__exp__casez_tmp_0   =  core__ibuf__exp__io_in  [11:7];
         endcase 
       end
  
   reg[4:0]  core__ibuf__exp__casez_tmp_1  ; 
  always @(*)
       begin 
         casez (  core__ibuf__exp___io_out_T_2  )
          5 'b00000: 
              core__ibuf__exp__casez_tmp_1   =5'h2;
          5 'b00001: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b00010: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b00011: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b00100: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b00101: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b00110: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b00111: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b01000: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [11:7];
          5 'b01001: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [11:7];
          5 'b01010: 
              core__ibuf__exp__casez_tmp_1   =5'h0;
          5 'b01011: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [11:7];
          5 'b01100: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b01101: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b01110: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b01111: 
              core__ibuf__exp__casez_tmp_1   ={2'h1,  core__ibuf__exp__io_in  [9:7]};
          5 'b10000: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [11:7];
          5 'b10001: 
              core__ibuf__exp__casez_tmp_1   =5'h2;
          5 'b10010: 
              core__ibuf__exp__casez_tmp_1   =5'h2;
          5 'b10011: 
              core__ibuf__exp__casez_tmp_1   =5'h2;
          5 'b10100: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [12]|~(|(  core__ibuf__exp__io_in  [6:2])) ?   core__ibuf__exp__io_in  [11:7]:5'h0;
          5 'b10101: 
              core__ibuf__exp__casez_tmp_1   =5'h2;
          5 'b10110: 
              core__ibuf__exp__casez_tmp_1   =5'h2;
          5 'b10111: 
              core__ibuf__exp__casez_tmp_1   =5'h2;
          5 'b11000: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
          5 'b11001: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
          5 'b11010: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
          5 'b11011: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
          5 'b11100: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
          5 'b11101: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
          5 'b11110: 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
          default : 
              core__ibuf__exp__casez_tmp_1   =  core__ibuf__exp__io_in  [19:15];
         endcase 
       end
  
  assign   core__ibuf__exp__io_out_bits  =(&  core__ibuf__exp___io_out_T_2  )|  core__ibuf__exp___io_out_T_61  |  core__ibuf__exp___io_out_T_59  |  core__ibuf__exp___io_out_T_57  |  core__ibuf__exp___io_out_T_55  |  core__ibuf__exp___io_out_T_53  |  core__ibuf__exp___io_out_T_51  |  core__ibuf__exp___io_out_T_49   ?   core__ibuf__exp__io_in  :  core__ibuf__exp___io_out_T_47   ? {3'h0,  core__ibuf__exp__io_in  [9:7],  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:2],8'h13,  core__ibuf__exp__io_in  [11:10],10'h23}:  core__ibuf__exp___io_out_T_45   ? {4'h0,  core__ibuf__exp__io_in  [8:7],  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:2],8'h12,  core__ibuf__exp__io_in  [11:9],9'h23}:  core__ibuf__exp___io_out_T_43   ? {3'h0,  core__ibuf__exp__io_in  [9:7],  core__ibuf__exp__io_in  [12],  core__ibuf__exp__io_in  [6:2],8'h13,  core__ibuf__exp__io_in  [11:10],10'h27}:  core__ibuf__exp___io_out_T_42_bits  ; 
  assign   core__ibuf__exp__io_out_rd  =  core__ibuf__exp__casez_tmp_0  ; 
  assign   core__ibuf__exp__io_out_rs1  =  core__ibuf__exp__casez_tmp_1  ; 
  assign   core__ibuf__exp__io_out_rs2  =(&  core__ibuf__exp___io_out_T_2  )|  core__ibuf__exp___io_out_T_61  |  core__ibuf__exp___io_out_T_59  |  core__ibuf__exp___io_out_T_57  |  core__ibuf__exp___io_out_T_55  |  core__ibuf__exp___io_out_T_53  |  core__ibuf__exp___io_out_T_51  |  core__ibuf__exp___io_out_T_49   ?   core__ibuf__exp__io_in  [24:20]:  core__ibuf__exp___io_out_T_47  |  core__ibuf__exp___io_out_T_45  |  core__ibuf__exp___io_out_T_43  |  core__ibuf__exp___io_out_T_41  |  core__ibuf__exp___io_out_T_39  |  core__ibuf__exp___io_out_T_37  |  core__ibuf__exp___io_out_T_35  |  core__ibuf__exp___io_out_T_33   ?   core__ibuf__exp__io_in  [6:2]:  core__ibuf__exp___io_out_T_31  |  core__ibuf__exp___io_out_T_29   ? 5'h0:{2'h1,  core__ibuf__exp__io_in  [4:2]}; 
  assign   core__ibuf__exp__io_rvc  =  core__ibuf__exp__io_in  [1:0]!=2'h3;
assign core__ibuf__exp__io_in = core__ibuf__inst;
assign core__ibuf__io_inst_0_bits_inst_bits = core__ibuf__exp__io_out_bits;
assign core__ibuf__io_inst_0_bits_inst_rd = core__ibuf__exp__io_out_rd;
assign core__ibuf__io_inst_0_bits_inst_rs1 = core__ibuf__exp__io_out_rs1;
assign core__ibuf__io_inst_0_bits_inst_rs2 = core__ibuf__exp__io_out_rs2;
assign core__ibuf___exp_io_rvc = core__ibuf__exp__io_rvc;
 
  assign   core__ibuf__io_imem_ready  =  core__ibuf__io_inst_0_ready  &  core__ibuf___nBufValid_T  &(  core__ibuf___nICReady_T  >=  core__ibuf___nIC_T_2  |~(  core__ibuf___nBufValid_T_6  [1])); 
  assign   core__ibuf__io_pc  =  core__ibuf__nBufValid   ?   core__ibuf__buf_pc  :  core__ibuf__io_imem_bits_pc  ; 
  assign   core__ibuf__io_inst_0_valid  =  core__ibuf___valid_T_1  [0]&  core__ibuf__full_insn  ; 
  assign   core__ibuf__io_inst_0_bits_xcpt0_pf_inst  =  core__ibuf___bufMask_T_1  [0] ?   core__ibuf__buf_xcpt_pf_inst  :  core__ibuf__io_imem_bits_xcpt_pf_inst  ; 
  assign   core__ibuf__io_inst_0_bits_xcpt0_gf_inst  =  core__ibuf___bufMask_T_1  [0] ?   core__ibuf__buf_xcpt_gf_inst  :  core__ibuf__io_imem_bits_xcpt_gf_inst  ; 
  assign   core__ibuf__io_inst_0_bits_xcpt0_ae_inst  =  core__ibuf___bufMask_T_1  [0] ?   core__ibuf__buf_xcpt_ae_inst  :  core__ibuf__io_imem_bits_xcpt_ae_inst  ; 
  assign   core__ibuf__io_inst_0_bits_xcpt1_pf_inst  =  core__ibuf___io_inst_0_bits_xcpt1_T_5  [2]; 
  assign   core__ibuf__io_inst_0_bits_xcpt1_gf_inst  =  core__ibuf___io_inst_0_bits_xcpt1_T_5  [1]; 
  assign   core__ibuf__io_inst_0_bits_xcpt1_ae_inst  =  core__ibuf___io_inst_0_bits_xcpt1_T_5  [0]; 
  assign   core__ibuf__io_inst_0_bits_replay  =  core__ibuf__ic_replay  [0]|~  core__ibuf___exp_io_rvc  &  core__ibuf__ic_replay  [1]; 
  assign   core__ibuf__io_inst_0_bits_rvc  =  core__ibuf___exp_io_rvc  ; 
  assign   core__ibuf__io_inst_0_bits_raw  =  core__ibuf__inst  ;
assign core__ibuf__clock = core__clock;
assign core__ibuf__reset = core__reset;
assign core__io_imem_resp_ready = core__ibuf__io_imem_ready;
assign core__ibuf__io_imem_valid = core__io_imem_resp_valid;
assign core__ibuf__io_imem_bits_pc = core__io_imem_resp_bits_pc;
assign core__ibuf__io_imem_bits_data = core__io_imem_resp_bits_data;
assign core__ibuf__io_imem_bits_xcpt_pf_inst = core__io_imem_resp_bits_xcpt_pf_inst;
assign core__ibuf__io_imem_bits_xcpt_gf_inst = core__io_imem_resp_bits_xcpt_gf_inst;
assign core__ibuf__io_imem_bits_xcpt_ae_inst = core__io_imem_resp_bits_xcpt_ae_inst;
assign core__ibuf__io_imem_bits_replay = core__io_imem_resp_bits_replay;
assign core__ibuf__io_kill = core__ibuf_io_kill;
assign core___ibuf_io_pc = core__ibuf__io_pc;
assign core__ibuf__io_inst_0_ready = ~core___ctrl_stalld_T_28;
assign core___ibuf_io_inst_0_valid = core__ibuf__io_inst_0_valid;
assign core___ibuf_io_inst_0_bits_xcpt0_pf_inst = core__ibuf__io_inst_0_bits_xcpt0_pf_inst;
assign core___ibuf_io_inst_0_bits_xcpt0_gf_inst = core__ibuf__io_inst_0_bits_xcpt0_gf_inst;
assign core___ibuf_io_inst_0_bits_xcpt0_ae_inst = core__ibuf__io_inst_0_bits_xcpt0_ae_inst;
assign core___ibuf_io_inst_0_bits_xcpt1_pf_inst = core__ibuf__io_inst_0_bits_xcpt1_pf_inst;
assign core___ibuf_io_inst_0_bits_xcpt1_gf_inst = core__ibuf__io_inst_0_bits_xcpt1_gf_inst;
assign core___ibuf_io_inst_0_bits_xcpt1_ae_inst = core__ibuf__io_inst_0_bits_xcpt1_ae_inst;
assign core___ibuf_io_inst_0_bits_replay = core__ibuf__io_inst_0_bits_replay;
assign core___ibuf_io_inst_0_bits_rvc = core__ibuf__io_inst_0_bits_rvc;
assign core___ibuf_io_inst_0_bits_inst_bits = core__ibuf__io_inst_0_bits_inst_bits;
assign core___ibuf_io_inst_0_bits_inst_rd = core__ibuf__io_inst_0_bits_inst_rd;
assign core___ibuf_io_inst_0_bits_inst_rs1 = core__ibuf__io_inst_0_bits_inst_rs1;
assign core___ibuf_io_inst_0_bits_inst_rs2 = core__ibuf__io_inst_0_bits_inst_rs2;
assign core___ibuf_io_inst_0_bits_raw = core__ibuf__io_inst_0_bits_raw;
  
  rf_31x64    core__rf_ext  (. R0_addr (~  core___ibuf_io_inst_0_bits_inst_rs2  ),. R0_en (1'h1),. R0_clk (  core__clock  ),. R0_data (  core___rf_ext_R0_data  ),. R1_addr (~  core___ibuf_io_inst_0_bits_inst_rs1  ),. R1_en (1'h1),. R1_clk (  core__clock  ),. R1_data (  core___rf_ext_R1_data  ),. W0_addr (~  core__rf_waddr  ),. W0_en (  core__rf_wen  &(|  core__rf_waddr  )),. W0_clk (  core__clock  ),. W0_data (  core__rf_wdata  ));  
  CSRFile    core__csr  (. clock (  core__clock  ),. reset (  core__reset  ),. io_ungated_clock (  core__clock  ),. io_interrupts_debug (  core__io_interrupts_debug  ),. io_interrupts_mtip (  core__io_interrupts_mtip  ),. io_interrupts_msip (  core__io_interrupts_msip  ),. io_interrupts_meip (  core__io_interrupts_meip  ),. io_hartid (  core__io_hartid  ),. io_rw_addr (  core__wb_reg_inst  [31:20]),. io_rw_cmd (  core__wb_ctrl_csr  &{  core__wb_reg_valid  ,2'h3}),. io_rw_rdata (  core___csr_io_rw_rdata  ),. io_rw_wdata (  core__wb_reg_wdata  ),. io_decode_0_inst (  core___ibuf_io_inst_0_bits_inst_bits  ),. io_decode_0_read_illegal (  core___csr_io_decode_0_read_illegal  ),. io_decode_0_write_illegal (  core___csr_io_decode_0_write_illegal  ),. io_decode_0_write_flush (  core___csr_io_decode_0_write_flush  ),. io_decode_0_system_illegal (  core___csr_io_decode_0_system_illegal  ),. io_decode_0_virtual_access_illegal (  core___csr_io_decode_0_virtual_access_illegal  ),. io_decode_0_virtual_system_illegal (  core___csr_io_decode_0_virtual_system_illegal  ),. io_csr_stall (  core___csr_io_csr_stall  ),. io_eret (  core___csr_io_eret  ),. io_singleStep (  core___csr_io_singleStep  ),. io_status_debug (  core___csr_io_status_debug  ),. io_status_wfi (  core__io_wfi  ),. io_status_isa (  core___csr_io_status_isa  ),. io_status_dv (  core___csr_io_status_dv  ),. io_status_v (  core___csr_io_status_v  ),. io_evec (  core___csr_io_evec  ),. io_exception (  core__wb_xcpt  ),. io_retire (  core__wb_valid  ),. io_cause (  core__wb_reg_xcpt   ?   core__wb_reg_cause  :{59'h0,  core___GEN_0   ? 5'hF:  core___GEN_1   ? 5'hD:{2'h0,  core___GEN_2   ? 3'h7:  core___GEN_3   ? 3'h5:{1'h1,  core___GEN_4  ,1'h0}}}),. io_pc (  core__wb_reg_pc  ),. io_tval (  core__wb_xcpt  &(  core__tval_any_addr  |  core__wb_reg_cause  ==64'h2) ? {  core__wb_reg_wdata  [63:33]==31'h0|(&(  core__wb_reg_wdata  [63:33])) ?   core__wb_reg_wdata  [33]:~(  core__wb_reg_wdata  [32]),  core__wb_reg_wdata  [32:0]}:34'h0),. io_gva (  core__wb_xcpt  &(  core__tval_any_addr  &  core___csr_io_status_v  |~  core__wb_reg_xcpt  &  core__wb_reg_hls_or_dv  )),. io_time (  core___csr_io_time  ),. io_interrupt (  core___csr_io_interrupt  ),. io_interrupt_cause (  core___csr_io_interrupt_cause  ),. io_bp_0_control_action (  core___csr_io_bp_0_control_action  ),. io_bp_0_control_tmatch (  core___csr_io_bp_0_control_tmatch  ),. io_bp_0_control_x (  core___csr_io_bp_0_control_x  ),. io_bp_0_control_w (  core___csr_io_bp_0_control_w  ),. io_bp_0_control_r (  core___csr_io_bp_0_control_r  ),. io_bp_0_address (  core___csr_io_bp_0_address  ),. io_pmp_cfg_l_0 (  core__io_ptw_pmp_cfg_l_0  ),. io_pmp_cfg_l_1 (  core__io_ptw_pmp_cfg_l_1  ),. io_pmp_cfg_l_2 (  core__io_ptw_pmp_cfg_l_2  ),. io_pmp_cfg_l_3 (  core__io_ptw_pmp_cfg_l_3  ),. io_pmp_cfg_l_4 (  core__io_ptw_pmp_cfg_l_4  ),. io_pmp_cfg_l_5 (  core__io_ptw_pmp_cfg_l_5  ),. io_pmp_cfg_l_6 (  core__io_ptw_pmp_cfg_l_6  ),. io_pmp_cfg_l_7 (  core__io_ptw_pmp_cfg_l_7  ),. io_pmp_cfg_a_0 (  core__io_ptw_pmp_cfg_a_0  ),. io_pmp_cfg_a_1 (  core__io_ptw_pmp_cfg_a_1  ),. io_pmp_cfg_a_2 (  core__io_ptw_pmp_cfg_a_2  ),. io_pmp_cfg_a_3 (  core__io_ptw_pmp_cfg_a_3  ),. io_pmp_cfg_a_4 (  core__io_ptw_pmp_cfg_a_4  ),. io_pmp_cfg_a_5 (  core__io_ptw_pmp_cfg_a_5  ),. io_pmp_cfg_a_6 (  core__io_ptw_pmp_cfg_a_6  ),. io_pmp_cfg_a_7 (  core__io_ptw_pmp_cfg_a_7  ),. io_pmp_cfg_x_0 (  core__io_ptw_pmp_cfg_x_0  ),. io_pmp_cfg_x_1 (  core__io_ptw_pmp_cfg_x_1  ),. io_pmp_cfg_x_2 (  core__io_ptw_pmp_cfg_x_2  ),. io_pmp_cfg_x_3 (  core__io_ptw_pmp_cfg_x_3  ),. io_pmp_cfg_x_4 (  core__io_ptw_pmp_cfg_x_4  ),. io_pmp_cfg_x_5 (  core__io_ptw_pmp_cfg_x_5  ),. io_pmp_cfg_x_6 (  core__io_ptw_pmp_cfg_x_6  ),. io_pmp_cfg_x_7 (  core__io_ptw_pmp_cfg_x_7  ),. io_pmp_cfg_w_0 (  core__io_ptw_pmp_cfg_w_0  ),. io_pmp_cfg_w_1 (  core__io_ptw_pmp_cfg_w_1  ),. io_pmp_cfg_w_2 (  core__io_ptw_pmp_cfg_w_2  ),. io_pmp_cfg_w_3 (  core__io_ptw_pmp_cfg_w_3  ),. io_pmp_cfg_w_4 (  core__io_ptw_pmp_cfg_w_4  ),. io_pmp_cfg_w_5 (  core__io_ptw_pmp_cfg_w_5  ),. io_pmp_cfg_w_6 (  core__io_ptw_pmp_cfg_w_6  ),. io_pmp_cfg_w_7 (  core__io_ptw_pmp_cfg_w_7  ),. io_pmp_cfg_r_0 (  core__io_ptw_pmp_cfg_r_0  ),. io_pmp_cfg_r_1 (  core__io_ptw_pmp_cfg_r_1  ),. io_pmp_cfg_r_2 (  core__io_ptw_pmp_cfg_r_2  ),. io_pmp_cfg_r_3 (  core__io_ptw_pmp_cfg_r_3  ),. io_pmp_cfg_r_4 (  core__io_ptw_pmp_cfg_r_4  ),. io_pmp_cfg_r_5 (  core__io_ptw_pmp_cfg_r_5  ),. io_pmp_cfg_r_6 (  core__io_ptw_pmp_cfg_r_6  ),. io_pmp_cfg_r_7 (  core__io_ptw_pmp_cfg_r_7  ),. io_pmp_addr_0 (  core__io_ptw_pmp_addr_0  ),. io_pmp_addr_1 (  core__io_ptw_pmp_addr_1  ),. io_pmp_addr_2 (  core__io_ptw_pmp_addr_2  ),. io_pmp_addr_3 (  core__io_ptw_pmp_addr_3  ),. io_pmp_addr_4 (  core__io_ptw_pmp_addr_4  ),. io_pmp_addr_5 (  core__io_ptw_pmp_addr_5  ),. io_pmp_addr_6 (  core__io_ptw_pmp_addr_6  ),. io_pmp_addr_7 (  core__io_ptw_pmp_addr_7  ),. io_pmp_mask_0 (  core__io_ptw_pmp_mask_0  ),. io_pmp_mask_1 (  core__io_ptw_pmp_mask_1  ),. io_pmp_mask_2 (  core__io_ptw_pmp_mask_2  ),. io_pmp_mask_3 (  core__io_ptw_pmp_mask_3  ),. io_pmp_mask_4 (  core__io_ptw_pmp_mask_4  ),. io_pmp_mask_5 (  core__io_ptw_pmp_mask_5  ),. io_pmp_mask_6 (  core__io_ptw_pmp_mask_6  ),. io_pmp_mask_7 (  core__io_ptw_pmp_mask_7  ),. io_inhibit_cycle (  core___csr_io_inhibit_cycle  ),. io_inst_0 ({(&(  core__wb_reg_raw_inst  [1:0])) ?   core__wb_reg_inst  [31:16]:16'h0,  core__wb_reg_raw_inst  [15:0]}),. io_trace_valid_0 (  core___csr_io_trace_valid_0  ),. io_trace_iaddr_0 (  core___csr_io_trace_iaddr_0  ),. io_trace_insn_0 (  core___csr_io_trace_insn_0  ),. io_trace_exception_0 (  core___csr_io_trace_exception_0  ),. io_customCSRs_0_value (  core___csr_io_customCSRs_0_value  ));  
  BreakpointUnit    core__bpu  (. io_status_debug (  core___csr_io_status_debug  ),. io_bp_0_control_action (  core___csr_io_bp_0_control_action  ),. io_bp_0_control_tmatch (  core___csr_io_bp_0_control_tmatch  ),. io_bp_0_control_x (  core___csr_io_bp_0_control_x  ),. io_bp_0_control_w (  core___csr_io_bp_0_control_w  ),. io_bp_0_control_r (  core___csr_io_bp_0_control_r  ),. io_bp_0_address (  core___csr_io_bp_0_address  ),. io_pc (  core___ibuf_io_pc  [32:0]),. io_ea (  core__mem_reg_wdata  [32:0]),. io_xcpt_if (  core___bpu_io_xcpt_if  ),. io_xcpt_ld (  core___bpu_io_xcpt_ld  ),. io_xcpt_st (  core___bpu_io_xcpt_st  ),. io_debug_if (  core___bpu_io_debug_if  ),. io_debug_ld (  core___bpu_io_debug_ld  ),. io_debug_st (  core___bpu_io_debug_st  ));  
  ALU    core__alu  (. io_dw (  core__ex_ctrl_alu_dw  ),. io_fn (  core__ex_ctrl_alu_fn  ),. io_in2 (  core__casez_tmp_1  ),. io_in1 (  core__ex_ctrl_sel_alu1  ==2'h2 ? {{30{  core__ex_reg_pc  [33]}},  core__ex_reg_pc  }:  core__ex_ctrl_sel_alu1  ==2'h1 ?   core__ex_rs_0  :64'h0),. io_out (  core___alu_io_out  ),. io_adder_out (  core___alu_io_adder_out  ),. io_cmp_out (  core___alu_io_cmp_out  ));  
  MulDiv    core__div  (. clock (  core__clock  ),. reset (  core__reset  ),. io_req_ready (  core___div_io_req_ready  ),. io_req_valid (  core__div_io_req_valid  ),. io_req_bits_fn (  core__ex_ctrl_alu_fn  ),. io_req_bits_dw (  core__ex_ctrl_alu_dw  ),. io_req_bits_in1 (  core__ex_rs_0  ),. io_req_bits_in2 (  core__ex_rs_1  ),. io_req_bits_tag (  core__ex_reg_inst  [11:7]),. io_kill (  core__killm_common  &  core__div_io_kill_REG  ),. io_resp_ready (  core__div_io_resp_ready  ),. io_resp_valid (  core___div_io_resp_valid  ),. io_resp_bits_data (  core___div_io_resp_bits_data  ),. io_resp_bits_tag (  core___div_io_resp_bits_tag  ));  
  PlusArgTimeout    core__PlusArgTimeout  (. clock (  core__clock  ),. reset (  core__reset  ),. io_count (  core___csr_io_time  [31:0])); 
  assign   core__io_imem_might_request  =  core__imem_might_request_reg  ; 
  assign   core__io_imem_req_valid  =  core__ibuf_io_kill  ; 
  assign   core__io_imem_req_bits_pc  =  core__wb_xcpt  |  core___csr_io_eret   ?   core___csr_io_evec  :  core___replay_wb_T   ?   core__wb_reg_pc  :  core__mem_npc  ; 
  assign   core__io_imem_req_bits_speculative  =~  core__take_pc_wb  ; 
  assign   core__io_imem_btb_update_valid  =  core__mem_reg_valid  &~  core__take_pc_wb  &(  core__ex_pc_valid   ?   core__mem_npc  !=  core__ex_reg_pc  :~(  core___ibuf_io_inst_0_valid  |  core__io_imem_resp_valid  )|  core__mem_npc  !=  core___ibuf_io_pc  )&(~(  core__mem_ctrl_branch  |  core__mem_ctrl_jalr  |  core__mem_ctrl_jal  )|  core__mem_cfi_taken  ); 
  assign   core__io_imem_bht_update_valid  =  core__mem_reg_valid  &~  core__take_pc_wb  ; 
  assign   core__io_imem_flush_icache  =  core__wb_reg_valid  &  core__wb_ctrl_fence_i  &~  core__io_dmem_s2_nack  ; 
  assign   core__io_dmem_req_valid  =  core__io_dmem_req_valid_0  ; 
  assign   core__io_dmem_req_bits_addr  ={  core__ex_rs_0  [63:33]==31'h0|(&(  core__ex_rs_0  [63:33])) ?   core___alu_io_adder_out  [33]:~(  core___alu_io_adder_out  [32]),  core___alu_io_adder_out  [32:0]}; 
  assign   core__io_dmem_req_bits_tag  ={  core__ex_reg_inst  [11:7],  core__ex_ctrl_fp  }; 
  assign   core__io_dmem_req_bits_cmd  =  core__ex_ctrl_mem_cmd  ; 
  assign   core__io_dmem_req_bits_size  =  core__ex_reg_mem_size  ; 
  assign   core__io_dmem_req_bits_signed  =~(  core__ex_reg_inst  [14]); 
  assign   core__io_dmem_req_bits_dv  =  core___csr_io_status_dv  ; 
  assign   core__io_dmem_s1_kill  =  core__killm_common  |  core__mem_ldst_xcpt  ; 
  assign   core__io_dmem_s1_data_data  =  core__mem_reg_rs2  ; 
  assign   core__io_ptw_status_debug  =  core___csr_io_status_debug  ; 
  assign   core__io_ptw_customCSRs_csrs_0_value  =  core___csr_io_customCSRs_0_value  ;
assign core__clock = clock;
assign core__reset = reset;
assign core__io_hartid = auto_hartid_in;
assign core__io_interrupts_debug = _intXbar_auto_int_out_0;
assign core__io_interrupts_mtip = _intXbar_auto_int_out_2;
assign core__io_interrupts_msip = _intXbar_auto_int_out_1;
assign core__io_interrupts_meip = _intXbar_auto_int_out_3;
assign _core_io_imem_might_request = core__io_imem_might_request;
assign _core_io_imem_req_valid = core__io_imem_req_valid;
assign _core_io_imem_req_bits_pc = core__io_imem_req_bits_pc;
assign _core_io_imem_req_bits_speculative = core__io_imem_req_bits_speculative;
assign _core_io_imem_resp_ready = core__io_imem_resp_ready;
assign core__io_imem_resp_valid = _frontend_io_cpu_resp_valid;
assign core__io_imem_resp_bits_pc = _frontend_io_cpu_resp_bits_pc;
assign core__io_imem_resp_bits_data = _frontend_io_cpu_resp_bits_data;
assign core__io_imem_resp_bits_xcpt_pf_inst = _frontend_io_cpu_resp_bits_xcpt_pf_inst;
assign core__io_imem_resp_bits_xcpt_gf_inst = _frontend_io_cpu_resp_bits_xcpt_gf_inst;
assign core__io_imem_resp_bits_xcpt_ae_inst = _frontend_io_cpu_resp_bits_xcpt_ae_inst;
assign core__io_imem_resp_bits_replay = _frontend_io_cpu_resp_bits_replay;
assign _core_io_imem_btb_update_valid = core__io_imem_btb_update_valid;
assign _core_io_imem_bht_update_valid = core__io_imem_bht_update_valid;
assign _core_io_imem_flush_icache = core__io_imem_flush_icache;
assign core__io_dmem_req_ready = _dcacheArb_io_requestor_0_req_ready;
assign _core_io_dmem_req_valid = core__io_dmem_req_valid;
assign _core_io_dmem_req_bits_addr = core__io_dmem_req_bits_addr;
assign _core_io_dmem_req_bits_tag = core__io_dmem_req_bits_tag;
assign _core_io_dmem_req_bits_cmd = core__io_dmem_req_bits_cmd;
assign _core_io_dmem_req_bits_size = core__io_dmem_req_bits_size;
assign _core_io_dmem_req_bits_signed = core__io_dmem_req_bits_signed;
assign _core_io_dmem_req_bits_dv = core__io_dmem_req_bits_dv;
assign _core_io_dmem_s1_kill = core__io_dmem_s1_kill;
assign _core_io_dmem_s1_data_data = core__io_dmem_s1_data_data;
assign core__io_dmem_s2_nack = _dcacheArb_io_requestor_0_s2_nack;
assign core__io_dmem_resp_valid = _dcacheArb_io_requestor_0_resp_valid;
assign core__io_dmem_resp_bits_tag = _dcacheArb_io_requestor_0_resp_bits_tag;
assign core__io_dmem_resp_bits_data = _dcacheArb_io_requestor_0_resp_bits_data;
assign core__io_dmem_resp_bits_replay = _dcacheArb_io_requestor_0_resp_bits_replay;
assign core__io_dmem_resp_bits_has_data = _dcacheArb_io_requestor_0_resp_bits_has_data;
assign core__io_dmem_resp_bits_data_word_bypass = _dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
assign core__io_dmem_replay_next = _dcacheArb_io_requestor_0_replay_next;
assign core__io_dmem_s2_xcpt_ma_ld = _dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
assign core__io_dmem_s2_xcpt_ma_st = _dcacheArb_io_requestor_0_s2_xcpt_ma_st;
assign core__io_dmem_s2_xcpt_pf_ld = _dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
assign core__io_dmem_s2_xcpt_pf_st = _dcacheArb_io_requestor_0_s2_xcpt_pf_st;
assign core__io_dmem_s2_xcpt_ae_ld = _dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
assign core__io_dmem_s2_xcpt_ae_st = _dcacheArb_io_requestor_0_s2_xcpt_ae_st;
assign core__io_dmem_ordered = _dcacheArb_io_requestor_0_ordered;
assign core__io_dmem_perf_release = _dcacheArb_io_requestor_0_perf_release;
assign core__io_dmem_perf_grant = _dcacheArb_io_requestor_0_perf_grant;
assign _core_io_ptw_status_debug = core__io_ptw_status_debug;
assign _core_io_ptw_pmp_cfg_l_0 = core__io_ptw_pmp_cfg_l_0;
assign _core_io_ptw_pmp_cfg_l_1 = core__io_ptw_pmp_cfg_l_1;
assign _core_io_ptw_pmp_cfg_l_2 = core__io_ptw_pmp_cfg_l_2;
assign _core_io_ptw_pmp_cfg_l_3 = core__io_ptw_pmp_cfg_l_3;
assign _core_io_ptw_pmp_cfg_l_4 = core__io_ptw_pmp_cfg_l_4;
assign _core_io_ptw_pmp_cfg_l_5 = core__io_ptw_pmp_cfg_l_5;
assign _core_io_ptw_pmp_cfg_l_6 = core__io_ptw_pmp_cfg_l_6;
assign _core_io_ptw_pmp_cfg_l_7 = core__io_ptw_pmp_cfg_l_7;
assign _core_io_ptw_pmp_cfg_a_0 = core__io_ptw_pmp_cfg_a_0;
assign _core_io_ptw_pmp_cfg_a_1 = core__io_ptw_pmp_cfg_a_1;
assign _core_io_ptw_pmp_cfg_a_2 = core__io_ptw_pmp_cfg_a_2;
assign _core_io_ptw_pmp_cfg_a_3 = core__io_ptw_pmp_cfg_a_3;
assign _core_io_ptw_pmp_cfg_a_4 = core__io_ptw_pmp_cfg_a_4;
assign _core_io_ptw_pmp_cfg_a_5 = core__io_ptw_pmp_cfg_a_5;
assign _core_io_ptw_pmp_cfg_a_6 = core__io_ptw_pmp_cfg_a_6;
assign _core_io_ptw_pmp_cfg_a_7 = core__io_ptw_pmp_cfg_a_7;
assign _core_io_ptw_pmp_cfg_x_0 = core__io_ptw_pmp_cfg_x_0;
assign _core_io_ptw_pmp_cfg_x_1 = core__io_ptw_pmp_cfg_x_1;
assign _core_io_ptw_pmp_cfg_x_2 = core__io_ptw_pmp_cfg_x_2;
assign _core_io_ptw_pmp_cfg_x_3 = core__io_ptw_pmp_cfg_x_3;
assign _core_io_ptw_pmp_cfg_x_4 = core__io_ptw_pmp_cfg_x_4;
assign _core_io_ptw_pmp_cfg_x_5 = core__io_ptw_pmp_cfg_x_5;
assign _core_io_ptw_pmp_cfg_x_6 = core__io_ptw_pmp_cfg_x_6;
assign _core_io_ptw_pmp_cfg_x_7 = core__io_ptw_pmp_cfg_x_7;
assign _core_io_ptw_pmp_cfg_w_0 = core__io_ptw_pmp_cfg_w_0;
assign _core_io_ptw_pmp_cfg_w_1 = core__io_ptw_pmp_cfg_w_1;
assign _core_io_ptw_pmp_cfg_w_2 = core__io_ptw_pmp_cfg_w_2;
assign _core_io_ptw_pmp_cfg_w_3 = core__io_ptw_pmp_cfg_w_3;
assign _core_io_ptw_pmp_cfg_w_4 = core__io_ptw_pmp_cfg_w_4;
assign _core_io_ptw_pmp_cfg_w_5 = core__io_ptw_pmp_cfg_w_5;
assign _core_io_ptw_pmp_cfg_w_6 = core__io_ptw_pmp_cfg_w_6;
assign _core_io_ptw_pmp_cfg_w_7 = core__io_ptw_pmp_cfg_w_7;
assign _core_io_ptw_pmp_cfg_r_0 = core__io_ptw_pmp_cfg_r_0;
assign _core_io_ptw_pmp_cfg_r_1 = core__io_ptw_pmp_cfg_r_1;
assign _core_io_ptw_pmp_cfg_r_2 = core__io_ptw_pmp_cfg_r_2;
assign _core_io_ptw_pmp_cfg_r_3 = core__io_ptw_pmp_cfg_r_3;
assign _core_io_ptw_pmp_cfg_r_4 = core__io_ptw_pmp_cfg_r_4;
assign _core_io_ptw_pmp_cfg_r_5 = core__io_ptw_pmp_cfg_r_5;
assign _core_io_ptw_pmp_cfg_r_6 = core__io_ptw_pmp_cfg_r_6;
assign _core_io_ptw_pmp_cfg_r_7 = core__io_ptw_pmp_cfg_r_7;
assign _core_io_ptw_pmp_addr_0 = core__io_ptw_pmp_addr_0;
assign _core_io_ptw_pmp_addr_1 = core__io_ptw_pmp_addr_1;
assign _core_io_ptw_pmp_addr_2 = core__io_ptw_pmp_addr_2;
assign _core_io_ptw_pmp_addr_3 = core__io_ptw_pmp_addr_3;
assign _core_io_ptw_pmp_addr_4 = core__io_ptw_pmp_addr_4;
assign _core_io_ptw_pmp_addr_5 = core__io_ptw_pmp_addr_5;
assign _core_io_ptw_pmp_addr_6 = core__io_ptw_pmp_addr_6;
assign _core_io_ptw_pmp_addr_7 = core__io_ptw_pmp_addr_7;
assign _core_io_ptw_pmp_mask_0 = core__io_ptw_pmp_mask_0;
assign _core_io_ptw_pmp_mask_1 = core__io_ptw_pmp_mask_1;
assign _core_io_ptw_pmp_mask_2 = core__io_ptw_pmp_mask_2;
assign _core_io_ptw_pmp_mask_3 = core__io_ptw_pmp_mask_3;
assign _core_io_ptw_pmp_mask_4 = core__io_ptw_pmp_mask_4;
assign _core_io_ptw_pmp_mask_5 = core__io_ptw_pmp_mask_5;
assign _core_io_ptw_pmp_mask_6 = core__io_ptw_pmp_mask_6;
assign _core_io_ptw_pmp_mask_7 = core__io_ptw_pmp_mask_7;
assign _core_io_ptw_customCSRs_csrs_0_value = core__io_ptw_customCSRs_csrs_0_value;
assign _core_io_wfi = core__io_wfi;
 
  assign auto_wfi_out_0=wfiNodeOut_0_REG; 
endmodule
 
module TLMonitor_25 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [3:0] io_in_a_bits_size,
  input [1:0] io_in_a_bits_source,
  input [31:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_b_ready,
  input io_in_b_valid,
  input [2:0] io_in_b_bits_opcode,
  input [1:0] io_in_b_bits_param,
  input [3:0] io_in_b_bits_size,
  input [1:0] io_in_b_bits_source,
  input [31:0] io_in_b_bits_address,
  input [7:0] io_in_b_bits_mask,
  input io_in_b_bits_corrupt,
  input io_in_c_ready,
  input io_in_c_valid,
  input [2:0] io_in_c_bits_opcode,
  input [2:0] io_in_c_bits_param,
  input [3:0] io_in_c_bits_size,
  input [1:0] io_in_c_bits_source,
  input [31:0] io_in_c_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [3:0] io_in_d_bits_size,
  input [1:0] io_in_d_bits_source,
  input [1:0] io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt,
  input io_in_e_ready,
  input io_in_e_valid,
  input [1:0] io_in_e_bits_sink) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire [26:0] _GEN={23'h0,io_in_a_bits_size} ;  
   wire [26:0] _GEN_0={23'h0,io_in_c_bits_size} ;  
   wire _a_first_T_1=io_in_a_ready&io_in_a_valid ;  
   reg [8:0] a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [3:0] size ;  
   reg [1:0] source ;  
   reg [31:0] address ;  
   wire _d_first_T_3=io_in_d_ready&io_in_d_valid ;  
   reg [8:0] d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [3:0] size_1 ;  
   reg [1:0] source_1 ;  
   reg [1:0] sink ;  
   reg denied ;  
   reg [8:0] b_first_counter ;  
   reg [2:0] opcode_2 ;  
   reg [1:0] param_2 ;  
   reg [3:0] size_2 ;  
   reg [1:0] source_2 ;  
   reg [31:0] address_1 ;  
   wire _c_first_T_1=io_in_c_ready&io_in_c_valid ;  
   reg [8:0] c_first_counter ;  
   reg [2:0] opcode_3 ;  
   reg [2:0] param_3 ;  
   reg [3:0] size_3 ;  
   reg [1:0] source_3 ;  
   reg [31:0] address_2 ;  
   reg [2:0] inflight ;  
   reg [11:0] inflight_opcodes ;  
   reg [23:0] inflight_sizes ;  
   reg [8:0] a_first_counter_1 ;  
   wire a_first_1=a_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_1 ;  
   wire d_first_1=d_first_counter_1==9'h0 ;  
   wire [11:0] _a_opcode_lookup_T_1=inflight_opcodes>>{8'h0,io_in_d_bits_source,2'h0} ;  
   wire [3:0] _GEN_1={2'h0,io_in_a_bits_source} ;  
   wire _GEN_2=_a_first_T_1&a_first_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [3:0] _GEN_3={2'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [2:0] inflight_1 ;  
   reg [23:0] inflight_sizes_1 ;  
   reg [8:0] c_first_counter_1 ;  
   wire c_first_1=c_first_counter_1==9'h0 ;  
   reg [8:0] d_first_counter_2 ;  
   wire d_first_2=d_first_counter_2==9'h0 ;  
   wire _GEN_4=io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1] ;  
   wire [3:0] _GEN_5={2'h0,io_in_c_bits_source} ;  
   wire _GEN_6=_c_first_T_1&c_first_1&_GEN_4 ;  
   reg [31:0] watchdog_1 ;  
   reg [3:0] inflight_2 ;  
   reg [8:0] d_first_counter_3 ;  
   wire d_first_3=d_first_counter_3==9'h0 ;  
   wire _GEN_7=_d_first_T_3&d_first_3&io_in_d_bits_opcode[2]&~(io_in_d_bits_opcode[1]) ;  
   wire [3:0] _GEN_8={2'h0,io_in_d_bits_sink} ;  
   wire [3:0] d_set=_GEN_7 ? 4'h1<<_GEN_8:4'h0 ;  
   wire _GEN_9=io_in_e_ready&io_in_e_valid ;  
   wire [3:0] _GEN_10={2'h0,io_in_e_bits_sink} ;  
   wire _source_ok_T=io_in_a_bits_source==2'h0 ;  
   wire _source_ok_T_1=io_in_a_bits_source==2'h1 ;  
   wire _source_ok_T_2=io_in_a_bits_source==2'h2 ;  
   wire source_ok=_source_ok_T|_source_ok_T_1|_source_ok_T_2 ;  
   wire [26:0] _is_aligned_mask_T_1=27'hFFF<<_GEN ;  
   wire [11:0] _GEN_11=io_in_a_bits_address[11:0]&~(_is_aligned_mask_T_1[11:0]) ;  
   wire _mask_T=io_in_a_bits_size>4'h2 ;  
   wire mask_size=io_in_a_bits_size[1:0]==2'h2 ;  
   wire mask_acc=_mask_T|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=_mask_T|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size[1:0]==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_12=io_in_a_bits_size<4'hD ;  
   wire _GEN_13=_GEN_12&(_source_ok_T|_source_ok_T_1|_source_ok_T_2) ;  
   wire _GEN_14=io_in_a_bits_size<4'h7 ;  
   wire _GEN_15=io_in_a_bits_address[31:28]==4'h8 ;  
   wire _GEN_16=_GEN_13&_GEN_14&_GEN_15 ;  
   wire _GEN_17=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_18=io_in_a_bits_address[31:12]==20'h0 ;  
   wire _GEN_19={io_in_a_bits_address[31:14],~(io_in_a_bits_address[13:12])}==20'h0 ;  
   wire _GEN_20={io_in_a_bits_address[31:17],~(io_in_a_bits_address[16])}==16'h0 ;  
   wire _GEN_21={io_in_a_bits_address[31:26],io_in_a_bits_address[25:16]^10'h200}==16'h0 ;  
   wire _GEN_22={io_in_a_bits_address[31:28],~(io_in_a_bits_address[27:26])}==6'h0 ;  
   wire _GEN_23={io_in_a_bits_address[31],~(io_in_a_bits_address[30:29])}==3'h0 ;  
   wire _GEN_24=_GEN_18|_GEN_19 ;  
   wire _GEN_25=_source_ok_T&io_in_a_bits_size==4'h6&_GEN_12&(_GEN_24|_GEN_20|_GEN_21|_GEN_22|_GEN_23|_GEN_15) ;  
   wire _GEN_26=io_in_a_bits_param>3'h2 ;  
   wire _GEN_27=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_28=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_29=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_30=_GEN_12&_GEN_19 ;  
   wire _GEN_31=io_in_a_bits_mask!=mask ;  
   wire _GEN_32=_GEN_13&(_GEN_30|_GEN_14&(_GEN_18|_GEN_21|_GEN_22|_GEN_15)|io_in_a_bits_size<4'h9&_GEN_23) ;  
   wire _GEN_33=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_34=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_35=_GEN_13&io_in_a_bits_size<4'h4&(_GEN_24|_GEN_21|_GEN_22) ;  
   wire _GEN_36=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_37=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_38=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire source_ok_1=io_in_d_bits_source==2'h0|io_in_d_bits_source==2'h1|io_in_d_bits_source==2'h2 ;  
   wire _GEN_39=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_40=io_in_d_bits_size<4'h3 ;  
   wire _GEN_41=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_42=io_in_d_bits_param==2'h2 ;  
   wire _GEN_43=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_44=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_45=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_46=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_47=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire [19:0] _GEN_48={io_in_b_bits_address[31:14],~(io_in_b_bits_address[13:12])} ;  
   wire [5:0] _GEN_49={io_in_b_bits_address[31:28],~(io_in_b_bits_address[27:26])} ;  
   wire [15:0] _GEN_50={io_in_b_bits_address[31:26],io_in_b_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_51={io_in_b_bits_address[31:17],~(io_in_b_bits_address[16])} ;  
   wire _GEN_52=io_in_b_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_53={io_in_b_bits_address[31],~(io_in_b_bits_address[30:29])} ;  
   wire address_ok=~(|_GEN_48)|~(|_GEN_49)|~(|_GEN_50)|~(|(io_in_b_bits_address[31:12]))|~(|_GEN_51)|~_GEN_52|~(|_GEN_53) ;  
   wire [26:0] _is_aligned_mask_T_4=27'hFFF<<io_in_b_bits_size ;  
   wire [11:0] _GEN_54=io_in_b_bits_address[11:0]&~(_is_aligned_mask_T_4[11:0]) ;  
   wire _mask_T_1=io_in_b_bits_size>4'h2 ;  
   wire mask_size_3=io_in_b_bits_size[1:0]==2'h2 ;  
   wire mask_acc_14=_mask_T_1|mask_size_3&~(io_in_b_bits_address[2]) ;  
   wire mask_acc_15=_mask_T_1|mask_size_3&io_in_b_bits_address[2] ;  
   wire mask_size_4=io_in_b_bits_size[1:0]==2'h1 ;  
   wire mask_eq_16=~(io_in_b_bits_address[2])&~(io_in_b_bits_address[1]) ;  
   wire mask_acc_16=mask_acc_14|mask_size_4&mask_eq_16 ;  
   wire mask_eq_17=~(io_in_b_bits_address[2])&io_in_b_bits_address[1] ;  
   wire mask_acc_17=mask_acc_14|mask_size_4&mask_eq_17 ;  
   wire mask_eq_18=io_in_b_bits_address[2]&~(io_in_b_bits_address[1]) ;  
   wire mask_acc_18=mask_acc_15|mask_size_4&mask_eq_18 ;  
   wire mask_eq_19=io_in_b_bits_address[2]&io_in_b_bits_address[1] ;  
   wire mask_acc_19=mask_acc_15|mask_size_4&mask_eq_19 ;  
   wire [7:0] mask_1={mask_acc_19|mask_eq_19&io_in_b_bits_address[0],mask_acc_19|mask_eq_19&~(io_in_b_bits_address[0]),mask_acc_18|mask_eq_18&io_in_b_bits_address[0],mask_acc_18|mask_eq_18&~(io_in_b_bits_address[0]),mask_acc_17|mask_eq_17&io_in_b_bits_address[0],mask_acc_17|mask_eq_17&~(io_in_b_bits_address[0]),mask_acc_16|mask_eq_16&io_in_b_bits_address[0],mask_acc_16|mask_eq_16&~(io_in_b_bits_address[0])} ;  
   wire _GEN_55=io_in_b_valid&io_in_b_bits_opcode==3'h6&~reset ;  
   wire _GEN_56={io_in_b_bits_source==2'h2,io_in_b_bits_source==2'h1}!=io_in_b_bits_source ;  
   wire _GEN_57=io_in_b_bits_mask!=mask_1 ;  
   wire _GEN_58=io_in_b_valid&io_in_b_bits_opcode==3'h4&~reset ;  
   wire _GEN_59=io_in_b_valid&io_in_b_bits_opcode==3'h0&~reset ;  
   wire _GEN_60=io_in_b_valid&io_in_b_bits_opcode==3'h1&~reset ;  
   wire _GEN_61=io_in_b_valid&io_in_b_bits_opcode==3'h2&~reset ;  
   wire _GEN_62=io_in_b_valid&io_in_b_bits_opcode==3'h3&~reset ;  
   wire _GEN_63=io_in_b_valid&io_in_b_bits_opcode==3'h5&~reset ;  
   wire _source_ok_T_8=io_in_c_bits_source==2'h0 ;  
   wire _source_ok_T_9=io_in_c_bits_source==2'h1 ;  
   wire _source_ok_T_10=io_in_c_bits_source==2'h2 ;  
   wire source_ok_2=_source_ok_T_8|_source_ok_T_9|_source_ok_T_10 ;  
   wire [26:0] _is_aligned_mask_T_7=27'hFFF<<_GEN_0 ;  
   wire [11:0] _GEN_64=io_in_c_bits_address[11:0]&~(_is_aligned_mask_T_7[11:0]) ;  
   wire [19:0] _GEN_65={io_in_c_bits_address[31:14],~(io_in_c_bits_address[13:12])} ;  
   wire [5:0] _GEN_66={io_in_c_bits_address[31:28],~(io_in_c_bits_address[27:26])} ;  
   wire [15:0] _GEN_67={io_in_c_bits_address[31:26],io_in_c_bits_address[25:16]^10'h200} ;  
   wire [15:0] _GEN_68={io_in_c_bits_address[31:17],~(io_in_c_bits_address[16])} ;  
   wire _GEN_69=io_in_c_bits_address[31:28]!=4'h8 ;  
   wire [2:0] _GEN_70={io_in_c_bits_address[31],~(io_in_c_bits_address[30:29])} ;  
   wire address_ok_1=~(|_GEN_65)|~(|_GEN_66)|~(|_GEN_67)|~(|(io_in_c_bits_address[31:12]))|~(|_GEN_68)|~_GEN_69|~(|_GEN_70) ;  
   wire _GEN_71=io_in_c_valid&io_in_c_bits_opcode==3'h4&~reset ;  
   wire _GEN_72=io_in_c_bits_size<4'h3 ;  
   wire _GEN_73=io_in_c_valid&io_in_c_bits_opcode==3'h5&~reset ;  
   wire _GEN_74=io_in_c_bits_size<4'hD ;  
   wire _GEN_75=_GEN_74&(_source_ok_T_8|_source_ok_T_9|_source_ok_T_10)&io_in_c_bits_size<4'h7&~_GEN_69 ;  
   wire _GEN_76=io_in_c_valid&io_in_c_bits_opcode==3'h6&~reset ;  
   wire _GEN_77=_source_ok_T_8&io_in_c_bits_size==4'h6&_GEN_74&(~(|(io_in_c_bits_address[31:12]))|~(|_GEN_65)|~(|_GEN_68)|~(|_GEN_67)|~(|_GEN_66)|~(|_GEN_70)|~_GEN_69) ;  
   wire _GEN_78=io_in_c_valid&(&io_in_c_bits_opcode)&~reset ;  
   wire _GEN_79=io_in_c_valid&io_in_c_bits_opcode==3'h0&~reset ;  
   wire _GEN_80=io_in_c_valid&io_in_c_bits_opcode==3'h1&~reset ;  
   wire _GEN_81=io_in_c_valid&io_in_c_bits_opcode==3'h2&~reset ;  
   wire _GEN_82=io_in_a_valid&(|a_first_counter)&~reset ;  
   wire _GEN_83=io_in_d_valid&(|d_first_counter)&~reset ;  
   wire _GEN_84=io_in_b_valid&(|b_first_counter)&~reset ;  
   wire _GEN_85=io_in_c_valid&(|c_first_counter)&~reset ;  
   wire [23:0] _GEN_86={19'h0,io_in_d_bits_source,3'h0} ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&a_first_1 ;  
   wire [3:0] _a_set_wo_ready_T=4'h1<<_GEN_1 ;  
   wire [2:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[2:0]:3'h0 ;  
   wire _GEN_87=io_in_d_valid&d_first_1 ;  
   wire _GEN_88=_GEN_87&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [2:0] _GEN_89={1'h0,io_in_d_bits_source} ;  
   wire _GEN_90=_GEN_88&same_cycle_resp&~reset ;  
   wire _GEN_91=_GEN_88&~same_cycle_resp&~reset ;  
   wire [7:0] _GEN_92={4'h0,io_in_d_bits_size} ;  
   wire _same_cycle_resp_T_3=io_in_c_valid&c_first_1 ;  
   wire [3:0] _c_set_wo_ready_T=4'h1<<_GEN_5 ;  
   wire [2:0] c_set_wo_ready=_same_cycle_resp_T_3&_GEN_4 ? _c_set_wo_ready_T[2:0]:3'h0 ;  
   wire _GEN_93=io_in_d_valid&d_first_2 ;  
   wire _GEN_94=_GEN_93&d_release_ack ;  
   wire same_cycle_resp_1=_same_cycle_resp_T_3&io_in_c_bits_opcode[2]&io_in_c_bits_opcode[1]&io_in_c_bits_source==io_in_d_bits_source ;  
   wire [2:0] _GEN_95=inflight>>io_in_a_bits_source ;  
   wire [2:0] _GEN_96=inflight>>_GEN_89 ;  
   wire [23:0] _a_size_lookup_T_1=inflight_sizes>>_GEN_86 ;  
   wire [3:0] _d_clr_wo_ready_T=4'h1<<_GEN_3 ;  
   wire [2:0] _GEN_97=inflight_1>>io_in_c_bits_source ;  
   wire [2:0] _GEN_98=inflight_1>>_GEN_89 ;  
   wire [23:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN_86 ;  
   wire [3:0] _d_clr_wo_ready_T_1=4'h1<<_GEN_3 ;  
   wire [3:0] _GEN_99=inflight_2>>_GEN_8 ;  
   wire [3:0] _GEN_100=(d_set|inflight_2)>>_GEN_10 ;  
  always @( posedge clock)
       begin 
         if (_GEN_17&~_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_GEN_25)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~_mask_T)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_26)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_27)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~(_GEN_30|_GEN_14&(_GEN_18|_GEN_20|_GEN_21|_GEN_22|_GEN_23|_GEN_15)))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_33&_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~_GEN_32)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_34&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~_GEN_35)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_36&_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~_GEN_35)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_37&_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&~(_GEN_13&_GEN_30))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&~source_ok)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&(|_GEN_11))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_38&_GEN_31)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&_GEN_40)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_39&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&_GEN_40)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&_GEN_42)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_41&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&_GEN_40)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&_GEN_42)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_43&~_GEN_44)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_45&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_46&~_GEN_44)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&~source_ok_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_47&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_b_valid&~reset&(&io_in_b_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'B' channel has invalid opcode (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&~(io_in_b_bits_source==2'h0&io_in_b_bits_size==4'h6&io_in_b_bits_size<4'hD&(~(|(io_in_b_bits_address[31:12]))|~(|_GEN_48)|~(|_GEN_51)|~(|_GEN_50)|~(|_GEN_49)|~(|_GEN_53)|~_GEN_52)))
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries source that is not first source (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&(&io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe carries invalid cap param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&_GEN_57)
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_55&io_in_b_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'B' channel Probe is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Get carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel Get carries source that is not first source (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'B' channel Get address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&(|io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel Get carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&_GEN_57)
            begin 
              if (1)$display("Assertion failed: 'B' channel Get contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_58&io_in_b_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'B' channel Get is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull carries source that is not first source (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&(|io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_59&_GEN_57)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutFull contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&(|io_in_b_bits_param))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_60&(|(io_in_b_bits_mask&~mask_1)))
            begin 
              if (1)$display("Assertion failed: 'B' channel PutPartial contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_61&_GEN_57)
            begin 
              if (1)$display("Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_62)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Logical type unsupported by client (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_62&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_62&_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical carries source that is not first source (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_62&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_62&_GEN_57)
            begin 
              if (1)$display("Assertion failed: 'B' channel Logical contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63)
            begin 
              if (1)$display("Assertion failed: 'B' channel carries Hint type unsupported by client (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&~address_ok)
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&_GEN_56)
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint carries source that is not first source (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&(|_GEN_54))
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&_GEN_57)
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint contains invalid mask (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_63&io_in_b_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'B' channel Hint is corrupt (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&_GEN_72)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(|_GEN_64))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_71&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&_GEN_72)
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&(|_GEN_64))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_73&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&~_GEN_75)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&~_GEN_77)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&_GEN_72)
            begin 
              if (1)$display("Assertion failed: 'C' channel Release smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&(|_GEN_64))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_76&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel Release carries invalid report param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&~_GEN_75)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&~_GEN_77)
            begin 
              if (1)$display("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&_GEN_72)
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&(|_GEN_64))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_78&(&(io_in_c_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_79&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_79&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_79&(|_GEN_64))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_79&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&(|_GEN_64))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_80&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&~address_ok_1)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&~source_ok_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&(|_GEN_64))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck address not aligned to size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_81&(|io_in_c_bits_param))
            begin 
              if (1)$display("Assertion failed: 'C' channel HintAck carries invalid param (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_82&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_83&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&io_in_b_bits_opcode!=opcode_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&io_in_b_bits_param!=param_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel param changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&io_in_b_bits_size!=size_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&io_in_b_bits_source!=source_2)
            begin 
              if (1)$display("Assertion failed: 'B' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_84&io_in_b_bits_address!=address_1)
            begin 
              if (1)$display("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_85&io_in_c_bits_opcode!=opcode_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_85&io_in_c_bits_param!=param_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel param changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_85&io_in_c_bits_size!=size_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel size changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_85&io_in_c_bits_source!=source_3)
            begin 
              if (1)$display("Assertion failed: 'C' channel source changed within multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_85&io_in_c_bits_address!=address_2)
            begin 
              if (1)$display("Assertion failed: 'C' channel address changed with multibeat operation (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~reset&_GEN_95[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_88&~reset&~(_GEN_96[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_90&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_90&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_91&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_91&_GEN_92!={1'h0,_a_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_87&a_first_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_88 ? _d_clr_wo_ready_T[2:0]:3'h0)|a_set_wo_ready==3'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==3'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~reset&_GEN_97[0])
            begin 
              if (1)$display("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_94&~reset&~(_GEN_98[0]|same_cycle_resp_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_94&same_cycle_resp_1&~reset&io_in_d_bits_size!=io_in_c_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_94&~same_cycle_resp_1&~reset&_GEN_92!={1'h0,_c_size_lookup_T_1[7:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_93&c_first_1&io_in_c_valid&io_in_c_bits_source==io_in_d_bits_source&d_release_ack&~(io_in_c_bits_opcode==3'h4|io_in_c_bits_opcode==3'h5)&~reset&~(~io_in_d_ready|io_in_c_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if ((|c_set_wo_ready)&~reset&c_set_wo_ready==(_GEN_94 ? _d_clr_wo_ready_T_1[2:0]:3'h0))
            begin 
              if (1)$display("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==3'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~reset&_GEN_99[0])
            begin 
              if (1)$display("Assertion failed: 'D' channel re-used a sink ID (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~reset&~(_GEN_100[0]))
            begin 
              if (1)$display("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at src/main/scala/tilelink/CrossingHelper.scala:61:80)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [26:0] _a_first_beats1_decode_T_1=27'hFFF<<_GEN ;  
   wire [26:0] _a_first_beats1_decode_T_5=27'hFFF<<_GEN ;  
   wire [26:0] _GEN_101={23'h0,io_in_d_bits_size} ;  
   wire [26:0] _d_first_beats1_decode_T_1=27'hFFF<<_GEN_101 ;  
   wire [26:0] _d_first_beats1_decode_T_5=27'hFFF<<_GEN_101 ;  
   wire [26:0] _d_first_beats1_decode_T_9=27'hFFF<<_GEN_101 ;  
   wire [26:0] _d_first_beats1_decode_T_13=27'hFFF<<_GEN_101 ;  
   wire [26:0] _c_first_beats1_decode_T_1=27'hFFF<<_GEN_0 ;  
   wire [26:0] _c_first_beats1_decode_T_5=27'hFFF<<_GEN_0 ;  
   wire _GEN_102=_d_first_T_3&d_first_1&~d_release_ack ;  
   wire [46:0] _GEN_103={42'h0,io_in_d_bits_source,3'h0} ;  
   wire _GEN_104=_d_first_T_3&d_first_2&d_release_ack ;  
   wire [3:0] _d_clr_T=4'h1<<_GEN_3 ;  
   wire [3:0] _a_set_T=4'h1<<_GEN_1 ;  
   wire [46:0] _d_opcodes_clr_T_5=47'hF<<{43'h0,io_in_d_bits_source,2'h0} ;  
   wire [34:0] _a_opcodes_set_T_1={31'h0,_GEN_2 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{31'h0,io_in_a_bits_source,2'h0} ;  
   wire [46:0] _d_sizes_clr_T_5=47'hFF<<_GEN_103 ;  
   wire [35:0] _a_sizes_set_T_1={31'h0,_GEN_2 ? {io_in_a_bits_size,1'h1}:5'h0}<<{31'h0,io_in_a_bits_source,3'h0} ;  
   wire [3:0] _d_clr_T_1=4'h1<<_GEN_3 ;  
   wire [3:0] _c_set_T=4'h1<<_GEN_5 ;  
   wire [46:0] _d_sizes_clr_T_11=47'hFF<<_GEN_103 ;  
   wire [35:0] _c_sizes_set_T_1={31'h0,_GEN_6 ? {io_in_c_bits_size,1'h1}:5'h0}<<{31'h0,io_in_c_bits_source,3'h0} ;  
   wire b_first_done=io_in_b_ready&io_in_b_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=9'h0;
              d_first_counter <=9'h0;
              b_first_counter <=9'h0;
              c_first_counter <=9'h0;
              inflight <=3'h0;
              inflight_opcodes <=12'h0;
              inflight_sizes <=24'h0;
              a_first_counter_1 <=9'h0;
              d_first_counter_1 <=9'h0;
              watchdog <=32'h0;
              inflight_1 <=3'h0;
              inflight_sizes_1 <=24'h0;
              c_first_counter_1 <=9'h0;
              d_first_counter_2 <=9'h0;
              watchdog_1 <=32'h0;
              inflight_2 <=4'h0;
              d_first_counter_3 <=9'h0;
            end 
          else 
            begin 
              if (_a_first_T_1)
                 begin 
                   if (|a_first_counter)
                      a_first_counter <=a_first_counter-9'h1;
                    else 
                      a_first_counter <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_1[11:3]);
                   if (a_first_1)
                      a_first_counter_1 <=io_in_a_bits_opcode[2] ? 9'h0:~(_a_first_beats1_decode_T_5[11:3]);
                    else 
                      a_first_counter_1 <=a_first_counter_1-9'h1;
                 end 
              if (_d_first_T_3)
                 begin 
                   if (|d_first_counter)
                      d_first_counter <=d_first_counter-9'h1;
                    else 
                      d_first_counter <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_1[11:3]):9'h0;
                   if (d_first_1)
                      d_first_counter_1 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      d_first_counter_1 <=d_first_counter_1-9'h1;
                   if (d_first_2)
                      d_first_counter_2 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_9[11:3]):9'h0;
                    else 
                      d_first_counter_2 <=d_first_counter_2-9'h1;
                   if (d_first_3)
                      d_first_counter_3 <=io_in_d_bits_opcode[0] ? ~(_d_first_beats1_decode_T_13[11:3]):9'h0;
                    else 
                      d_first_counter_3 <=d_first_counter_3-9'h1;
                 end 
              if (b_first_done)
                 begin 
                   if (|b_first_counter)
                      b_first_counter <=b_first_counter-9'h1;
                    else 
                      b_first_counter <=9'h0;
                 end 
              if (_c_first_T_1)
                 begin 
                   if (|c_first_counter)
                      c_first_counter <=c_first_counter-9'h1;
                    else 
                      c_first_counter <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_1[11:3]):9'h0;
                   if (c_first_1)
                      c_first_counter_1 <=io_in_c_bits_opcode[0] ? ~(_c_first_beats1_decode_T_5[11:3]):9'h0;
                    else 
                      c_first_counter_1 <=c_first_counter_1-9'h1;
                 end 
              inflight <=(inflight|(_GEN_2 ? _a_set_T[2:0]:3'h0))&~(_GEN_102 ? _d_clr_T[2:0]:3'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_2 ? _a_opcodes_set_T_1[11:0]:12'h0))&~(_GEN_102 ? _d_opcodes_clr_T_5[11:0]:12'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_2 ? _a_sizes_set_T_1[23:0]:24'h0))&~(_GEN_102 ? _d_sizes_clr_T_5[23:0]:24'h0);
              if (_a_first_T_1|_d_first_T_3)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=(inflight_1|(_GEN_6 ? _c_set_T[2:0]:3'h0))&~(_GEN_104 ? _d_clr_T_1[2:0]:3'h0);
              inflight_sizes_1 <=(inflight_sizes_1|(_GEN_6 ? _c_sizes_set_T_1[23:0]:24'h0))&~(_GEN_104 ? _d_sizes_clr_T_11[23:0]:24'h0);
              if (_c_first_T_1|_d_first_T_3)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
              inflight_2 <=(inflight_2|d_set)&~(_GEN_9 ? 4'h1<<_GEN_10:4'h0);
            end 
         if (_a_first_T_1&~(|a_first_counter))
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (_d_first_T_3&~(|d_first_counter))
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
         if (b_first_done&~(|b_first_counter))
            begin 
              opcode_2 <=io_in_b_bits_opcode;
              param_2 <=io_in_b_bits_param;
              size_2 <=io_in_b_bits_size;
              source_2 <=io_in_b_bits_source;
              address_1 <=io_in_b_bits_address;
            end 
         if (_c_first_T_1&~(|c_first_counter))
            begin 
              opcode_3 <=io_in_c_bits_opcode;
              param_3 <=io_in_c_bits_param;
              size_3 <=io_in_c_bits_size;
              source_3 <=io_in_c_bits_source;
              address_2 <=io_in_c_bits_address;
            end 
       end
  
endmodule
 
module Queue_78 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [1:0] io_enq_bits_source,
  input [31:0] io_enq_bits_address,
  input [7:0] io_enq_bits_mask,
  input [63:0] io_enq_bits_data,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [1:0] io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output [63:0] io_deq_bits_data,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x3 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_2x2 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_addr_2x32 ram_address_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_address),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_address)); 
  ram_2x8 ram_mask_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_mask),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_mask)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(1'h0)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_79 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [1:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [1:0] io_enq_bits_source,
  input [1:0] io_enq_bits_sink,
  input io_enq_bits_denied,
  input [63:0] io_enq_bits_data,
  input io_enq_bits_corrupt,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [1:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [1:0] io_deq_bits_source,
  output [1:0] io_deq_bits_sink,
  output io_deq_bits_denied,
  output [63:0] io_deq_bits_data,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x2 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_2x2 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_2x2 ram_sink_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_sink),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_sink)); 
  ram_2x1 ram_denied_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_denied),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_denied)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_corrupt)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module ram_2x52 (
  input R0_addr,
  input R0_en,
  input R0_clk,
  output [51:0] R0_data,
  input W0_addr,
  input W0_en,
  input W0_clk,
  input [51:0] W0_data) ; 
   reg [51:0] Memory[0:1] ;  
  always @( posedge W0_clk)
       begin 
         if (W0_en&1'h1)
            Memory [W0_addr]<=W0_data;
       end
  
  assign R0_data=R0_en ? Memory[R0_addr]:52'bx; 
endmodule
 
module Queue_80 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [1:0] io_enq_bits_param,
  input [31:0] io_enq_bits_address,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [1:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [1:0] io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0] io_deq_bits_mask,
  output io_deq_bits_corrupt) ; 
   wire [51:0] _ram_ext_R0_data ;  
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x52 ram_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(_ram_ext_R0_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data({9'hFF,io_enq_bits_address,6'h6,io_enq_bits_param,3'h6})); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
  assign io_deq_bits_opcode=_ram_ext_R0_data[2:0]; 
  assign io_deq_bits_param=_ram_ext_R0_data[4:3]; 
  assign io_deq_bits_size=_ram_ext_R0_data[8:5]; 
  assign io_deq_bits_source=_ram_ext_R0_data[10:9]; 
  assign io_deq_bits_address=_ram_ext_R0_data[42:11]; 
  assign io_deq_bits_mask=_ram_ext_R0_data[50:43]; 
  assign io_deq_bits_corrupt=_ram_ext_R0_data[51]; 
endmodule
 
module Queue_81 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [2:0] io_enq_bits_param,
  input [3:0] io_enq_bits_size,
  input [1:0] io_enq_bits_source,
  input [31:0] io_enq_bits_address,
  input [63:0] io_enq_bits_data,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [1:0] io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [63:0] io_deq_bits_data,
  output io_deq_bits_corrupt) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x3 ram_opcode_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_opcode),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_opcode)); 
  ram_2x3 ram_param_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_param),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_param)); 
  ram_2x4 ram_size_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_size),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_size)); 
  ram_2x2 ram_source_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_source),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_source)); 
  ram_addr_2x32 ram_address_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_address),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_address)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x1 ram_corrupt_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_corrupt),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(1'h0)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_82 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [1:0] io_enq_bits_sink,
  output io_deq_valid,
  output [1:0] io_deq_bits_sink) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (~empty)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==~empty))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x2 ram_sink_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_sink),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_sink)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module TLBuffer_10 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [3:0] auto_in_a_bits_size,
  input [1:0] auto_in_a_bits_source,
  input [31:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [2:0] auto_in_b_bits_opcode,
  output [1:0] auto_in_b_bits_param,
  output [3:0] auto_in_b_bits_size,
  output [1:0] auto_in_b_bits_source,
  output [31:0] auto_in_b_bits_address,
  output [7:0] auto_in_b_bits_mask,
  output auto_in_b_bits_corrupt,
  output auto_in_c_ready,
  input auto_in_c_valid,
  input [2:0] auto_in_c_bits_opcode,
  input [2:0] auto_in_c_bits_param,
  input [3:0] auto_in_c_bits_size,
  input [1:0] auto_in_c_bits_source,
  input [31:0] auto_in_c_bits_address,
  input [63:0] auto_in_c_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [3:0] auto_in_d_bits_size,
  output [1:0] auto_in_d_bits_source,
  output [1:0] auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [63:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  output auto_in_e_ready,
  input auto_in_e_valid,
  input [1:0] auto_in_e_bits_sink,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [3:0] auto_out_a_bits_size,
  output [1:0] auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0] auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [1:0] auto_out_b_bits_param,
  input [31:0] auto_out_b_bits_address,
  input auto_out_c_ready,
  output auto_out_c_valid,
  output [2:0] auto_out_c_bits_opcode,
  output [2:0] auto_out_c_bits_param,
  output [3:0] auto_out_c_bits_size,
  output [1:0] auto_out_c_bits_source,
  output [31:0] auto_out_c_bits_address,
  output [63:0] auto_out_c_bits_data,
  output auto_out_c_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_param,
  input [3:0] auto_out_d_bits_size,
  input [1:0] auto_out_d_bits_source,
  input [1:0] auto_out_d_bits_sink,
  input auto_out_d_bits_denied,
  input [63:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt,
  output auto_out_e_valid,
  output [1:0] auto_out_e_bits_sink) ; 
   wire _nodeOut_e_q_io_enq_ready ;  
   wire _nodeOut_c_q_io_enq_ready ;  
   wire _nodeIn_b_q_io_deq_valid ;  
   wire [2:0] _nodeIn_b_q_io_deq_bits_opcode ;  
   wire [1:0] _nodeIn_b_q_io_deq_bits_param ;  
   wire [3:0] _nodeIn_b_q_io_deq_bits_size ;  
   wire [1:0] _nodeIn_b_q_io_deq_bits_source ;  
   wire [31:0] _nodeIn_b_q_io_deq_bits_address ;  
   wire [7:0] _nodeIn_b_q_io_deq_bits_mask ;  
   wire _nodeIn_b_q_io_deq_bits_corrupt ;  
   wire _nodeIn_d_q_io_deq_valid ;  
   wire [2:0] _nodeIn_d_q_io_deq_bits_opcode ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_param ;  
   wire [3:0] _nodeIn_d_q_io_deq_bits_size ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_source ;  
   wire [1:0] _nodeIn_d_q_io_deq_bits_sink ;  
   wire _nodeIn_d_q_io_deq_bits_denied ;  
   wire _nodeIn_d_q_io_deq_bits_corrupt ;  
   wire _nodeOut_a_q_io_enq_ready ;  
  TLMonitor_25 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_nodeOut_a_q_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_b_ready(auto_in_b_ready),.io_in_b_valid(_nodeIn_b_q_io_deq_valid),.io_in_b_bits_opcode(_nodeIn_b_q_io_deq_bits_opcode),.io_in_b_bits_param(_nodeIn_b_q_io_deq_bits_param),.io_in_b_bits_size(_nodeIn_b_q_io_deq_bits_size),.io_in_b_bits_source(_nodeIn_b_q_io_deq_bits_source),.io_in_b_bits_address(_nodeIn_b_q_io_deq_bits_address),.io_in_b_bits_mask(_nodeIn_b_q_io_deq_bits_mask),.io_in_b_bits_corrupt(_nodeIn_b_q_io_deq_bits_corrupt),.io_in_c_ready(_nodeOut_c_q_io_enq_ready),.io_in_c_valid(auto_in_c_valid),.io_in_c_bits_opcode(auto_in_c_bits_opcode),.io_in_c_bits_param(auto_in_c_bits_param),.io_in_c_bits_size(auto_in_c_bits_size),.io_in_c_bits_source(auto_in_c_bits_source),.io_in_c_bits_address(auto_in_c_bits_address),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(_nodeIn_d_q_io_deq_valid),.io_in_d_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_in_d_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_in_d_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_in_d_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_in_d_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_in_d_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_in_d_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt),.io_in_e_ready(_nodeOut_e_q_io_enq_ready),.io_in_e_valid(auto_in_e_valid),.io_in_e_bits_sink(auto_in_e_bits_sink)); 
  Queue_78 nodeOut_a_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_a_q_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_param(auto_in_a_bits_param),.io_enq_bits_size(auto_in_a_bits_size),.io_enq_bits_source(auto_in_a_bits_source),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_data(auto_in_a_bits_data),.io_deq_ready(auto_out_a_ready),.io_deq_valid(auto_out_a_valid),.io_deq_bits_opcode(auto_out_a_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(auto_out_a_bits_size),.io_deq_bits_source(auto_out_a_bits_source),.io_deq_bits_address(auto_out_a_bits_address),.io_deq_bits_mask(auto_out_a_bits_mask),.io_deq_bits_data(auto_out_a_bits_data),.io_deq_bits_corrupt(auto_out_a_bits_corrupt)); 
  Queue_79 nodeIn_d_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_d_ready),.io_enq_valid(auto_out_d_valid),.io_enq_bits_opcode(auto_out_d_bits_opcode),.io_enq_bits_param(auto_out_d_bits_param),.io_enq_bits_size(auto_out_d_bits_size),.io_enq_bits_source(auto_out_d_bits_source),.io_enq_bits_sink(auto_out_d_bits_sink),.io_enq_bits_denied(auto_out_d_bits_denied),.io_enq_bits_data(auto_out_d_bits_data),.io_enq_bits_corrupt(auto_out_d_bits_corrupt),.io_deq_ready(auto_in_d_ready),.io_deq_valid(_nodeIn_d_q_io_deq_valid),.io_deq_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),.io_deq_bits_param(_nodeIn_d_q_io_deq_bits_param),.io_deq_bits_size(_nodeIn_d_q_io_deq_bits_size),.io_deq_bits_source(_nodeIn_d_q_io_deq_bits_source),.io_deq_bits_sink(_nodeIn_d_q_io_deq_bits_sink),.io_deq_bits_denied(_nodeIn_d_q_io_deq_bits_denied),.io_deq_bits_data(auto_in_d_bits_data),.io_deq_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)); 
  Queue_80 nodeIn_b_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_b_ready),.io_enq_valid(auto_out_b_valid),.io_enq_bits_param(auto_out_b_bits_param),.io_enq_bits_address(auto_out_b_bits_address),.io_deq_ready(auto_in_b_ready),.io_deq_valid(_nodeIn_b_q_io_deq_valid),.io_deq_bits_opcode(_nodeIn_b_q_io_deq_bits_opcode),.io_deq_bits_param(_nodeIn_b_q_io_deq_bits_param),.io_deq_bits_size(_nodeIn_b_q_io_deq_bits_size),.io_deq_bits_source(_nodeIn_b_q_io_deq_bits_source),.io_deq_bits_address(_nodeIn_b_q_io_deq_bits_address),.io_deq_bits_mask(_nodeIn_b_q_io_deq_bits_mask),.io_deq_bits_corrupt(_nodeIn_b_q_io_deq_bits_corrupt)); 
  Queue_81 nodeOut_c_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_c_q_io_enq_ready),.io_enq_valid(auto_in_c_valid),.io_enq_bits_opcode(auto_in_c_bits_opcode),.io_enq_bits_param(auto_in_c_bits_param),.io_enq_bits_size(auto_in_c_bits_size),.io_enq_bits_source(auto_in_c_bits_source),.io_enq_bits_address(auto_in_c_bits_address),.io_enq_bits_data(auto_in_c_bits_data),.io_deq_ready(auto_out_c_ready),.io_deq_valid(auto_out_c_valid),.io_deq_bits_opcode(auto_out_c_bits_opcode),.io_deq_bits_param(auto_out_c_bits_param),.io_deq_bits_size(auto_out_c_bits_size),.io_deq_bits_source(auto_out_c_bits_source),.io_deq_bits_address(auto_out_c_bits_address),.io_deq_bits_data(auto_out_c_bits_data),.io_deq_bits_corrupt(auto_out_c_bits_corrupt)); 
  Queue_82 nodeOut_e_q(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_e_q_io_enq_ready),.io_enq_valid(auto_in_e_valid),.io_enq_bits_sink(auto_in_e_bits_sink),.io_deq_valid(auto_out_e_valid),.io_deq_bits_sink(auto_out_e_bits_sink)); 
  assign auto_in_a_ready=_nodeOut_a_q_io_enq_ready; 
  assign auto_in_b_valid=_nodeIn_b_q_io_deq_valid; 
  assign auto_in_b_bits_opcode=_nodeIn_b_q_io_deq_bits_opcode; 
  assign auto_in_b_bits_param=_nodeIn_b_q_io_deq_bits_param; 
  assign auto_in_b_bits_size=_nodeIn_b_q_io_deq_bits_size; 
  assign auto_in_b_bits_source=_nodeIn_b_q_io_deq_bits_source; 
  assign auto_in_b_bits_address=_nodeIn_b_q_io_deq_bits_address; 
  assign auto_in_b_bits_mask=_nodeIn_b_q_io_deq_bits_mask; 
  assign auto_in_b_bits_corrupt=_nodeIn_b_q_io_deq_bits_corrupt; 
  assign auto_in_c_ready=_nodeOut_c_q_io_enq_ready; 
  assign auto_in_d_valid=_nodeIn_d_q_io_deq_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_q_io_deq_bits_opcode; 
  assign auto_in_d_bits_param=_nodeIn_d_q_io_deq_bits_param; 
  assign auto_in_d_bits_size=_nodeIn_d_q_io_deq_bits_size; 
  assign auto_in_d_bits_source=_nodeIn_d_q_io_deq_bits_source; 
  assign auto_in_d_bits_sink=_nodeIn_d_q_io_deq_bits_sink; 
  assign auto_in_d_bits_denied=_nodeIn_d_q_io_deq_bits_denied; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_q_io_deq_bits_corrupt; 
  assign auto_in_e_ready=_nodeOut_e_q_io_enq_ready; 
endmodule
 
module SynchronizerShiftReg_w1_d3 (
  input clock,
  input io_d,
  output io_q) ; 
  NonSyncResetSynchronizerPrimitiveShiftReg_d3 output_chain(.clock(clock),.io_d(io_d),.io_q(io_q)); 
endmodule
 
module IntSyncAsyncCrossingSink_1 (
  input clock,
  input auto_in_sync_0,
  output auto_out_0) ; 
  SynchronizerShiftReg_w1_d3 chain(.clock(clock),.io_d(auto_in_sync_0),.io_q(auto_out_0)); 
endmodule
 
module IntSyncSyncCrossingSink (
  input auto_in_sync_0,
  input auto_in_sync_1,
  output auto_out_0,
  output auto_out_1) ; 
  assign auto_out_0=auto_in_sync_0; 
  assign auto_out_1=auto_in_sync_1; 
endmodule
 
module IntSyncSyncCrossingSink_1 (
  input auto_in_sync_0,
  output auto_out_0) ; 
  assign auto_out_0=auto_in_sync_0; 
endmodule
 
module AsyncResetRegVec_w1_i0 (
  input clock,
  input reset,
  input io_d,
  output io_q) ; 
   reg reg_0 ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            reg_0 <=1'h0;
          else 
            reg_0 <=io_d;
       end
  
  assign io_q=reg_0; 
endmodule
 
module IntSyncCrossingSource_1 (
  input clock,
  input reset,
  input auto_in_0,
  output auto_out_sync_0) ; 
  AsyncResetRegVec_w1_i0 reg_0(.clock(clock),.reset(reset),.io_d(auto_in_0),.io_q(auto_out_sync_0)); 
endmodule
 
module TilePRCIDomain (
  input auto_intsink_in_sync_0,
  input auto_tile_reset_domain_tile_hartid_in,
  input auto_int_in_clock_xing_in_1_sync_0,
  input auto_int_in_clock_xing_in_0_sync_0,
  input auto_int_in_clock_xing_in_0_sync_1,
  input auto_tl_master_clock_xing_out_a_ready,
  output auto_tl_master_clock_xing_out_a_valid,
  output [2:0] auto_tl_master_clock_xing_out_a_bits_opcode,
  output [2:0] auto_tl_master_clock_xing_out_a_bits_param,
  output [3:0] auto_tl_master_clock_xing_out_a_bits_size,
  output [1:0] auto_tl_master_clock_xing_out_a_bits_source,
  output [31:0] auto_tl_master_clock_xing_out_a_bits_address,
  output [7:0] auto_tl_master_clock_xing_out_a_bits_mask,
  output [63:0] auto_tl_master_clock_xing_out_a_bits_data,
  output auto_tl_master_clock_xing_out_a_bits_corrupt,
  output auto_tl_master_clock_xing_out_b_ready,
  input auto_tl_master_clock_xing_out_b_valid,
  input [1:0] auto_tl_master_clock_xing_out_b_bits_param,
  input [31:0] auto_tl_master_clock_xing_out_b_bits_address,
  input auto_tl_master_clock_xing_out_c_ready,
  output auto_tl_master_clock_xing_out_c_valid,
  output [2:0] auto_tl_master_clock_xing_out_c_bits_opcode,
  output [2:0] auto_tl_master_clock_xing_out_c_bits_param,
  output [3:0] auto_tl_master_clock_xing_out_c_bits_size,
  output [1:0] auto_tl_master_clock_xing_out_c_bits_source,
  output [31:0] auto_tl_master_clock_xing_out_c_bits_address,
  output [63:0] auto_tl_master_clock_xing_out_c_bits_data,
  output auto_tl_master_clock_xing_out_c_bits_corrupt,
  output auto_tl_master_clock_xing_out_d_ready,
  input auto_tl_master_clock_xing_out_d_valid,
  input [2:0] auto_tl_master_clock_xing_out_d_bits_opcode,
  input [1:0] auto_tl_master_clock_xing_out_d_bits_param,
  input [3:0] auto_tl_master_clock_xing_out_d_bits_size,
  input [1:0] auto_tl_master_clock_xing_out_d_bits_source,
  input [1:0] auto_tl_master_clock_xing_out_d_bits_sink,
  input auto_tl_master_clock_xing_out_d_bits_denied,
  input [63:0] auto_tl_master_clock_xing_out_d_bits_data,
  input auto_tl_master_clock_xing_out_d_bits_corrupt,
  output auto_tl_master_clock_xing_out_e_valid,
  output [1:0] auto_tl_master_clock_xing_out_e_bits_sink,
  input auto_tap_clock_in_clock,
  input auto_tap_clock_in_reset) ; 
   wire _intsink_2_auto_out_0 ;  
   wire _intsink_1_auto_out_0 ;  
   wire _intsink_1_auto_out_1 ;  
   wire _intsink_auto_out_0 ;  
   wire _buffer_auto_in_a_ready ;  
   wire _buffer_auto_in_b_valid ;  
   wire [2:0] _buffer_auto_in_b_bits_opcode ;  
   wire [1:0] _buffer_auto_in_b_bits_param ;  
   wire [3:0] _buffer_auto_in_b_bits_size ;  
   wire [1:0] _buffer_auto_in_b_bits_source ;  
   wire [31:0] _buffer_auto_in_b_bits_address ;  
   wire [7:0] _buffer_auto_in_b_bits_mask ;  
   wire _buffer_auto_in_b_bits_corrupt ;  
   wire _buffer_auto_in_c_ready ;  
   wire _buffer_auto_in_d_valid ;  
   wire [2:0] _buffer_auto_in_d_bits_opcode ;  
   wire [1:0] _buffer_auto_in_d_bits_param ;  
   wire [3:0] _buffer_auto_in_d_bits_size ;  
   wire [1:0] _buffer_auto_in_d_bits_source ;  
   wire [1:0] _buffer_auto_in_d_bits_sink ;  
   wire _buffer_auto_in_d_bits_denied ;  
   wire [63:0] _buffer_auto_in_d_bits_data ;  
   wire _buffer_auto_in_d_bits_corrupt ;  
   wire _buffer_auto_in_e_ready ;  
   wire _tile_reset_domain_tile_auto_buffer_out_a_valid ;  
   wire [2:0] _tile_reset_domain_tile_auto_buffer_out_a_bits_opcode ;  
   wire [2:0] _tile_reset_domain_tile_auto_buffer_out_a_bits_param ;  
   wire [3:0] _tile_reset_domain_tile_auto_buffer_out_a_bits_size ;  
   wire [1:0] _tile_reset_domain_tile_auto_buffer_out_a_bits_source ;  
   wire [31:0] _tile_reset_domain_tile_auto_buffer_out_a_bits_address ;  
   wire [7:0] _tile_reset_domain_tile_auto_buffer_out_a_bits_mask ;  
   wire [63:0] _tile_reset_domain_tile_auto_buffer_out_a_bits_data ;  
   wire _tile_reset_domain_tile_auto_buffer_out_b_ready ;  
   wire _tile_reset_domain_tile_auto_buffer_out_c_valid ;  
   wire [2:0] _tile_reset_domain_tile_auto_buffer_out_c_bits_opcode ;  
   wire [2:0] _tile_reset_domain_tile_auto_buffer_out_c_bits_param ;  
   wire [3:0] _tile_reset_domain_tile_auto_buffer_out_c_bits_size ;  
   wire [1:0] _tile_reset_domain_tile_auto_buffer_out_c_bits_source ;  
   wire [31:0] _tile_reset_domain_tile_auto_buffer_out_c_bits_address ;  
   wire [63:0] _tile_reset_domain_tile_auto_buffer_out_c_bits_data ;  
   wire _tile_reset_domain_tile_auto_buffer_out_d_ready ;  
   wire _tile_reset_domain_tile_auto_buffer_out_e_valid ;  
   wire [1:0] _tile_reset_domain_tile_auto_buffer_out_e_bits_sink ;  
   wire _tile_reset_domain_tile_auto_wfi_out_0 ;  
  RocketTile tile_reset_domain_tile(.clock(auto_tap_clock_in_clock),.reset(auto_tap_clock_in_reset),.auto_buffer_out_a_ready(_buffer_auto_in_a_ready),.auto_buffer_out_a_valid(_tile_reset_domain_tile_auto_buffer_out_a_valid),.auto_buffer_out_a_bits_opcode(_tile_reset_domain_tile_auto_buffer_out_a_bits_opcode),.auto_buffer_out_a_bits_param(_tile_reset_domain_tile_auto_buffer_out_a_bits_param),.auto_buffer_out_a_bits_size(_tile_reset_domain_tile_auto_buffer_out_a_bits_size),.auto_buffer_out_a_bits_source(_tile_reset_domain_tile_auto_buffer_out_a_bits_source),.auto_buffer_out_a_bits_address(_tile_reset_domain_tile_auto_buffer_out_a_bits_address),.auto_buffer_out_a_bits_mask(_tile_reset_domain_tile_auto_buffer_out_a_bits_mask),.auto_buffer_out_a_bits_data(_tile_reset_domain_tile_auto_buffer_out_a_bits_data),.auto_buffer_out_b_ready(_tile_reset_domain_tile_auto_buffer_out_b_ready),.auto_buffer_out_b_valid(_buffer_auto_in_b_valid),.auto_buffer_out_b_bits_opcode(_buffer_auto_in_b_bits_opcode),.auto_buffer_out_b_bits_param(_buffer_auto_in_b_bits_param),.auto_buffer_out_b_bits_size(_buffer_auto_in_b_bits_size),.auto_buffer_out_b_bits_source(_buffer_auto_in_b_bits_source),.auto_buffer_out_b_bits_address(_buffer_auto_in_b_bits_address),.auto_buffer_out_b_bits_mask(_buffer_auto_in_b_bits_mask),.auto_buffer_out_b_bits_corrupt(_buffer_auto_in_b_bits_corrupt),.auto_buffer_out_c_ready(_buffer_auto_in_c_ready),.auto_buffer_out_c_valid(_tile_reset_domain_tile_auto_buffer_out_c_valid),.auto_buffer_out_c_bits_opcode(_tile_reset_domain_tile_auto_buffer_out_c_bits_opcode),.auto_buffer_out_c_bits_param(_tile_reset_domain_tile_auto_buffer_out_c_bits_param),.auto_buffer_out_c_bits_size(_tile_reset_domain_tile_auto_buffer_out_c_bits_size),.auto_buffer_out_c_bits_source(_tile_reset_domain_tile_auto_buffer_out_c_bits_source),.auto_buffer_out_c_bits_address(_tile_reset_domain_tile_auto_buffer_out_c_bits_address),.auto_buffer_out_c_bits_data(_tile_reset_domain_tile_auto_buffer_out_c_bits_data),.auto_buffer_out_d_ready(_tile_reset_domain_tile_auto_buffer_out_d_ready),.auto_buffer_out_d_valid(_buffer_auto_in_d_valid),.auto_buffer_out_d_bits_opcode(_buffer_auto_in_d_bits_opcode),.auto_buffer_out_d_bits_param(_buffer_auto_in_d_bits_param),.auto_buffer_out_d_bits_size(_buffer_auto_in_d_bits_size),.auto_buffer_out_d_bits_source(_buffer_auto_in_d_bits_source),.auto_buffer_out_d_bits_sink(_buffer_auto_in_d_bits_sink),.auto_buffer_out_d_bits_denied(_buffer_auto_in_d_bits_denied),.auto_buffer_out_d_bits_data(_buffer_auto_in_d_bits_data),.auto_buffer_out_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt),.auto_buffer_out_e_ready(_buffer_auto_in_e_ready),.auto_buffer_out_e_valid(_tile_reset_domain_tile_auto_buffer_out_e_valid),.auto_buffer_out_e_bits_sink(_tile_reset_domain_tile_auto_buffer_out_e_bits_sink),.auto_wfi_out_0(_tile_reset_domain_tile_auto_wfi_out_0),.auto_int_local_in_2_0(_intsink_2_auto_out_0),.auto_int_local_in_1_0(_intsink_1_auto_out_0),.auto_int_local_in_1_1(_intsink_1_auto_out_1),.auto_int_local_in_0_0(_intsink_auto_out_0),.auto_hartid_in(auto_tile_reset_domain_tile_hartid_in)); 
  TLBuffer_10 buffer(.clock(auto_tap_clock_in_clock),.reset(auto_tap_clock_in_reset),.auto_in_a_ready(_buffer_auto_in_a_ready),.auto_in_a_valid(_tile_reset_domain_tile_auto_buffer_out_a_valid),.auto_in_a_bits_opcode(_tile_reset_domain_tile_auto_buffer_out_a_bits_opcode),.auto_in_a_bits_param(_tile_reset_domain_tile_auto_buffer_out_a_bits_param),.auto_in_a_bits_size(_tile_reset_domain_tile_auto_buffer_out_a_bits_size),.auto_in_a_bits_source(_tile_reset_domain_tile_auto_buffer_out_a_bits_source),.auto_in_a_bits_address(_tile_reset_domain_tile_auto_buffer_out_a_bits_address),.auto_in_a_bits_mask(_tile_reset_domain_tile_auto_buffer_out_a_bits_mask),.auto_in_a_bits_data(_tile_reset_domain_tile_auto_buffer_out_a_bits_data),.auto_in_b_ready(_tile_reset_domain_tile_auto_buffer_out_b_ready),.auto_in_b_valid(_buffer_auto_in_b_valid),.auto_in_b_bits_opcode(_buffer_auto_in_b_bits_opcode),.auto_in_b_bits_param(_buffer_auto_in_b_bits_param),.auto_in_b_bits_size(_buffer_auto_in_b_bits_size),.auto_in_b_bits_source(_buffer_auto_in_b_bits_source),.auto_in_b_bits_address(_buffer_auto_in_b_bits_address),.auto_in_b_bits_mask(_buffer_auto_in_b_bits_mask),.auto_in_b_bits_corrupt(_buffer_auto_in_b_bits_corrupt),.auto_in_c_ready(_buffer_auto_in_c_ready),.auto_in_c_valid(_tile_reset_domain_tile_auto_buffer_out_c_valid),.auto_in_c_bits_opcode(_tile_reset_domain_tile_auto_buffer_out_c_bits_opcode),.auto_in_c_bits_param(_tile_reset_domain_tile_auto_buffer_out_c_bits_param),.auto_in_c_bits_size(_tile_reset_domain_tile_auto_buffer_out_c_bits_size),.auto_in_c_bits_source(_tile_reset_domain_tile_auto_buffer_out_c_bits_source),.auto_in_c_bits_address(_tile_reset_domain_tile_auto_buffer_out_c_bits_address),.auto_in_c_bits_data(_tile_reset_domain_tile_auto_buffer_out_c_bits_data),.auto_in_d_ready(_tile_reset_domain_tile_auto_buffer_out_d_ready),.auto_in_d_valid(_buffer_auto_in_d_valid),.auto_in_d_bits_opcode(_buffer_auto_in_d_bits_opcode),.auto_in_d_bits_param(_buffer_auto_in_d_bits_param),.auto_in_d_bits_size(_buffer_auto_in_d_bits_size),.auto_in_d_bits_source(_buffer_auto_in_d_bits_source),.auto_in_d_bits_sink(_buffer_auto_in_d_bits_sink),.auto_in_d_bits_denied(_buffer_auto_in_d_bits_denied),.auto_in_d_bits_data(_buffer_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt),.auto_in_e_ready(_buffer_auto_in_e_ready),.auto_in_e_valid(_tile_reset_domain_tile_auto_buffer_out_e_valid),.auto_in_e_bits_sink(_tile_reset_domain_tile_auto_buffer_out_e_bits_sink),.auto_out_a_ready(auto_tl_master_clock_xing_out_a_ready),.auto_out_a_valid(auto_tl_master_clock_xing_out_a_valid),.auto_out_a_bits_opcode(auto_tl_master_clock_xing_out_a_bits_opcode),.auto_out_a_bits_param(auto_tl_master_clock_xing_out_a_bits_param),.auto_out_a_bits_size(auto_tl_master_clock_xing_out_a_bits_size),.auto_out_a_bits_source(auto_tl_master_clock_xing_out_a_bits_source),.auto_out_a_bits_address(auto_tl_master_clock_xing_out_a_bits_address),.auto_out_a_bits_mask(auto_tl_master_clock_xing_out_a_bits_mask),.auto_out_a_bits_data(auto_tl_master_clock_xing_out_a_bits_data),.auto_out_a_bits_corrupt(auto_tl_master_clock_xing_out_a_bits_corrupt),.auto_out_b_ready(auto_tl_master_clock_xing_out_b_ready),.auto_out_b_valid(auto_tl_master_clock_xing_out_b_valid),.auto_out_b_bits_param(auto_tl_master_clock_xing_out_b_bits_param),.auto_out_b_bits_address(auto_tl_master_clock_xing_out_b_bits_address),.auto_out_c_ready(auto_tl_master_clock_xing_out_c_ready),.auto_out_c_valid(auto_tl_master_clock_xing_out_c_valid),.auto_out_c_bits_opcode(auto_tl_master_clock_xing_out_c_bits_opcode),.auto_out_c_bits_param(auto_tl_master_clock_xing_out_c_bits_param),.auto_out_c_bits_size(auto_tl_master_clock_xing_out_c_bits_size),.auto_out_c_bits_source(auto_tl_master_clock_xing_out_c_bits_source),.auto_out_c_bits_address(auto_tl_master_clock_xing_out_c_bits_address),.auto_out_c_bits_data(auto_tl_master_clock_xing_out_c_bits_data),.auto_out_c_bits_corrupt(auto_tl_master_clock_xing_out_c_bits_corrupt),.auto_out_d_ready(auto_tl_master_clock_xing_out_d_ready),.auto_out_d_valid(auto_tl_master_clock_xing_out_d_valid),.auto_out_d_bits_opcode(auto_tl_master_clock_xing_out_d_bits_opcode),.auto_out_d_bits_param(auto_tl_master_clock_xing_out_d_bits_param),.auto_out_d_bits_size(auto_tl_master_clock_xing_out_d_bits_size),.auto_out_d_bits_source(auto_tl_master_clock_xing_out_d_bits_source),.auto_out_d_bits_sink(auto_tl_master_clock_xing_out_d_bits_sink),.auto_out_d_bits_denied(auto_tl_master_clock_xing_out_d_bits_denied),.auto_out_d_bits_data(auto_tl_master_clock_xing_out_d_bits_data),.auto_out_d_bits_corrupt(auto_tl_master_clock_xing_out_d_bits_corrupt),.auto_out_e_valid(auto_tl_master_clock_xing_out_e_valid),.auto_out_e_bits_sink(auto_tl_master_clock_xing_out_e_bits_sink)); 
  IntSyncAsyncCrossingSink_1 intsink(.clock(auto_tap_clock_in_clock),.auto_in_sync_0(auto_intsink_in_sync_0),.auto_out_0(_intsink_auto_out_0)); 
  IntSyncSyncCrossingSink intsink_1(.auto_in_sync_0(auto_int_in_clock_xing_in_0_sync_0),.auto_in_sync_1(auto_int_in_clock_xing_in_0_sync_1),.auto_out_0(_intsink_1_auto_out_0),.auto_out_1(_intsink_1_auto_out_1)); 
  IntSyncSyncCrossingSink_1 intsink_2(.auto_in_sync_0(auto_int_in_clock_xing_in_1_sync_0),.auto_out_0(_intsink_2_auto_out_0)); 
  IntSyncCrossingSource_1 intsource_1(.clock(auto_tap_clock_in_clock),.reset(auto_tap_clock_in_reset),.auto_in_0(1'h0),.auto_out_sync_0()); 
  IntSyncCrossingSource_1 intsource_2(.clock(auto_tap_clock_in_clock),.reset(auto_tap_clock_in_reset),.auto_in_0(_tile_reset_domain_tile_auto_wfi_out_0),.auto_out_sync_0()); 
  IntSyncCrossingSource_1 intsource_3(.clock(auto_tap_clock_in_clock),.reset(auto_tap_clock_in_reset),.auto_in_0(1'h0),.auto_out_sync_0()); 
endmodule
 
module TLMonitor_26 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [1:0] io_in_a_bits_size,
  input [8:0] io_in_a_bits_source,
  input [27:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_size,
  input [8:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [1:0] size ;  
   reg [8:0] source ;  
   reg [27:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] size_1 ;  
   reg [8:0] source_1 ;  
   reg [303:0] inflight ;  
   reg [1215:0] inflight_opcodes ;  
   reg [1215:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire [1215:0] _GEN={1205'h0,io_in_d_bits_source,2'h0} ;  
   wire [1215:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire [511:0] _GEN_0={503'h0,io_in_a_bits_source} ;  
   wire _GEN_1=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   wire [511:0] _GEN_2={503'h0,io_in_d_bits_source} ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [303:0] inflight_1 ;  
   reg [1215:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire [5:0] _is_aligned_mask_T_1=6'h7<<io_in_a_bits_size ;  
   wire [2:0] _GEN_3=io_in_a_bits_address[2:0]&~(_is_aligned_mask_T_1[2:0]) ;  
   wire mask_size=io_in_a_bits_size==2'h2 ;  
   wire mask_acc=(&io_in_a_bits_size)|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=(&io_in_a_bits_size)|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_4=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_5=io_in_a_bits_source>9'h12F ;  
   wire _GEN_6=io_in_a_bits_param>3'h2 ;  
   wire _GEN_7=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_8=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_9=io_in_a_bits_source<9'h130 ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_11=io_in_a_bits_address[27:26]!=2'h3 ;  
   wire _GEN_12=io_in_a_bits_mask!=mask ;  
   wire _GEN_13=_GEN_9&~_GEN_11 ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_17=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_18=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_19=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_20=io_in_d_bits_source>9'h12F ;  
   wire _GEN_21=io_in_d_bits_size!=2'h3 ;  
   wire _GEN_22=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_23=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_24=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_25=io_in_d_valid&d_first_counter&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&~a_first_counter_1 ;  
   wire [511:0] _a_set_wo_ready_T=512'h1<<_GEN_0 ;  
   wire [303:0] a_set_wo_ready=_same_cycle_resp_T_1 ? _a_set_wo_ready_T[303:0]:304'h0 ;  
   wire _GEN_26=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_27=_GEN_26&~d_release_ack ;  
   wire same_cycle_resp=_same_cycle_resp_T_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [303:0] _GEN_28={295'h0,io_in_d_bits_source} ;  
   wire _GEN_29=_GEN_27&same_cycle_resp&~reset ;  
   wire _GEN_30=_GEN_27&~same_cycle_resp&~reset ;  
   wire [3:0] _GEN_31={2'h0,io_in_d_bits_size} ;  
   wire _GEN_32=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
   wire [303:0] _GEN_33=inflight>>io_in_a_bits_source ;  
   wire [303:0] _GEN_34=inflight>>_GEN_28 ;  
   wire [1215:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
   wire [511:0] _d_clr_wo_ready_T=512'h1<<_GEN_2 ;  
   wire [303:0] _GEN_35=inflight_1>>_GEN_28 ;  
   wire [1215:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|_GEN_3))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&~reset&_GEN_33[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~reset&~(_GEN_34[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_29&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_31!={1'h0,_a_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~a_first_counter_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_27 ? _d_clr_wo_ready_T[303:0]:304'h0)|a_set_wo_ready==304'h0))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==304'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&~(_GEN_35[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_32&_GEN_31!={1'h0,_c_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==304'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/Plic.scala:364:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [4110:0] _GEN_36={4100'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _d_clr_T=512'h1<<_GEN_2 ;  
   wire [511:0] _a_set_T=512'h1<<_GEN_0 ;  
   wire [4110:0] _d_opcodes_clr_T_5=4111'hF<<_GEN_36 ;  
   wire [4098:0] _a_opcodes_set_T_1={4095'h0,_GEN_1 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{4088'h0,io_in_a_bits_source,2'h0} ;  
   wire [4110:0] _d_sizes_clr_T_5=4111'hF<<_GEN_36 ;  
   wire [4097:0] _a_sizes_set_T_1={4095'h0,_GEN_1 ? {io_in_a_bits_size,1'h1}:3'h0}<<{4087'h0,io_in_a_bits_source,2'h0} ;  
   wire [511:0] _d_clr_T_1=512'h1<<_GEN_2 ;  
   wire [4110:0] _d_sizes_clr_T_11=4111'hF<<_GEN_36 ;  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_37=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire _GEN_38=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=304'h0;
              inflight_opcodes <=1216'h0;
              inflight_sizes <=1216'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=304'h0;
              inflight_sizes_1 <=1216'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|(_GEN_1 ? _a_set_T[303:0]:304'h0))&~(_GEN_37 ? _d_clr_T[303:0]:304'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_1 ? _a_opcodes_set_T_1[1215:0]:1216'h0))&~(_GEN_37 ? _d_opcodes_clr_T_5[1215:0]:1216'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_1 ? _a_sizes_set_T_1[1215:0]:1216'h0))&~(_GEN_37 ? _d_sizes_clr_T_5[1215:0]:1216'h0);
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_38 ? _d_clr_T_1[303:0]:304'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_38 ? _d_sizes_clr_T_11[1215:0]:1216'h0);
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module LevelGateway (
  input clock,
  input reset,
  input io_interrupt,
  output io_plic_valid,
  input io_plic_ready,
  input io_plic_complete) ; 
   reg inFlight ;  
  always @( posedge clock)
       begin 
         if (reset)
            inFlight <=1'h0;
          else 
            inFlight <=~io_plic_complete&(io_interrupt&io_plic_ready|inFlight);
       end
  
  assign io_plic_valid=io_interrupt&~inFlight; 
endmodule
 
module PLICFanIn (
  input [1:0] io_prio_0,
  input [1:0] io_prio_1,
  input [1:0] io_ip,
  output [1:0] io_dev,
  output [1:0] io_max) ; 
   wire [2:0] effectivePriority_1={io_ip[0],io_prio_0} ;  
   wire _GEN=effectivePriority_1<3'h5 ;  
   wire [2:0] _GEN_0=_GEN ? 3'h4:effectivePriority_1 ;  
   wire _GEN_1=_GEN_0>={io_ip[1],io_prio_1} ;  
  assign io_dev=_GEN_1 ? {1'h0,~_GEN}:2'h2; 
  assign io_max=_GEN_1 ? _GEN_0[1:0]:io_prio_1; 
endmodule
 
module Queue_83 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input io_enq_bits_read,
  input [22:0] io_enq_bits_index,
  input [63:0] io_enq_bits_data,
  input [7:0] io_enq_bits_mask,
  input [8:0] io_enq_bits_extra_tlrr_extra_source,
  input [1:0] io_enq_bits_extra_tlrr_extra_size,
  input io_deq_ready,
  output io_deq_valid,
  output io_deq_bits_read,
  output [22:0] io_deq_bits_index,
  output [63:0] io_deq_bits_data,
  output [7:0] io_deq_bits_mask,
  output [8:0] io_deq_bits_extra_tlrr_extra_source,
  output [1:0] io_deq_bits_extra_tlrr_extra_size) ; 
   reg [106:0] ram ;  
   reg full ;  
   wire do_enq=~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            ram <={io_enq_bits_extra_tlrr_extra_size,io_enq_bits_extra_tlrr_extra_source,io_enq_bits_mask,io_enq_bits_data,io_enq_bits_index,io_enq_bits_read};
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(io_deq_ready&full)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=full; 
  assign io_deq_bits_read=ram[0]; 
  assign io_deq_bits_index=ram[23:1]; 
  assign io_deq_bits_data=ram[87:24]; 
  assign io_deq_bits_mask=ram[95:88]; 
  assign io_deq_bits_extra_tlrr_extra_source=ram[104:96]; 
  assign io_deq_bits_extra_tlrr_extra_size=ram[106:105]; 
endmodule
 
module TLPLIC (
  input clock,
  input reset,
  input auto_int_in_0,
  input auto_int_in_1,
  output auto_int_out_0,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [1:0] auto_in_a_bits_size,
  input [8:0] auto_in_a_bits_source,
  input [27:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_size,
  output [8:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data) ; 
   wire out_woready_6 ;  
   wire _out_wofireMux_T ;  
   wire out_backSel_8 ;  
   wire completer_0 ;  
   wire [1:0] completerDev ;  
   wire _out_back_q_io_enq_ready ;  
   wire _out_back_q_io_deq_valid ;  
   wire _out_back_q_io_deq_bits_read ;  
   wire [22:0] _out_back_q_io_deq_bits_index ;  
   wire [63:0] _out_back_q_io_deq_bits_data ;  
   wire [7:0] _out_back_q_io_deq_bits_mask ;  
   wire [8:0] _out_back_q_io_deq_bits_extra_tlrr_extra_source ;  
   wire [1:0] _out_back_q_io_deq_bits_extra_tlrr_extra_size ;  
   wire [1:0] _fanin_io_dev ;  
   wire [1:0] _fanin_io_max ;  
   wire _gateways_gateway_1_io_plic_valid ;  
   wire _gateways_gateway_io_plic_valid ;  
   reg [1:0] priority_0 ;  
   reg [1:0] priority_1 ;  
   reg [1:0] threshold_0 ;  
   reg pending_0 ;  
   reg pending_1 ;  
   reg [1:0] enables_0_0 ;  
   reg [1:0] maxDevs_0 ;  
   reg [1:0] intnodeOut_0_REG ;  
   wire [3:0] _completedDevs_T=4'h1<<completerDev ;  
   wire [1:0] completedDevs=completer_0 ? _completedDevs_T[2:1]:2'h0 ;  
   wire _out_T_9={_out_back_q_io_deq_bits_index[22:19],_out_back_q_io_deq_bits_index[17:11],_out_back_q_io_deq_bits_index[8:1]}==19'h0 ;  
   wire [31:0] _out_womask_T_6={{8{_out_back_q_io_deq_bits_mask[7]}},{8{_out_back_q_io_deq_bits_mask[6]}},{8{_out_back_q_io_deq_bits_mask[5]}},{8{_out_back_q_io_deq_bits_mask[4]}}} ;  
   wire claimer_0=_out_wofireMux_T&_out_back_q_io_deq_bits_read&out_backSel_8&_out_T_9&(|_out_womask_T_6) ;  
  assign completerDev=_out_back_q_io_deq_bits_data[33:32]; 
  always @( posedge clock)
       begin 
         if (~reset&claimer_0&claimer_0-1'h1)
            begin 
              if (1)$display("Assertion failed\n    at Plic.scala:246 assert((claimer.asUInt & (claimer.asUInt - 1.U)) === 0.U) // One-Hot\n");
              if (1)$display("");
            end 
         if (~reset&completer_0&completer_0-1'h1)
            begin 
              if (1)$display("Assertion failed\n    at Plic.scala:263 assert((completer.asUInt & (completer.asUInt - 1.U)) === 0.U) // One-Hot\n");
              if (1)$display("");
            end 
       end
  
   wire [2:0] _out_completer_0_T={enables_0_0,1'h0}>>completerDev ;  
  assign completer_0=out_woready_6&(&_out_womask_T_6)&_out_completer_0_T[0]; 
   wire [3:0] out_oindex={_out_back_q_io_deq_bits_index[18],_out_back_q_io_deq_bits_index[10:9],_out_back_q_io_deq_bits_index[0]} ;  
   wire [3:0] _GEN={_out_back_q_io_deq_bits_index[18],_out_back_q_io_deq_bits_index[10:9],_out_back_q_io_deq_bits_index[0]} ;  
  assign out_backSel_8=_GEN==4'h8; 
  assign _out_wofireMux_T=_out_back_q_io_deq_valid&auto_in_d_ready; 
   wire _out_wofireMux_T_2=_out_wofireMux_T&~_out_back_q_io_deq_bits_read ;  
  assign out_woready_6=_out_wofireMux_T_2&out_backSel_8&_out_T_9; 
   wire _out_out_bits_data_T_5=out_oindex==4'h0 ;  
   wire [2:0] nodeIn_d_bits_opcode={2'h0,_out_back_q_io_deq_bits_read} ;  
   wire [1:0] claiming=claimer_0 ? maxDevs_0:2'h0 ;  
   wire claimedDevs_1=claiming==2'h1 ;  
   wire claimedDevs_2=claiming==2'h2 ;  
  always @( posedge clock)
       begin 
         if (_out_wofireMux_T_2&_GEN==4'h0&_out_T_9&_out_back_q_io_deq_bits_mask[4])
            priority_0 <=_out_back_q_io_deq_bits_data[33:32];
         if (_out_wofireMux_T_2&_GEN==4'h1&_out_T_9&_out_back_q_io_deq_bits_mask[0])
            priority_1 <=_out_back_q_io_deq_bits_data[1:0];
         if (out_woready_6&_out_back_q_io_deq_bits_mask[0])
            threshold_0 <=_out_back_q_io_deq_bits_data[1:0];
         if (_out_wofireMux_T_2&_GEN==4'h4&_out_T_9&_out_back_q_io_deq_bits_mask[0])
            enables_0_0 <=_out_back_q_io_deq_bits_data[2:1];
         maxDevs_0 <=_fanin_io_dev;
         intnodeOut_0_REG <=_fanin_io_max;
         if (reset)
            begin 
              pending_0 <=1'h0;
              pending_1 <=1'h0;
            end 
          else 
            begin 
              if (claimedDevs_1|_gateways_gateway_io_plic_valid)
                 pending_0 <=~claimedDevs_1;
              if (claimedDevs_2|_gateways_gateway_1_io_plic_valid)
                 pending_1 <=~claimedDevs_2;
            end 
       end
  
  TLMonitor_26 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_out_back_q_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(_out_back_q_io_deq_valid),.io_in_d_bits_opcode(nodeIn_d_bits_opcode),.io_in_d_bits_size(_out_back_q_io_deq_bits_extra_tlrr_extra_size),.io_in_d_bits_source(_out_back_q_io_deq_bits_extra_tlrr_extra_source)); 
  LevelGateway gateways_gateway(.clock(clock),.reset(reset),.io_interrupt(auto_int_in_0),.io_plic_valid(_gateways_gateway_io_plic_valid),.io_plic_ready(~pending_0),.io_plic_complete(completedDevs[0])); 
  LevelGateway gateways_gateway_1(.clock(clock),.reset(reset),.io_interrupt(auto_int_in_1),.io_plic_valid(_gateways_gateway_1_io_plic_valid),.io_plic_ready(~pending_1),.io_plic_complete(completedDevs[1])); 
  PLICFanIn fanin(.io_prio_0(priority_0),.io_prio_1(priority_1),.io_ip(enables_0_0&{pending_1,pending_0}),.io_dev(_fanin_io_dev),.io_max(_fanin_io_max)); 
  Queue_83 out_back_q(.clock(clock),.reset(reset),.io_enq_ready(_out_back_q_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_read(auto_in_a_bits_opcode==3'h4),.io_enq_bits_index(auto_in_a_bits_address[25:3]),.io_enq_bits_data(auto_in_a_bits_data),.io_enq_bits_mask(auto_in_a_bits_mask),.io_enq_bits_extra_tlrr_extra_source(auto_in_a_bits_source),.io_enq_bits_extra_tlrr_extra_size(auto_in_a_bits_size),.io_deq_ready(auto_in_d_ready),.io_deq_valid(_out_back_q_io_deq_valid),.io_deq_bits_read(_out_back_q_io_deq_bits_read),.io_deq_bits_index(_out_back_q_io_deq_bits_index),.io_deq_bits_data(_out_back_q_io_deq_bits_data),.io_deq_bits_mask(_out_back_q_io_deq_bits_mask),.io_deq_bits_extra_tlrr_extra_source(_out_back_q_io_deq_bits_extra_tlrr_extra_source),.io_deq_bits_extra_tlrr_extra_size(_out_back_q_io_deq_bits_extra_tlrr_extra_size)); 
  assign auto_int_out_0=intnodeOut_0_REG>threshold_0; 
  assign auto_in_a_ready=_out_back_q_io_enq_ready; 
  assign auto_in_d_valid=_out_back_q_io_deq_valid; 
  assign auto_in_d_bits_opcode=nodeIn_d_bits_opcode; 
  assign auto_in_d_bits_size=_out_back_q_io_deq_bits_extra_tlrr_extra_size; 
  assign auto_in_d_bits_source=_out_back_q_io_deq_bits_extra_tlrr_extra_source; 
  assign auto_in_d_bits_data=~(_out_out_bits_data_T_5|out_oindex==4'h1|out_oindex==4'h2|out_oindex==4'h4|out_oindex==4'h8)|_out_T_9 ? (_out_out_bits_data_T_5 ? {30'h0,priority_0,32'h0}:out_oindex==4'h1 ? {62'h0,priority_1}:out_oindex==4'h2 ? {61'h0,pending_1,pending_0,1'h0}:out_oindex==4'h4 ? {61'h0,enables_0_0,1'h0}:out_oindex==4'h8 ? {30'h0,maxDevs_0,30'h0,threshold_0}:64'h0):64'h0; 
endmodule
 
module ClockSinkDomain (
  input auto_plic_int_in_0,
  input auto_plic_int_in_1,
  output auto_plic_int_out_0,
  output auto_plic_in_a_ready,
  input auto_plic_in_a_valid,
  input [2:0] auto_plic_in_a_bits_opcode,
  input [2:0] auto_plic_in_a_bits_param,
  input [1:0] auto_plic_in_a_bits_size,
  input [8:0] auto_plic_in_a_bits_source,
  input [27:0] auto_plic_in_a_bits_address,
  input [7:0] auto_plic_in_a_bits_mask,
  input [63:0] auto_plic_in_a_bits_data,
  input auto_plic_in_a_bits_corrupt,
  input auto_plic_in_d_ready,
  output auto_plic_in_d_valid,
  output [2:0] auto_plic_in_d_bits_opcode,
  output [1:0] auto_plic_in_d_bits_size,
  output [8:0] auto_plic_in_d_bits_source,
  output [63:0] auto_plic_in_d_bits_data,
  input auto_clock_in_clock,
  input auto_clock_in_reset) ; 
  TLPLIC plic(.clock(auto_clock_in_clock),.reset(auto_clock_in_reset),.auto_int_in_0(auto_plic_int_in_0),.auto_int_in_1(auto_plic_int_in_1),.auto_int_out_0(auto_plic_int_out_0),.auto_in_a_ready(auto_plic_in_a_ready),.auto_in_a_valid(auto_plic_in_a_valid),.auto_in_a_bits_opcode(auto_plic_in_a_bits_opcode),.auto_in_a_bits_param(auto_plic_in_a_bits_param),.auto_in_a_bits_size(auto_plic_in_a_bits_size),.auto_in_a_bits_source(auto_plic_in_a_bits_source),.auto_in_a_bits_address(auto_plic_in_a_bits_address),.auto_in_a_bits_mask(auto_plic_in_a_bits_mask),.auto_in_a_bits_data(auto_plic_in_a_bits_data),.auto_in_a_bits_corrupt(auto_plic_in_a_bits_corrupt),.auto_in_d_ready(auto_plic_in_d_ready),.auto_in_d_valid(auto_plic_in_d_valid),.auto_in_d_bits_opcode(auto_plic_in_d_bits_opcode),.auto_in_d_bits_size(auto_plic_in_d_bits_size),.auto_in_d_bits_source(auto_plic_in_d_bits_source),.auto_in_d_bits_data(auto_plic_in_d_bits_data)); 
endmodule
 
module TLMonitor_27 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [1:0] io_in_a_bits_size,
  input [8:0] io_in_a_bits_source,
  input [25:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_size,
  input [8:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [1:0] size ;  
   reg [8:0] source ;  
   reg [25:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] size_1 ;  
   reg [8:0] source_1 ;  
   reg [303:0] inflight ;  
   reg [1215:0] inflight_opcodes ;  
   reg [1215:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire [1215:0] _GEN={1205'h0,io_in_d_bits_source,2'h0} ;  
   wire [1215:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire _GEN_0=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [303:0] inflight_1 ;  
   reg [1215:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire [5:0] _is_aligned_mask_T_1=6'h7<<io_in_a_bits_size ;  
   wire [2:0] _GEN_1=io_in_a_bits_address[2:0]&~(_is_aligned_mask_T_1[2:0]) ;  
   wire mask_size=io_in_a_bits_size==2'h2 ;  
   wire mask_acc=(&io_in_a_bits_size)|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=(&io_in_a_bits_size)|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_3=io_in_a_bits_source>9'h12F ;  
   wire _GEN_4=io_in_a_bits_param>3'h2 ;  
   wire _GEN_5=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_6=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_7=io_in_a_bits_source<9'h130 ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_9=io_in_a_bits_address[25:16]!=10'h200 ;  
   wire _GEN_10=io_in_a_bits_mask!=mask ;  
   wire _GEN_11=_GEN_7&~_GEN_9 ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_16=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_18=io_in_d_bits_source>9'h12F ;  
   wire _GEN_19=io_in_d_bits_size!=2'h3 ;  
   wire _GEN_20=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_21=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_22=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_23=io_in_d_valid&d_first_counter&~reset ;  
   wire _GEN_24=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_25=_GEN_24&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&~a_first_counter_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [303:0] _GEN_26={295'h0,io_in_d_bits_source} ;  
   wire _GEN_27=_GEN_25&same_cycle_resp&~reset ;  
   wire _GEN_28=_GEN_25&~same_cycle_resp&~reset ;  
   wire [3:0] _GEN_29={2'h0,io_in_d_bits_size} ;  
   wire _GEN_30=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
   wire [303:0] _GEN_31=inflight>>io_in_a_bits_source ;  
   wire [303:0] _GEN_32=inflight>>_GEN_26 ;  
   wire [1215:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
   wire [303:0] _GEN_33=inflight_1>>_GEN_26 ;  
   wire [1215:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&_GEN_19)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&_GEN_31[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~reset&~(_GEN_32[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_28&_GEN_29!={1'h0,_a_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~a_first_counter_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==304'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&~(_GEN_33[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_30&_GEN_29!={1'h0,_c_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==304'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/CLINT.scala:108:16)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [511:0] _GEN_34={503'h0,io_in_d_bits_source} ;  
   wire [4110:0] _GEN_35={4100'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _d_clr_T=512'h1<<_GEN_34 ;  
   wire [511:0] _a_set_T=512'h1<<io_in_a_bits_source ;  
   wire [4110:0] _d_opcodes_clr_T_5=4111'hF<<_GEN_35 ;  
   wire [4098:0] _a_opcodes_set_T_1={4095'h0,_GEN_0 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{4088'h0,io_in_a_bits_source,2'h0} ;  
   wire [4110:0] _d_sizes_clr_T_5=4111'hF<<_GEN_35 ;  
   wire [4097:0] _a_sizes_set_T_1={4095'h0,_GEN_0 ? {io_in_a_bits_size,1'h1}:3'h0}<<{4087'h0,io_in_a_bits_source,2'h0} ;  
   wire [511:0] _d_clr_T_1=512'h1<<_GEN_34 ;  
   wire [4110:0] _d_sizes_clr_T_11=4111'hF<<_GEN_35 ;  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_36=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire _GEN_37=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=304'h0;
              inflight_opcodes <=1216'h0;
              inflight_sizes <=1216'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=304'h0;
              inflight_sizes_1 <=1216'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|(_GEN_0 ? _a_set_T[303:0]:304'h0))&~(_GEN_36 ? _d_clr_T[303:0]:304'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_0 ? _a_opcodes_set_T_1[1215:0]:1216'h0))&~(_GEN_36 ? _d_opcodes_clr_T_5[1215:0]:1216'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_0 ? _a_sizes_set_T_1[1215:0]:1216'h0))&~(_GEN_36 ? _d_sizes_clr_T_5[1215:0]:1216'h0);
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_37 ? _d_clr_T_1[303:0]:304'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_37 ? _d_sizes_clr_T_11[1215:0]:1216'h0);
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module CLINT (
  input clock,
  input reset,
  output auto_int_out_0,
  output auto_int_out_1,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [1:0] auto_in_a_bits_size,
  input [8:0] auto_in_a_bits_source,
  input [25:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input [63:0] auto_in_a_bits_data,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_size,
  output [8:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data,
  input io_rtcTick) ; 
   wire out_woready_9 ;  
   wire out_woready_17 ;  
   reg [63:0] time_0 ;  
   reg [63:0] pad ;  
   reg ipi_0 ;  
   wire in_bits_read=auto_in_a_bits_opcode==3'h4 ;  
   wire _out_T_5=auto_in_a_bits_address[13:3]==11'h0 ;  
   wire valids_1_0=out_woready_9&auto_in_a_bits_mask[0] ;  
   wire valids_1_1=out_woready_9&auto_in_a_bits_mask[1] ;  
   wire valids_1_2=out_woready_9&auto_in_a_bits_mask[2] ;  
   wire valids_1_3=out_woready_9&auto_in_a_bits_mask[3] ;  
   wire valids_1_4=out_woready_9&auto_in_a_bits_mask[4] ;  
   wire valids_1_5=out_woready_9&auto_in_a_bits_mask[5] ;  
   wire valids_1_6=out_woready_9&auto_in_a_bits_mask[6] ;  
   wire valids_1_7=out_woready_9&auto_in_a_bits_mask[7] ;  
   wire valids_0=out_woready_17&auto_in_a_bits_mask[0] ;  
   wire valids_1=out_woready_17&auto_in_a_bits_mask[1] ;  
   wire valids_2=out_woready_17&auto_in_a_bits_mask[2] ;  
   wire valids_3=out_woready_17&auto_in_a_bits_mask[3] ;  
   wire valids_4=out_woready_17&auto_in_a_bits_mask[4] ;  
   wire valids_5=out_woready_17&auto_in_a_bits_mask[5] ;  
   wire valids_6=out_woready_17&auto_in_a_bits_mask[6] ;  
   wire valids_7=out_woready_17&auto_in_a_bits_mask[7] ;  
   wire _out_wofireMux_T_2=auto_in_a_valid&auto_in_d_ready&~in_bits_read ;  
  assign out_woready_17=_out_wofireMux_T_2&auto_in_a_bits_address[15:14]==2'h1&_out_T_5; 
  assign out_woready_9=_out_wofireMux_T_2&auto_in_a_bits_address[15:14]==2'h2&(&(auto_in_a_bits_address[13:3])); 
   reg casez_tmp ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_address[15:14])
          2 'b00:
             casez_tmp =_out_T_5;
          2 'b01:
             casez_tmp =_out_T_5;
          2 'b10:
             casez_tmp =&(auto_in_a_bits_address[13:3]);
          default :
             casez_tmp =1'h1;
         endcase 
       end
  
   reg [63:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_address[15:14])
          2 'b00:
             casez_tmp_0 ={63'h0,ipi_0};
          2 'b01:
             casez_tmp_0 =pad;
          2 'b10:
             casez_tmp_0 =time_0;
          default :
             casez_tmp_0 =64'h0;
         endcase 
       end
  
   wire [2:0] nodeIn_d_bits_opcode={2'h0,in_bits_read} ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              time_0 <=64'h0;
              ipi_0 <=1'h0;
            end 
          else 
            begin 
              if (valids_1_0|valids_1_1|valids_1_2|valids_1_3|valids_1_4|valids_1_5|valids_1_6|valids_1_7)
                 time_0 <={valids_1_7 ? auto_in_a_bits_data[63:56]:time_0[63:56],valids_1_6 ? auto_in_a_bits_data[55:48]:time_0[55:48],valids_1_5 ? auto_in_a_bits_data[47:40]:time_0[47:40],valids_1_4 ? auto_in_a_bits_data[39:32]:time_0[39:32],valids_1_3 ? auto_in_a_bits_data[31:24]:time_0[31:24],valids_1_2 ? auto_in_a_bits_data[23:16]:time_0[23:16],valids_1_1 ? auto_in_a_bits_data[15:8]:time_0[15:8],valids_1_0 ? auto_in_a_bits_data[7:0]:time_0[7:0]};
               else 
                 if (io_rtcTick)
                    time_0 <=time_0+64'h1;
              if (_out_wofireMux_T_2&auto_in_a_bits_address[15:14]==2'h0&_out_T_5&auto_in_a_bits_mask[0])
                 ipi_0 <=auto_in_a_bits_data[0];
            end 
         if (valids_0|valids_1|valids_2|valids_3|valids_4|valids_5|valids_6|valids_7)
            pad <={valids_7 ? auto_in_a_bits_data[63:56]:pad[63:56],valids_6 ? auto_in_a_bits_data[55:48]:pad[55:48],valids_5 ? auto_in_a_bits_data[47:40]:pad[47:40],valids_4 ? auto_in_a_bits_data[39:32]:pad[39:32],valids_3 ? auto_in_a_bits_data[31:24]:pad[31:24],valids_2 ? auto_in_a_bits_data[23:16]:pad[23:16],valids_1 ? auto_in_a_bits_data[15:8]:pad[15:8],valids_0 ? auto_in_a_bits_data[7:0]:pad[7:0]};
       end
  
  TLMonitor_27 monitor(.clock(clock),.reset(reset),.io_in_a_ready(auto_in_d_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_in_a_valid),.io_in_d_bits_opcode(nodeIn_d_bits_opcode),.io_in_d_bits_size(auto_in_a_bits_size),.io_in_d_bits_source(auto_in_a_bits_source)); 
  assign auto_int_out_0=ipi_0; 
  assign auto_int_out_1=time_0>=pad; 
  assign auto_in_a_ready=auto_in_d_ready; 
  assign auto_in_d_valid=auto_in_a_valid; 
  assign auto_in_d_bits_opcode=nodeIn_d_bits_opcode; 
  assign auto_in_d_bits_size=auto_in_a_bits_size; 
  assign auto_in_d_bits_source=auto_in_a_bits_source; 
  assign auto_in_d_bits_data=casez_tmp ? casez_tmp_0:64'h0; 
endmodule
 
module BundleBridgeNexus_15 (
  output auto_out) ; 
   wire outputs_0=1'h0 ;  
  assign auto_out=outputs_0; 
endmodule
 
module TLMonitor_28 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [8:0] io_in_a_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [1:0] io_in_d_bits_size,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [8:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [1:0] size_1 ;  
   reg sink ;  
   reg denied ;  
   reg inflight ;  
   reg [3:0] inflight_opcodes ;  
   reg [3:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire a_set=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg inflight_1 ;  
   reg [3:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire _GEN=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_0=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_1=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_3=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_4=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_5=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_7=io_in_d_bits_param==2'h2 ;  
   wire _GEN_8=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_9=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_10=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_11=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_12=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_13=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_14=io_in_d_valid&d_first_counter&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&~a_first_counter_1 ;  
   wire _GEN_15=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_16=_GEN_15&~d_release_ack ;  
   wire _GEN_17=_GEN_16&_same_cycle_resp_T_1&~reset ;  
   wire _GEN_18=_GEN_16&~_same_cycle_resp_T_1&~reset ;  
   wire [3:0] _GEN_19={2'h0,io_in_d_bits_size} ;  
   wire _GEN_20=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
  always @( posedge clock)
       begin 
         if (_GEN)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (a_set&~reset&inflight)
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~reset&~(inflight|_same_cycle_resp_T_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_size!=2'h2)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_19!={1'h0,inflight_sizes[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&~a_first_counter_1&io_in_a_valid&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~inflight_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&_GEN_19!={1'h0,inflight_sizes_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight_1|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:674:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire d_clr=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire [3:0] d_sizes_clr={4{d_clr}} ;  
   wire d_clr_1=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=1'h0;
              inflight_opcodes <=4'h0;
              inflight_sizes <=4'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=1'h0;
              inflight_sizes_1 <=4'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|a_set)&~d_clr;
              inflight_opcodes <=(inflight_opcodes|(a_set ? {io_in_a_bits_opcode,1'h1}:4'h0))&~d_sizes_clr;
              inflight_sizes <=(inflight_sizes|(a_set ? {1'h0,a_set ? 3'h5:3'h0}:4'h0))&~d_sizes_clr;
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~d_clr_1;
              inflight_sizes_1 <=inflight_sizes_1&~{4{d_clr_1}};
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLXbar_10 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [8:0] auto_in_a_bits_address,
  input [31:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output auto_in_d_bits_denied,
  output [31:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_1_a_ready,
  output auto_out_1_a_valid,
  output [2:0] auto_out_1_a_bits_opcode,
  output [6:0] auto_out_1_a_bits_address,
  output [31:0] auto_out_1_a_bits_data,
  output auto_out_1_d_ready,
  input auto_out_1_d_valid,
  input [2:0] auto_out_1_d_bits_opcode,
  input [31:0] auto_out_1_d_bits_data,
  input auto_out_0_a_ready,
  output auto_out_0_a_valid,
  output [2:0] auto_out_0_a_bits_opcode,
  output [8:0] auto_out_0_a_bits_address,
  output [31:0] auto_out_0_a_bits_data,
  output auto_out_0_d_ready,
  input auto_out_0_d_valid,
  input [2:0] auto_out_0_d_bits_opcode,
  input [1:0] auto_out_0_d_bits_param,
  input [1:0] auto_out_0_d_bits_size,
  input auto_out_0_d_bits_sink,
  input auto_out_0_d_bits_denied,
  input [31:0] auto_out_0_d_bits_data,
  input auto_out_0_d_bits_corrupt) ; 
   wire [4:0] _GEN=auto_in_a_bits_address[6:2]^5'h11 ;  
   wire requestAIO_0_0=auto_in_a_bits_address[8:6]==3'h0|{auto_in_a_bits_address[8:7],_GEN[4:2],_GEN[0]}==6'h0|{auto_in_a_bits_address[8:7],auto_in_a_bits_address[6:3]^4'hB}==6'h0|{auto_in_a_bits_address[8:7],~(auto_in_a_bits_address[6:5])}==4'h0|{auto_in_a_bits_address[8],~(auto_in_a_bits_address[7])}==2'h0|auto_in_a_bits_address[8] ;  
   wire requestAIO_0_1={auto_in_a_bits_address[8:7],auto_in_a_bits_address[6:4]^3'h4,auto_in_a_bits_address[2]}==6'h0|{auto_in_a_bits_address[8:7],auto_in_a_bits_address[6:3]^4'hA}==6'h0 ;  
   wire _portsAOI_in_0_a_ready_T_2=requestAIO_0_0&auto_out_0_a_ready|requestAIO_0_1&auto_out_1_a_ready ;  
   reg beatsLeft ;  
   wire [1:0] readys_valid={auto_out_1_d_valid,auto_out_0_d_valid} ;  
   reg [1:0] readys_mask ;  
   wire [1:0] _readys_filter_T_1=readys_valid&~readys_mask ;  
   wire [1:0] readys_readys=~({readys_mask[1],_readys_filter_T_1[1]|readys_mask[0]}&({_readys_filter_T_1[0],auto_out_1_d_valid}|_readys_filter_T_1)) ;  
   wire winner_0=readys_readys[0]&auto_out_0_d_valid ;  
   wire winner_1=readys_readys[1]&auto_out_1_d_valid ;  
   wire _in_0_d_valid_T=auto_out_0_d_valid|auto_out_1_d_valid ;  
  always @( posedge clock)
       begin 
         if (~reset&~(~winner_0|~winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
              if (1)$display("");
            end 
         if (~reset&~(~_in_0_d_valid_T|winner_0|winner_1))
            begin 
              if (1)$display("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
              if (1)$display("");
            end 
       end
  
   reg state_0 ;  
   reg state_1 ;  
   wire muxState_0=beatsLeft ? state_0:winner_0 ;  
   wire muxState_1=beatsLeft ? state_1:winner_1 ;  
   wire in_0_d_valid=beatsLeft ? state_0&auto_out_0_d_valid|state_1&auto_out_1_d_valid:_in_0_d_valid_T ;  
   wire _in_0_d_bits_T=muxState_0&auto_out_0_d_bits_corrupt ;  
   wire _in_0_d_bits_T_6=muxState_0&auto_out_0_d_bits_denied ;  
   wire [1:0] _readys_mask_T=readys_readys&readys_valid ;  
   wire latch=~beatsLeft&auto_in_d_ready ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              beatsLeft <=1'h0;
              readys_mask <=2'h3;
              state_0 <=1'h0;
              state_1 <=1'h0;
            end 
          else 
            begin 
              beatsLeft <=~latch&beatsLeft-(auto_in_d_ready&in_0_d_valid);
              if (latch&(|readys_valid))
                 readys_mask <=_readys_mask_T|{_readys_mask_T[0],1'h0};
              if (beatsLeft)
                 begin 
                 end 
               else 
                 begin 
                   state_0 <=winner_0;
                   state_1 <=winner_1;
                 end 
            end 
       end
  
  TLMonitor_28 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_portsAOI_in_0_a_ready_T_2),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(in_0_d_valid),.io_in_d_bits_opcode((muxState_0 ? auto_out_0_d_bits_opcode:3'h0)|(muxState_1 ? auto_out_1_d_bits_opcode:3'h0)),.io_in_d_bits_param(muxState_0 ? auto_out_0_d_bits_param:2'h0),.io_in_d_bits_size((muxState_0 ? auto_out_0_d_bits_size:2'h0)|{muxState_1,1'h0}),.io_in_d_bits_sink(muxState_0&auto_out_0_d_bits_sink),.io_in_d_bits_denied(_in_0_d_bits_T_6),.io_in_d_bits_corrupt(_in_0_d_bits_T)); 
  assign auto_in_a_ready=_portsAOI_in_0_a_ready_T_2; 
  assign auto_in_d_valid=in_0_d_valid; 
  assign auto_in_d_bits_denied=_in_0_d_bits_T_6; 
  assign auto_in_d_bits_data=(muxState_0 ? auto_out_0_d_bits_data:32'h0)|(muxState_1 ? auto_out_1_d_bits_data:32'h0); 
  assign auto_in_d_bits_corrupt=_in_0_d_bits_T; 
  assign auto_out_1_a_valid=auto_in_a_valid&requestAIO_0_1; 
  assign auto_out_1_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_1_a_bits_address=auto_in_a_bits_address[6:0]; 
  assign auto_out_1_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_1_d_ready=auto_in_d_ready&(beatsLeft ? state_1:readys_readys[1]); 
  assign auto_out_0_a_valid=auto_in_a_valid&requestAIO_0_0; 
  assign auto_out_0_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_0_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_0_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_0_d_ready=auto_in_d_ready&(beatsLeft ? state_0:readys_readys[0]); 
endmodule
 
module DMIToTL (
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [8:0] auto_out_a_bits_address,
  output [31:0] auto_out_a_bits_data,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input auto_out_d_bits_denied,
  input [31:0] auto_out_d_bits_data,
  input auto_out_d_bits_corrupt,
  output io_dmi_req_ready,
  input io_dmi_req_valid,
  input [6:0] io_dmi_req_bits_addr,
  input [31:0] io_dmi_req_bits_data,
  input [1:0] io_dmi_req_bits_op,
  input io_dmi_resp_ready,
  output io_dmi_resp_valid,
  output [31:0] io_dmi_resp_bits_data,
  output [1:0] io_dmi_resp_bits_resp) ; 
   wire _GEN=io_dmi_req_bits_op==2'h2 ;  
   wire _GEN_0=io_dmi_req_bits_op==2'h1 ;  
  assign auto_out_a_valid=io_dmi_req_valid; 
  assign auto_out_a_bits_opcode=_GEN ? 3'h0:{_GEN_0,2'h0}; 
  assign auto_out_a_bits_address=_GEN|_GEN_0 ? {io_dmi_req_bits_addr,2'h0}:9'h48; 
  assign auto_out_a_bits_data=_GEN ? io_dmi_req_bits_data:32'h0; 
  assign auto_out_d_ready=io_dmi_resp_ready; 
  assign io_dmi_req_ready=auto_out_a_ready; 
  assign io_dmi_resp_valid=auto_out_d_valid; 
  assign io_dmi_resp_bits_data=auto_out_d_bits_data; 
  assign io_dmi_resp_bits_resp={1'h0,auto_out_d_bits_corrupt|auto_out_d_bits_denied}; 
endmodule
 
module TLMonitor_29 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [6:0] io_in_a_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [6:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg inflight ;  
   reg [3:0] inflight_opcodes ;  
   reg [3:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire a_set=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg inflight_1 ;  
   reg [3:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire _GEN=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_0=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_1={io_in_a_bits_address[6:4]^3'h4,io_in_a_bits_address[2]}==4'h0|io_in_a_bits_address[6:3]==4'hA ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_3=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_4=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_6=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_7=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_8=io_in_a_valid&a_first_counter&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&~a_first_counter_1 ;  
   wire _GEN_9=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_10=_GEN_9&~d_release_ack ;  
   wire _GEN_11=_GEN_10&~_same_cycle_resp_T_1&~reset ;  
   wire _GEN_12=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
  always @( posedge clock)
       begin 
         if (_GEN)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&~_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&d_first_counter&~reset&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (a_set&~reset&inflight)
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~reset&~(inflight|_same_cycle_resp_T_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_same_cycle_resp_T_1&~reset&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&inflight_sizes[3:1]!=3'h2)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&~a_first_counter_1&io_in_a_valid&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~inflight_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&inflight_sizes_1[3:1]!=3'h2)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight_1|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:700:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire d_clr=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire [3:0] d_sizes_clr={4{d_clr}} ;  
   wire d_clr_1=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=1'h0;
              inflight_opcodes <=4'h0;
              inflight_sizes <=4'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=1'h0;
              inflight_sizes_1 <=4'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|a_set)&~d_clr;
              inflight_opcodes <=(inflight_opcodes|(a_set ? {io_in_a_bits_opcode,1'h1}:4'h0))&~d_sizes_clr;
              inflight_sizes <=(inflight_sizes|(a_set ? {1'h0,a_set ? 3'h5:3'h0}:4'h0))&~d_sizes_clr;
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~d_clr_1;
              inflight_sizes_1 <=inflight_sizes_1&~{4{d_clr_1}};
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            opcode_1 <=io_in_d_bits_opcode;
       end
  
endmodule
 
module TLDebugModuleOuter (
  input clock,
  input reset,
  output auto_dmi_in_a_ready,
  input auto_dmi_in_a_valid,
  input [2:0] auto_dmi_in_a_bits_opcode,
  input [6:0] auto_dmi_in_a_bits_address,
  input [31:0] auto_dmi_in_a_bits_data,
  input auto_dmi_in_d_ready,
  output auto_dmi_in_d_valid,
  output [2:0] auto_dmi_in_d_bits_opcode,
  output [31:0] auto_dmi_in_d_bits_data,
  output auto_int_out_0,
  output io_ctrl_ndreset,
  output io_ctrl_dmactive,
  input io_ctrl_dmactiveAck,
  input io_innerCtrl_ready,
  output io_innerCtrl_valid,
  output io_innerCtrl_bits_resumereq,
  output [9:0] io_innerCtrl_bits_hartsel,
  output io_innerCtrl_bits_ackhavereset,
  output io_innerCtrl_bits_hrmask_0,
  input io_hgDebugInt_0) ; 
   wire out_woready_9 ;  
   wire DMCONTROLWrData_setresethaltreq ;  
   wire DMCONTROLWrData_clrresethaltreq ;  
   reg DMCONTROLReg_haltreq ;  
   reg [9:0] DMCONTROLReg_hartsello ;  
   reg DMCONTROLReg_ndmreset ;  
   reg DMCONTROLReg_dmactive ;  
   reg hrmaskReg_0 ;  
   wire _GEN=DMCONTROLReg_hartsello==10'h0 ;  
   wire hrmaskNxt_0=~(~DMCONTROLReg_dmactive|out_woready_9&DMCONTROLWrData_clrresethaltreq&_GEN)&(out_woready_9&DMCONTROLWrData_setresethaltreq&_GEN|hrmaskReg_0) ;  
   wire in_bits_read=auto_dmi_in_a_bits_opcode==3'h4 ;  
   wire _out_T_3={auto_dmi_in_a_bits_address[4],auto_dmi_in_a_bits_address[2]}==2'h0 ;  
  assign DMCONTROLWrData_clrresethaltreq=auto_dmi_in_a_bits_data[2]; 
  assign DMCONTROLWrData_setresethaltreq=auto_dmi_in_a_bits_data[3]; 
  assign out_woready_9=auto_dmi_in_a_valid&auto_dmi_in_d_ready&~in_bits_read&~(auto_dmi_in_a_bits_address[3])&_out_T_3; 
   wire [2:0] dmiNodeIn_d_bits_opcode={2'h0,in_bits_read} ;  
   reg debugIntRegs_0 ;  
   reg innerCtrlValidReg ;  
   reg innerCtrlResumeReqReg ;  
   reg innerCtrlAckHaveResetReg ;  
   wire io_innerCtrl_valid_0=out_woready_9|innerCtrlValidReg ;  
   wire io_innerCtrl_bits_resumereq_0=out_woready_9&auto_dmi_in_a_bits_data[30]|innerCtrlResumeReqReg ;  
   wire io_innerCtrl_bits_ackhavereset_0=out_woready_9&auto_dmi_in_a_bits_data[28]|innerCtrlAckHaveResetReg ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              DMCONTROLReg_haltreq <=1'h0;
              DMCONTROLReg_hartsello <=10'h0;
              DMCONTROLReg_ndmreset <=1'h0;
              DMCONTROLReg_dmactive <=1'h0;
              hrmaskReg_0 <=1'h0;
              debugIntRegs_0 <=1'h0;
              innerCtrlValidReg <=1'h0;
              innerCtrlResumeReqReg <=1'h0;
              innerCtrlAckHaveResetReg <=1'h0;
            end 
          else 
            begin 
              DMCONTROLReg_haltreq <=DMCONTROLReg_dmactive&(out_woready_9 ? auto_dmi_in_a_bits_data[31]:DMCONTROLReg_haltreq);
              if (DMCONTROLReg_dmactive)
                 begin 
                 end 
               else 
                 DMCONTROLReg_hartsello <=10'h0;
              DMCONTROLReg_ndmreset <=DMCONTROLReg_dmactive&(out_woready_9 ? auto_dmi_in_a_bits_data[1]:DMCONTROLReg_ndmreset);
              if (out_woready_9)
                 DMCONTROLReg_dmactive <=auto_dmi_in_a_bits_data[0];
              hrmaskReg_0 <=hrmaskNxt_0;
              debugIntRegs_0 <=DMCONTROLReg_dmactive&(out_woready_9 ? auto_dmi_in_a_bits_data[31]:debugIntRegs_0);
              innerCtrlValidReg <=io_innerCtrl_valid_0&~io_innerCtrl_ready;
              innerCtrlResumeReqReg <=io_innerCtrl_bits_resumereq_0&~io_innerCtrl_ready;
              innerCtrlAckHaveResetReg <=io_innerCtrl_bits_ackhavereset_0&~io_innerCtrl_ready;
            end 
       end
  
  TLMonitor_29 monitor(.clock(clock),.reset(reset),.io_in_a_ready(auto_dmi_in_d_ready),.io_in_a_valid(auto_dmi_in_a_valid),.io_in_a_bits_opcode(auto_dmi_in_a_bits_opcode),.io_in_a_bits_address(auto_dmi_in_a_bits_address),.io_in_d_ready(auto_dmi_in_d_ready),.io_in_d_valid(auto_dmi_in_a_valid),.io_in_d_bits_opcode(dmiNodeIn_d_bits_opcode)); 
  assign auto_dmi_in_a_ready=auto_dmi_in_d_ready; 
  assign auto_dmi_in_d_valid=auto_dmi_in_a_valid; 
  assign auto_dmi_in_d_bits_opcode=dmiNodeIn_d_bits_opcode; 
  assign auto_dmi_in_d_bits_data=_out_T_3 ? (auto_dmi_in_a_bits_address[3] ? 32'h112380:{DMCONTROLReg_haltreq,29'h0,DMCONTROLReg_ndmreset,DMCONTROLReg_dmactive&io_ctrl_dmactiveAck}):32'h0; 
  assign auto_int_out_0=debugIntRegs_0|io_hgDebugInt_0; 
  assign io_ctrl_ndreset=DMCONTROLReg_ndmreset; 
  assign io_ctrl_dmactive=DMCONTROLReg_dmactive; 
  assign io_innerCtrl_valid=io_innerCtrl_valid_0; 
  assign io_innerCtrl_bits_resumereq=io_innerCtrl_bits_resumereq_0; 
  assign io_innerCtrl_bits_hartsel=DMCONTROLReg_hartsello; 
  assign io_innerCtrl_bits_ackhavereset=io_innerCtrl_bits_ackhavereset_0; 
  assign io_innerCtrl_bits_hrmask_0=hrmaskNxt_0; 
endmodule
 
module IntSyncCrossingSource_4 (
  input auto_in_0,
  output auto_out_sync_0) ; 
  assign auto_out_sync_0=auto_in_0; 
endmodule
 
module TLMonitor_30 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [8:0] io_in_a_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [1:0] io_in_d_bits_size,
  input io_in_d_bits_source,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [8:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [1:0] size_1 ;  
   reg source_1 ;  
   reg sink ;  
   reg denied ;  
   reg inflight ;  
   reg [3:0] inflight_opcodes ;  
   reg [3:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire [3:0] _GEN={1'h0,io_in_d_bits_source,2'h0} ;  
   wire [3:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire a_set=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg inflight_1 ;  
   reg [3:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire _GEN_0=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_1=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire [4:0] _GEN_2=io_in_a_bits_address[6:2]^5'h11 ;  
   wire _GEN_3=io_in_a_bits_address[8:6]==3'h0|{io_in_a_bits_address[8:7],_GEN_2[4:2],_GEN_2[0]}==6'h0|{io_in_a_bits_address[8:7],io_in_a_bits_address[6:3]^4'hB}==6'h0|{io_in_a_bits_address[8:7],~(io_in_a_bits_address[6:5])}==4'h0|{io_in_a_bits_address[8],~(io_in_a_bits_address[7])}==2'h0|io_in_a_bits_address[8] ;  
   wire _GEN_4=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_6=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_7=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_9=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_10=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_11=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_12=io_in_d_bits_param==2'h2 ;  
   wire _GEN_13=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_14=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_15=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_16=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_18=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_19=io_in_d_valid&d_first_counter&~reset ;  
   wire _GEN_20=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_21=_GEN_20&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&~a_first_counter_1&~io_in_d_bits_source ;  
   wire _GEN_22=_GEN_21&same_cycle_resp&~reset ;  
   wire _GEN_23=_GEN_21&~same_cycle_resp&~reset ;  
   wire [3:0] _GEN_24={2'h0,io_in_d_bits_size} ;  
   wire _GEN_25=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
   wire [3:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
   wire [3:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&~_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (a_set&~reset&inflight)
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~reset&~(inflight>>io_in_d_bits_source|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_d_bits_size!=2'h2)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_24!={1'h0,_a_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~a_first_counter_1&io_in_a_valid&~io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~(inflight_1>>io_in_d_bits_source))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_24!={1'h0,_c_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight_1|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/BusBypass.scala:32:12)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [30:0] _GEN_26={28'h0,io_in_d_bits_source,2'h0} ;  
   wire [30:0] _d_opcodes_clr_T_5=31'hF<<_GEN_26 ;  
   wire [30:0] _d_sizes_clr_T_5=31'hF<<_GEN_26 ;  
   wire [30:0] _d_sizes_clr_T_11=31'hF<<_GEN_26 ;  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_27=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire _GEN_28=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=1'h0;
              inflight_opcodes <=4'h0;
              inflight_sizes <=4'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=1'h0;
              inflight_sizes_1 <=4'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|a_set)&~(_GEN_27&~io_in_d_bits_source);
              inflight_opcodes <=(inflight_opcodes|(a_set ? {io_in_a_bits_opcode,1'h1}:4'h0))&~(_GEN_27 ? _d_opcodes_clr_T_5[3:0]:4'h0);
              inflight_sizes <=(inflight_sizes|(a_set ? {1'h0,a_set ? 3'h5:3'h0}:4'h0))&~(_GEN_27 ? _d_sizes_clr_T_5[3:0]:4'h0);
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_28&~io_in_d_bits_source);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_28 ? _d_sizes_clr_T_11[3:0]:4'h0);
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLBusBypassBar (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [8:0] auto_in_a_bits_address,
  input [31:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [1:0] auto_in_d_bits_size,
  output auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [31:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  input auto_out_1_a_ready,
  output auto_out_1_a_valid,
  output [2:0] auto_out_1_a_bits_opcode,
  output [8:0] auto_out_1_a_bits_address,
  output [31:0] auto_out_1_a_bits_data,
  output auto_out_1_d_ready,
  input auto_out_1_d_valid,
  input [2:0] auto_out_1_d_bits_opcode,
  input [1:0] auto_out_1_d_bits_param,
  input [1:0] auto_out_1_d_bits_size,
  input auto_out_1_d_bits_source,
  input auto_out_1_d_bits_sink,
  input auto_out_1_d_bits_denied,
  input [31:0] auto_out_1_d_bits_data,
  input auto_out_1_d_bits_corrupt,
  input auto_out_0_a_ready,
  output auto_out_0_a_valid,
  output [2:0] auto_out_0_a_bits_opcode,
  output [127:0] auto_out_0_a_bits_address,
  output auto_out_0_d_ready,
  input auto_out_0_d_valid,
  input [2:0] auto_out_0_d_bits_opcode,
  input [1:0] auto_out_0_d_bits_size,
  input auto_out_0_d_bits_denied,
  input auto_out_0_d_bits_corrupt,
  input io_bypass) ; 
   reg in_reset ;  
   reg bypass_reg ;  
   wire bypass=in_reset ? io_bypass:bypass_reg ;  
   reg [1:0] flight ;  
   reg counter ;  
   reg counter_3 ;  
   reg stall_counter ;  
   wire stall=bypass!=io_bypass&~stall_counter ;  
   wire nodeIn_a_ready=~stall&(bypass ? auto_out_0_a_ready:auto_out_1_a_ready) ;  
   wire nodeIn_d_valid=bypass ? auto_out_0_d_valid:auto_out_1_d_valid ;  
   wire [2:0] nodeIn_d_bits_opcode=bypass ? auto_out_0_d_bits_opcode:auto_out_1_d_bits_opcode ;  
   wire [1:0] nodeIn_d_bits_param=bypass ? 2'h0:auto_out_1_d_bits_param ;  
   wire [1:0] nodeIn_d_bits_size=bypass ? auto_out_0_d_bits_size:auto_out_1_d_bits_size ;  
   wire nodeIn_d_bits_sink=~bypass&auto_out_1_d_bits_sink ;  
   wire nodeIn_d_bits_denied=bypass ? auto_out_0_d_bits_denied:auto_out_1_d_bits_denied ;  
   wire nodeIn_d_bits_corrupt=bypass ? auto_out_0_d_bits_corrupt:auto_out_1_d_bits_corrupt ;  
   wire done=nodeIn_a_ready&auto_in_a_valid ;  
   wire d_dec=auto_in_d_ready&nodeIn_d_valid ;  
   wire [1:0] _next_flight_T_10=flight+{1'h0,d_dec&~counter_3&nodeIn_d_bits_opcode[2]&~(nodeIn_d_bits_opcode[1])}+{1'h0,done&~counter}-{1'h0,d_dec} ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              in_reset <=1'h1;
              flight <=2'h0;
              counter <=1'h0;
              counter_3 <=1'h0;
              stall_counter <=1'h0;
            end 
          else 
            begin 
              in_reset <=1'h0;
              flight <=_next_flight_T_10;
              counter <=(~done|counter-1'h1)&counter;
              counter_3 <=(~d_dec|counter_3-1'h1)&counter_3;
              stall_counter <=(~done|stall_counter-1'h1)&stall_counter;
            end 
         if (in_reset|_next_flight_T_10==2'h0)
            bypass_reg <=io_bypass;
       end
  
  TLMonitor_30 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(nodeIn_d_bits_opcode),.io_in_d_bits_param(nodeIn_d_bits_param),.io_in_d_bits_size(nodeIn_d_bits_size),.io_in_d_bits_source(~bypass&auto_out_1_d_bits_source),.io_in_d_bits_sink(nodeIn_d_bits_sink),.io_in_d_bits_denied(nodeIn_d_bits_denied),.io_in_d_bits_corrupt(nodeIn_d_bits_corrupt)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=nodeIn_d_bits_opcode; 
  assign auto_in_d_bits_param=nodeIn_d_bits_param; 
  assign auto_in_d_bits_size=nodeIn_d_bits_size; 
  assign auto_in_d_bits_sink=nodeIn_d_bits_sink; 
  assign auto_in_d_bits_denied=nodeIn_d_bits_denied; 
  assign auto_in_d_bits_data=bypass ? 32'h0:auto_out_1_d_bits_data; 
  assign auto_in_d_bits_corrupt=nodeIn_d_bits_corrupt; 
  assign auto_out_1_a_valid=~stall&auto_in_a_valid&~bypass; 
  assign auto_out_1_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_1_a_bits_address=auto_in_a_bits_address; 
  assign auto_out_1_a_bits_data=auto_in_a_bits_data; 
  assign auto_out_1_d_ready=auto_in_d_ready&~bypass; 
  assign auto_out_0_a_valid=~stall&auto_in_a_valid&bypass; 
  assign auto_out_0_a_bits_opcode=auto_in_a_bits_opcode; 
  assign auto_out_0_a_bits_address={119'h0,auto_in_a_bits_address}; 
  assign auto_out_0_d_ready=auto_in_d_ready&bypass; 
endmodule
 
module TLMonitor_31 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [127:0] io_in_a_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_size,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [127:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] size_1 ;  
   reg denied ;  
   reg inflight ;  
   reg [3:0] inflight_opcodes ;  
   reg [3:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire a_set=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (inflight_opcodes[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg inflight_1 ;  
   reg [3:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire _GEN=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_0=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_1=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_3=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_4=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_5=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_6=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_7=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_8=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_9=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_10=io_in_d_valid&d_first_counter&~reset ;  
   wire _same_cycle_resp_T_1=io_in_a_valid&~a_first_counter_1 ;  
   wire _GEN_11=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_12=_GEN_11&~d_release_ack ;  
   wire _GEN_13=_GEN_12&_same_cycle_resp_T_1&~reset ;  
   wire _GEN_14=_GEN_12&~_same_cycle_resp_T_1&~reset ;  
   wire [3:0] _GEN_15={2'h0,io_in_d_bits_size} ;  
   wire _GEN_16=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
  always @( posedge clock)
       begin 
         if (_GEN)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_3&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&~_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (a_set&~reset&inflight)
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&~reset&~(inflight|_same_cycle_resp_T_1))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_d_bits_size!=2'h2)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_15!={1'h0,inflight_sizes[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~a_first_counter_1&io_in_a_valid&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~inflight_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&_GEN_15!={1'h0,inflight_sizes_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight_1|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/BusBypass.scala:33:14)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire d_clr=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire [3:0] d_sizes_clr={4{d_clr}} ;  
   wire d_clr_1=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=1'h0;
              inflight_opcodes <=4'h0;
              inflight_sizes <=4'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=1'h0;
              inflight_sizes_1 <=4'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|a_set)&~d_clr;
              inflight_opcodes <=(inflight_opcodes|(a_set ? {io_in_a_bits_opcode,1'h1}:4'h0))&~d_sizes_clr;
              inflight_sizes <=(inflight_sizes|(a_set ? {1'h0,a_set ? 3'h5:3'h0}:4'h0))&~d_sizes_clr;
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~d_clr_1;
              inflight_sizes_1 <=inflight_sizes_1&~{4{d_clr_1}};
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module TLError_1 (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [127:0] auto_in_a_bits_address,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_size,
  output auto_in_d_bits_denied,
  output auto_in_d_bits_corrupt) ; 
   wire da_ready ;  
   reg [2:0] casez_tmp ;  
   reg idle ;  
   reg counter ;  
   wire nodeIn_a_ready=da_ready&idle ;  
   wire winner_1=auto_in_a_valid&idle ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg beatsLeft ;  
  always @( posedge clock)
       begin 
         if (~reset&~(idle|~counter))
            begin 
              if (1)$display("Assertion failed\n    at Error.scala:31 assert (idle || da_first) // we only send Grant, never GrantData => simplified flow control below\n");
              if (1)$display("");
            end 
       end
  
   reg state_1 ;  
   wire muxState_1=beatsLeft ? state_1:winner_1 ;  
  assign da_ready=auto_in_d_ready&(~beatsLeft|state_1); 
   wire nodeIn_d_valid=(~beatsLeft|state_1)&winner_1 ;  
   wire _nodeIn_d_bits_T_2=muxState_1&casez_tmp[0] ;  
   wire [1:0] _nodeIn_d_bits_T_17={muxState_1,1'h0} ;  
   wire [2:0] _nodeIn_d_bits_T_22=muxState_1 ? casez_tmp:3'h0 ;  
   wire done=da_ready&winner_1 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              idle <=1'h1;
              counter <=1'h0;
              beatsLeft <=1'h0;
              state_1 <=1'h0;
            end 
          else 
            begin 
              idle <=~(done&casez_tmp==3'h4)&idle;
              counter <=(~done|counter-1'h1)&counter;
              beatsLeft <=~(~beatsLeft&auto_in_d_ready)&beatsLeft-(auto_in_d_ready&nodeIn_d_valid);
              if (beatsLeft)
                 begin 
                 end 
               else 
                 state_1 <=winner_1;
            end 
       end
  
  TLMonitor_31 monitor(.clock(clock),.reset(reset),.io_in_a_ready(nodeIn_a_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(nodeIn_d_valid),.io_in_d_bits_opcode(_nodeIn_d_bits_T_22),.io_in_d_bits_size(_nodeIn_d_bits_T_17),.io_in_d_bits_denied(muxState_1),.io_in_d_bits_corrupt(_nodeIn_d_bits_T_2)); 
  assign auto_in_a_ready=nodeIn_a_ready; 
  assign auto_in_d_valid=nodeIn_d_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_bits_T_22; 
  assign auto_in_d_bits_size=_nodeIn_d_bits_T_17; 
  assign auto_in_d_bits_denied=muxState_1; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_bits_T_2; 
endmodule
 
module TLBusBypass (
  input clock,
  input reset,
  input auto_node_out_out_a_ready,
  output auto_node_out_out_a_valid,
  output [2:0] auto_node_out_out_a_bits_opcode,
  output [8:0] auto_node_out_out_a_bits_address,
  output [31:0] auto_node_out_out_a_bits_data,
  output auto_node_out_out_d_ready,
  input auto_node_out_out_d_valid,
  input [2:0] auto_node_out_out_d_bits_opcode,
  input [1:0] auto_node_out_out_d_bits_param,
  input [1:0] auto_node_out_out_d_bits_size,
  input auto_node_out_out_d_bits_source,
  input auto_node_out_out_d_bits_sink,
  input auto_node_out_out_d_bits_denied,
  input [31:0] auto_node_out_out_d_bits_data,
  input auto_node_out_out_d_bits_corrupt,
  output auto_node_in_in_a_ready,
  input auto_node_in_in_a_valid,
  input [2:0] auto_node_in_in_a_bits_opcode,
  input [8:0] auto_node_in_in_a_bits_address,
  input [31:0] auto_node_in_in_a_bits_data,
  input auto_node_in_in_d_ready,
  output auto_node_in_in_d_valid,
  output [2:0] auto_node_in_in_d_bits_opcode,
  output [1:0] auto_node_in_in_d_bits_param,
  output [1:0] auto_node_in_in_d_bits_size,
  output auto_node_in_in_d_bits_sink,
  output auto_node_in_in_d_bits_denied,
  output [31:0] auto_node_in_in_d_bits_data,
  output auto_node_in_in_d_bits_corrupt,
  input io_bypass) ; 
   wire _error_auto_in_a_ready ;  
   wire _error_auto_in_d_valid ;  
   wire [2:0] _error_auto_in_d_bits_opcode ;  
   wire [1:0] _error_auto_in_d_bits_size ;  
   wire _error_auto_in_d_bits_denied ;  
   wire _error_auto_in_d_bits_corrupt ;  
   wire _bar_auto_out_0_a_valid ;  
   wire [2:0] _bar_auto_out_0_a_bits_opcode ;  
   wire [127:0] _bar_auto_out_0_a_bits_address ;  
   wire _bar_auto_out_0_d_ready ;  
  TLBusBypassBar bar(.clock(clock),.reset(reset),.auto_in_a_ready(auto_node_in_in_a_ready),.auto_in_a_valid(auto_node_in_in_a_valid),.auto_in_a_bits_opcode(auto_node_in_in_a_bits_opcode),.auto_in_a_bits_address(auto_node_in_in_a_bits_address),.auto_in_a_bits_data(auto_node_in_in_a_bits_data),.auto_in_d_ready(auto_node_in_in_d_ready),.auto_in_d_valid(auto_node_in_in_d_valid),.auto_in_d_bits_opcode(auto_node_in_in_d_bits_opcode),.auto_in_d_bits_param(auto_node_in_in_d_bits_param),.auto_in_d_bits_size(auto_node_in_in_d_bits_size),.auto_in_d_bits_sink(auto_node_in_in_d_bits_sink),.auto_in_d_bits_denied(auto_node_in_in_d_bits_denied),.auto_in_d_bits_data(auto_node_in_in_d_bits_data),.auto_in_d_bits_corrupt(auto_node_in_in_d_bits_corrupt),.auto_out_1_a_ready(auto_node_out_out_a_ready),.auto_out_1_a_valid(auto_node_out_out_a_valid),.auto_out_1_a_bits_opcode(auto_node_out_out_a_bits_opcode),.auto_out_1_a_bits_address(auto_node_out_out_a_bits_address),.auto_out_1_a_bits_data(auto_node_out_out_a_bits_data),.auto_out_1_d_ready(auto_node_out_out_d_ready),.auto_out_1_d_valid(auto_node_out_out_d_valid),.auto_out_1_d_bits_opcode(auto_node_out_out_d_bits_opcode),.auto_out_1_d_bits_param(auto_node_out_out_d_bits_param),.auto_out_1_d_bits_size(auto_node_out_out_d_bits_size),.auto_out_1_d_bits_source(auto_node_out_out_d_bits_source),.auto_out_1_d_bits_sink(auto_node_out_out_d_bits_sink),.auto_out_1_d_bits_denied(auto_node_out_out_d_bits_denied),.auto_out_1_d_bits_data(auto_node_out_out_d_bits_data),.auto_out_1_d_bits_corrupt(auto_node_out_out_d_bits_corrupt),.auto_out_0_a_ready(_error_auto_in_a_ready),.auto_out_0_a_valid(_bar_auto_out_0_a_valid),.auto_out_0_a_bits_opcode(_bar_auto_out_0_a_bits_opcode),.auto_out_0_a_bits_address(_bar_auto_out_0_a_bits_address),.auto_out_0_d_ready(_bar_auto_out_0_d_ready),.auto_out_0_d_valid(_error_auto_in_d_valid),.auto_out_0_d_bits_opcode(_error_auto_in_d_bits_opcode),.auto_out_0_d_bits_size(_error_auto_in_d_bits_size),.auto_out_0_d_bits_denied(_error_auto_in_d_bits_denied),.auto_out_0_d_bits_corrupt(_error_auto_in_d_bits_corrupt),.io_bypass(io_bypass)); 
  TLError_1 error(.clock(clock),.reset(reset),.auto_in_a_ready(_error_auto_in_a_ready),.auto_in_a_valid(_bar_auto_out_0_a_valid),.auto_in_a_bits_opcode(_bar_auto_out_0_a_bits_opcode),.auto_in_a_bits_address(_bar_auto_out_0_a_bits_address),.auto_in_d_ready(_bar_auto_out_0_d_ready),.auto_in_d_valid(_error_auto_in_d_valid),.auto_in_d_bits_opcode(_error_auto_in_d_bits_opcode),.auto_in_d_bits_size(_error_auto_in_d_bits_size),.auto_in_d_bits_denied(_error_auto_in_d_bits_denied),.auto_in_d_bits_corrupt(_error_auto_in_d_bits_corrupt)); 
endmodule
 
module TLMonitor_32 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [8:0] io_in_a_bits_address,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_param,
  input [1:0] io_in_d_bits_size,
  input io_in_d_bits_source,
  input io_in_d_bits_sink,
  input io_in_d_bits_denied,
  input io_in_d_bits_corrupt) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [8:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] param_1 ;  
   reg [1:0] size_1 ;  
   reg source_1 ;  
   reg sink ;  
   reg denied ;  
   reg inflight ;  
   reg [3:0] inflight_opcodes ;  
   reg [3:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire [3:0] _GEN={1'h0,io_in_d_bits_source,2'h0} ;  
   wire [3:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire a_set=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg inflight_1 ;  
   reg [3:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire _GEN_0=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_1=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire [4:0] _GEN_2=io_in_a_bits_address[6:2]^5'h11 ;  
   wire _GEN_3=io_in_a_bits_address[8:6]==3'h0|{io_in_a_bits_address[8:7],_GEN_2[4:2],_GEN_2[0]}==6'h0|{io_in_a_bits_address[8:7],io_in_a_bits_address[6:3]^4'hB}==6'h0|{io_in_a_bits_address[8:7],~(io_in_a_bits_address[6:5])}==4'h0|{io_in_a_bits_address[8],~(io_in_a_bits_address[7])}==2'h0|io_in_a_bits_address[8] ;  
   wire _GEN_4=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_5=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_6=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_7=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_8=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_9=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_10=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_11=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_12=io_in_d_bits_param==2'h2 ;  
   wire _GEN_13=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_14=~io_in_d_bits_denied|io_in_d_bits_corrupt ;  
   wire _GEN_15=io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset ;  
   wire _GEN_16=io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset ;  
   wire _GEN_18=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_19=io_in_d_valid&d_first_counter&~reset ;  
   wire a_set_wo_ready=io_in_a_valid&~a_first_counter_1 ;  
   wire _GEN_20=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_21=_GEN_20&~d_release_ack ;  
   wire same_cycle_resp=a_set_wo_ready&~io_in_d_bits_source ;  
   wire _GEN_22=_GEN_21&same_cycle_resp&~reset ;  
   wire _GEN_23=_GEN_21&~same_cycle_resp&~reset ;  
   wire [3:0] _GEN_24={2'h0,io_in_d_bits_size} ;  
   wire _GEN_25=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
   wire [3:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
   wire [3:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_0)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_1)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&~_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_4&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|(io_in_a_bits_address[1:0])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant is denied (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(&io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData is denied (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck is denied (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData is denied (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&(|io_in_d_bits_param))
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck is denied (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_param!=param_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_sink!=sink)
            begin 
              if (1)$display("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_d_bits_denied!=denied)
            begin 
              if (1)$display("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (a_set&~reset&inflight)
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~reset&~(inflight>>io_in_d_bits_source|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&io_in_d_bits_size!=2'h2)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&_GEN_24!={1'h0,_a_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&~a_first_counter_1&io_in_a_valid&~io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(a_set_wo_ready!=(_GEN_21&~io_in_d_bits_source)|~a_set_wo_ready))
            begin 
              if (1)$display("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~(inflight_1>>io_in_d_bits_source))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_24!={1'h0,_c_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight_1|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:699:46)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [30:0] _GEN_26={28'h0,io_in_d_bits_source,2'h0} ;  
   wire [30:0] _d_opcodes_clr_T_5=31'hF<<_GEN_26 ;  
   wire [30:0] _d_sizes_clr_T_5=31'hF<<_GEN_26 ;  
   wire [30:0] _d_sizes_clr_T_11=31'hF<<_GEN_26 ;  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_27=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire _GEN_28=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=1'h0;
              inflight_opcodes <=4'h0;
              inflight_sizes <=4'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=1'h0;
              inflight_sizes_1 <=4'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|a_set)&~(_GEN_27&~io_in_d_bits_source);
              inflight_opcodes <=(inflight_opcodes|(a_set ? {io_in_a_bits_opcode,1'h1}:4'h0))&~(_GEN_27 ? _d_opcodes_clr_T_5[3:0]:4'h0);
              inflight_sizes <=(inflight_sizes|(a_set ? {1'h0,a_set ? 3'h5:3'h0}:4'h0))&~(_GEN_27 ? _d_sizes_clr_T_5[3:0]:4'h0);
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_28&~io_in_d_bits_source);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_28 ? _d_sizes_clr_T_11[3:0]:4'h0);
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              param_1 <=io_in_d_bits_param;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
              sink <=io_in_d_bits_sink;
              denied <=io_in_d_bits_denied;
            end 
       end
  
endmodule
 
module AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 (
  input clock,
  input reset,
  input io_d,
  output io_q) ; 
   reg sync_0 ;  
   reg sync_1 ;  
   reg sync_2 ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              sync_0 <=1'h0;
              sync_1 <=1'h0;
              sync_2 <=1'h0;
            end 
          else 
            begin 
              sync_0 <=sync_1;
              sync_1 <=sync_2;
              sync_2 <=io_d;
            end 
       end
  
  assign io_q=sync_0; 
endmodule
 
module AsyncResetSynchronizerShiftReg_w1_d3_i0 (
  input clock,
  input reset,
  input io_d,
  output io_q) ; 
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain(.clock(clock),.reset(reset),.io_d(io_d),.io_q(io_q)); 
endmodule
 
module AsyncResetSynchronizerShiftReg_w1_d3_i0_1 (
  input clock,
  input reset,
  input io_d,
  output io_q) ; 
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain(.clock(clock),.reset(reset),.io_d(io_d),.io_q(io_q)); 
endmodule
 
module AsyncValidSync (
  input io_in,
  output io_out,
  input clock,
  input reset) ; 
  AsyncResetSynchronizerShiftReg_w1_d3_i0_1 io_out_source_valid_0(.clock(clock),.reset(reset),.io_d(io_in),.io_q(io_out)); 
endmodule
 
module AsyncQueueSource (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [8:0] io_enq_bits_address,
  input [31:0] io_enq_bits_data,
  output [2:0] io_async_mem_0_opcode,
  output [8:0] io_async_mem_0_address,
  output [31:0] io_async_mem_0_data,
  input io_async_ridx,
  output io_async_widx,
  input io_async_safe_ridx_valid,
  output io_async_safe_widx_valid,
  output io_async_safe_source_reset_n,
  input io_async_safe_sink_reset_n) ; 
   wire io_enq_ready_0 ;  
   wire _sink_valid_io_out ;  
   wire _sink_extend_io_out ;  
   wire _source_valid_0_io_out ;  
   wire _ridx_ridx_gray_io_q ;  
   reg [2:0] mem_0_opcode ;  
   reg [8:0] mem_0_address ;  
   reg [31:0] mem_0_data ;  
   wire _widx_T_1=io_enq_ready_0&io_enq_valid ;  
   reg widx_widx_bin ;  
   reg ready_reg ;  
  assign io_enq_ready_0=ready_reg&_sink_valid_io_out; 
   reg widx_gray ;  
  always @( posedge clock)
       begin 
         if (_widx_T_1)
            begin 
              mem_0_opcode <=io_enq_bits_opcode;
              mem_0_address <=io_enq_bits_address;
              mem_0_data <=io_enq_bits_data;
            end 
       end
  
   wire widx=_sink_valid_io_out&widx_widx_bin+_widx_T_1 ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              widx_widx_bin <=1'h0;
              ready_reg <=1'h0;
              widx_gray <=1'h0;
            end 
          else 
            begin 
              widx_widx_bin <=widx;
              ready_reg <=_sink_valid_io_out&widx!=~_ridx_ridx_gray_io_q;
              widx_gray <=widx;
            end 
       end
  
  AsyncResetSynchronizerShiftReg_w1_d3_i0 ridx_ridx_gray(.clock(clock),.reset(reset),.io_d(io_async_ridx),.io_q(_ridx_ridx_gray_io_q)); 
  AsyncValidSync source_valid_0(.io_in(1'h1),.io_out(_source_valid_0_io_out),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync source_valid_1(.io_in(_source_valid_0_io_out),.io_out(io_async_safe_widx_valid),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync sink_extend(.io_in(io_async_safe_ridx_valid),.io_out(_sink_extend_io_out),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync sink_valid(.io_in(_sink_extend_io_out),.io_out(_sink_valid_io_out),.clock(clock),.reset(reset)); 
  assign io_enq_ready=io_enq_ready_0; 
  assign io_async_mem_0_opcode=mem_0_opcode; 
  assign io_async_mem_0_address=mem_0_address; 
  assign io_async_mem_0_data=mem_0_data; 
  assign io_async_widx=widx_gray; 
  assign io_async_safe_source_reset_n=~reset; 
endmodule
 
module ClockCrossingReg_w43 (
  input clock,
  input [42:0] io_d,
  output [42:0] io_q,
  input io_en) ; 
   reg [42:0] cdc_reg ;  
  always @( posedge clock)
       begin 
         if (io_en)
            cdc_reg <=io_d;
       end
  
  assign io_q=cdc_reg; 
endmodule
 
module AsyncQueueSink (
  input clock,
  input reset,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [1:0] io_deq_bits_param,
  output [1:0] io_deq_bits_size,
  output io_deq_bits_source,
  output io_deq_bits_sink,
  output io_deq_bits_denied,
  output [31:0] io_deq_bits_data,
  output io_deq_bits_corrupt,
  input [2:0] io_async_mem_0_opcode,
  input [1:0] io_async_mem_0_size,
  input io_async_mem_0_source,
  input [31:0] io_async_mem_0_data,
  output io_async_ridx,
  input io_async_widx,
  output io_async_safe_ridx_valid,
  input io_async_safe_widx_valid,
  input io_async_safe_source_reset_n,
  output io_async_safe_sink_reset_n) ; 
   wire io_deq_valid_0 ;  
   wire _source_valid_io_out ;  
   wire _source_extend_io_out ;  
   wire _sink_valid_0_io_out ;  
   wire [42:0] _io_deq_bits_deq_bits_reg_io_q ;  
   wire _widx_widx_gray_io_q ;  
   reg ridx_ridx_bin ;  
   wire ridx=_source_valid_io_out&ridx_ridx_bin+(io_deq_ready&io_deq_valid_0) ;  
   wire valid=_source_valid_io_out&ridx!=_widx_widx_gray_io_q ;  
   reg valid_reg ;  
  assign io_deq_valid_0=valid_reg&_source_valid_io_out; 
   reg ridx_gray ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              ridx_ridx_bin <=1'h0;
              valid_reg <=1'h0;
              ridx_gray <=1'h0;
            end 
          else 
            begin 
              ridx_ridx_bin <=ridx;
              valid_reg <=valid;
              ridx_gray <=ridx;
            end 
       end
  
  AsyncResetSynchronizerShiftReg_w1_d3_i0 widx_widx_gray(.clock(clock),.reset(reset),.io_d(io_async_widx),.io_q(_widx_widx_gray_io_q)); 
  ClockCrossingReg_w43 io_deq_bits_deq_bits_reg(.clock(clock),.io_d({io_async_mem_0_opcode,2'h0,io_async_mem_0_size,io_async_mem_0_source,2'h0,io_async_mem_0_data,1'h0}),.io_q(_io_deq_bits_deq_bits_reg_io_q),.io_en(valid)); 
  AsyncValidSync sink_valid_0(.io_in(1'h1),.io_out(_sink_valid_0_io_out),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync sink_valid_1(.io_in(_sink_valid_0_io_out),.io_out(io_async_safe_ridx_valid),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync source_extend(.io_in(io_async_safe_widx_valid),.io_out(_source_extend_io_out),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync source_valid(.io_in(_source_extend_io_out),.io_out(_source_valid_io_out),.clock(clock),.reset(reset)); 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_opcode=_io_deq_bits_deq_bits_reg_io_q[42:40]; 
  assign io_deq_bits_param=_io_deq_bits_deq_bits_reg_io_q[39:38]; 
  assign io_deq_bits_size=_io_deq_bits_deq_bits_reg_io_q[37:36]; 
  assign io_deq_bits_source=_io_deq_bits_deq_bits_reg_io_q[35]; 
  assign io_deq_bits_sink=_io_deq_bits_deq_bits_reg_io_q[34]; 
  assign io_deq_bits_denied=_io_deq_bits_deq_bits_reg_io_q[33]; 
  assign io_deq_bits_data=_io_deq_bits_deq_bits_reg_io_q[32:1]; 
  assign io_deq_bits_corrupt=_io_deq_bits_deq_bits_reg_io_q[0]; 
  assign io_async_ridx=ridx_gray; 
  assign io_async_safe_sink_reset_n=~reset; 
endmodule
 
module TLAsyncCrossingSource (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [8:0] auto_in_a_bits_address,
  input [31:0] auto_in_a_bits_data,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [2:0] auto_in_d_bits_opcode,
  output [1:0] auto_in_d_bits_param,
  output [1:0] auto_in_d_bits_size,
  output auto_in_d_bits_source,
  output auto_in_d_bits_sink,
  output auto_in_d_bits_denied,
  output [31:0] auto_in_d_bits_data,
  output auto_in_d_bits_corrupt,
  output [2:0] auto_out_a_mem_0_opcode,
  output [8:0] auto_out_a_mem_0_address,
  output [31:0] auto_out_a_mem_0_data,
  input auto_out_a_ridx,
  output auto_out_a_widx,
  input auto_out_a_safe_ridx_valid,
  output auto_out_a_safe_widx_valid,
  output auto_out_a_safe_source_reset_n,
  input auto_out_a_safe_sink_reset_n,
  input [2:0] auto_out_d_mem_0_opcode,
  input [1:0] auto_out_d_mem_0_size,
  input auto_out_d_mem_0_source,
  input [31:0] auto_out_d_mem_0_data,
  output auto_out_d_ridx,
  input auto_out_d_widx,
  output auto_out_d_safe_ridx_valid,
  input auto_out_d_safe_widx_valid,
  input auto_out_d_safe_source_reset_n,
  output auto_out_d_safe_sink_reset_n) ; 
   wire _nodeIn_d_sink_io_deq_valid ;  
   wire [2:0] _nodeIn_d_sink_io_deq_bits_opcode ;  
   wire [1:0] _nodeIn_d_sink_io_deq_bits_param ;  
   wire [1:0] _nodeIn_d_sink_io_deq_bits_size ;  
   wire _nodeIn_d_sink_io_deq_bits_source ;  
   wire _nodeIn_d_sink_io_deq_bits_sink ;  
   wire _nodeIn_d_sink_io_deq_bits_denied ;  
   wire _nodeIn_d_sink_io_deq_bits_corrupt ;  
   wire _nodeOut_a_source_io_enq_ready ;  
  TLMonitor_32 monitor(.clock(clock),.reset(reset),.io_in_a_ready(_nodeOut_a_source_io_enq_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(_nodeIn_d_sink_io_deq_valid),.io_in_d_bits_opcode(_nodeIn_d_sink_io_deq_bits_opcode),.io_in_d_bits_param(_nodeIn_d_sink_io_deq_bits_param),.io_in_d_bits_size(_nodeIn_d_sink_io_deq_bits_size),.io_in_d_bits_source(_nodeIn_d_sink_io_deq_bits_source),.io_in_d_bits_sink(_nodeIn_d_sink_io_deq_bits_sink),.io_in_d_bits_denied(_nodeIn_d_sink_io_deq_bits_denied),.io_in_d_bits_corrupt(_nodeIn_d_sink_io_deq_bits_corrupt)); 
  AsyncQueueSource nodeOut_a_source(.clock(clock),.reset(reset),.io_enq_ready(_nodeOut_a_source_io_enq_ready),.io_enq_valid(auto_in_a_valid),.io_enq_bits_opcode(auto_in_a_bits_opcode),.io_enq_bits_address(auto_in_a_bits_address),.io_enq_bits_data(auto_in_a_bits_data),.io_async_mem_0_opcode(auto_out_a_mem_0_opcode),.io_async_mem_0_address(auto_out_a_mem_0_address),.io_async_mem_0_data(auto_out_a_mem_0_data),.io_async_ridx(auto_out_a_ridx),.io_async_widx(auto_out_a_widx),.io_async_safe_ridx_valid(auto_out_a_safe_ridx_valid),.io_async_safe_widx_valid(auto_out_a_safe_widx_valid),.io_async_safe_source_reset_n(auto_out_a_safe_source_reset_n),.io_async_safe_sink_reset_n(auto_out_a_safe_sink_reset_n)); 
  AsyncQueueSink nodeIn_d_sink(.clock(clock),.reset(reset),.io_deq_ready(auto_in_d_ready),.io_deq_valid(_nodeIn_d_sink_io_deq_valid),.io_deq_bits_opcode(_nodeIn_d_sink_io_deq_bits_opcode),.io_deq_bits_param(_nodeIn_d_sink_io_deq_bits_param),.io_deq_bits_size(_nodeIn_d_sink_io_deq_bits_size),.io_deq_bits_source(_nodeIn_d_sink_io_deq_bits_source),.io_deq_bits_sink(_nodeIn_d_sink_io_deq_bits_sink),.io_deq_bits_denied(_nodeIn_d_sink_io_deq_bits_denied),.io_deq_bits_data(auto_in_d_bits_data),.io_deq_bits_corrupt(_nodeIn_d_sink_io_deq_bits_corrupt),.io_async_mem_0_opcode(auto_out_d_mem_0_opcode),.io_async_mem_0_size(auto_out_d_mem_0_size),.io_async_mem_0_source(auto_out_d_mem_0_source),.io_async_mem_0_data(auto_out_d_mem_0_data),.io_async_ridx(auto_out_d_ridx),.io_async_widx(auto_out_d_widx),.io_async_safe_ridx_valid(auto_out_d_safe_ridx_valid),.io_async_safe_widx_valid(auto_out_d_safe_widx_valid),.io_async_safe_source_reset_n(auto_out_d_safe_source_reset_n),.io_async_safe_sink_reset_n(auto_out_d_safe_sink_reset_n)); 
  assign auto_in_a_ready=_nodeOut_a_source_io_enq_ready; 
  assign auto_in_d_valid=_nodeIn_d_sink_io_deq_valid; 
  assign auto_in_d_bits_opcode=_nodeIn_d_sink_io_deq_bits_opcode; 
  assign auto_in_d_bits_param=_nodeIn_d_sink_io_deq_bits_param; 
  assign auto_in_d_bits_size=_nodeIn_d_sink_io_deq_bits_size; 
  assign auto_in_d_bits_source=_nodeIn_d_sink_io_deq_bits_source; 
  assign auto_in_d_bits_sink=_nodeIn_d_sink_io_deq_bits_sink; 
  assign auto_in_d_bits_denied=_nodeIn_d_sink_io_deq_bits_denied; 
  assign auto_in_d_bits_corrupt=_nodeIn_d_sink_io_deq_bits_corrupt; 
endmodule
 
module AsyncQueueSource_1 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input io_enq_bits_resumereq,
  input [9:0] io_enq_bits_hartsel,
  input io_enq_bits_ackhavereset,
  input io_enq_bits_hrmask_0,
  output io_async_mem_resumereq_0,
  output [9:0] io_async_mem_hartsel_0,
  output io_async_mem_ackhavereset_0,
  output io_async_mem_hrmask_0_0,
  input io_async_ridx,
  output io_async_widx,
  input io_async_safe_ridx_valid,
  output io_async_safe_widx_valid,
  output io_async_safe_source_reset_n,
  input io_async_safe_sink_reset_n) ; 
   wire io_enq_ready_0 ;  
   wire _sink_valid_io_out ;  
   wire _sink_extend_io_out ;  
   wire _source_valid_0_io_out ;  
   wire _ridx_ridx_gray_io_q ;  
   reg mem_resumereq_0 ;  
   reg [9:0] mem_hartsel_0 ;  
   reg mem_ackhavereset_0 ;  
   reg mem_hrmask_0_0 ;  
   wire _widx_T_1=io_enq_ready_0&io_enq_valid ;  
   reg widx_widx_bin ;  
   reg ready_reg ;  
  assign io_enq_ready_0=ready_reg&_sink_valid_io_out; 
   reg widx_gray ;  
  always @( posedge clock)
       begin 
         if (_widx_T_1)
            begin 
              mem_resumereq_0 <=io_enq_bits_resumereq;
              mem_hartsel_0 <=io_enq_bits_hartsel;
              mem_ackhavereset_0 <=io_enq_bits_ackhavereset;
              mem_hrmask_0_0 <=io_enq_bits_hrmask_0;
            end 
       end
  
   wire widx=_sink_valid_io_out&widx_widx_bin+_widx_T_1 ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              widx_widx_bin <=1'h0;
              ready_reg <=1'h0;
              widx_gray <=1'h0;
            end 
          else 
            begin 
              widx_widx_bin <=widx;
              ready_reg <=_sink_valid_io_out&widx!=~_ridx_ridx_gray_io_q;
              widx_gray <=widx;
            end 
       end
  
  AsyncResetSynchronizerShiftReg_w1_d3_i0 ridx_ridx_gray(.clock(clock),.reset(reset),.io_d(io_async_ridx),.io_q(_ridx_ridx_gray_io_q)); 
  AsyncValidSync source_valid_0(.io_in(1'h1),.io_out(_source_valid_0_io_out),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync source_valid_1(.io_in(_source_valid_0_io_out),.io_out(io_async_safe_widx_valid),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync sink_extend(.io_in(io_async_safe_ridx_valid),.io_out(_sink_extend_io_out),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync sink_valid(.io_in(_sink_extend_io_out),.io_out(_sink_valid_io_out),.clock(clock),.reset(reset)); 
  assign io_enq_ready=io_enq_ready_0; 
  assign io_async_mem_resumereq_0=mem_resumereq_0; 
  assign io_async_mem_hartsel_0=mem_hartsel_0; 
  assign io_async_mem_ackhavereset_0=mem_ackhavereset_0; 
  assign io_async_mem_hrmask_0_0=mem_hrmask_0_0; 
  assign io_async_widx=widx_gray; 
  assign io_async_safe_source_reset_n=~reset; 
endmodule
 
module TLDebugModuleOuterAsync (
  output [2:0] auto_asource_out_a_mem_0_opcode,
  output [8:0] auto_asource_out_a_mem_0_address,
  output [31:0] auto_asource_out_a_mem_0_data,
  input auto_asource_out_a_ridx,
  output auto_asource_out_a_widx,
  input auto_asource_out_a_safe_ridx_valid,
  output auto_asource_out_a_safe_widx_valid,
  output auto_asource_out_a_safe_source_reset_n,
  input auto_asource_out_a_safe_sink_reset_n,
  input [2:0] auto_asource_out_d_mem_0_opcode,
  input [1:0] auto_asource_out_d_mem_0_size,
  input auto_asource_out_d_mem_0_source,
  input [31:0] auto_asource_out_d_mem_0_data,
  output auto_asource_out_d_ridx,
  input auto_asource_out_d_widx,
  output auto_asource_out_d_safe_ridx_valid,
  input auto_asource_out_d_safe_widx_valid,
  input auto_asource_out_d_safe_source_reset_n,
  output auto_asource_out_d_safe_sink_reset_n,
  output auto_intsource_out_sync_0,
  input io_dmi_clock,
  input io_dmi_reset,
  output io_dmi_req_ready,
  input io_dmi_req_valid,
  input [6:0] io_dmi_req_bits_addr,
  input [31:0] io_dmi_req_bits_data,
  input [1:0] io_dmi_req_bits_op,
  input io_dmi_resp_ready,
  output io_dmi_resp_valid,
  output [31:0] io_dmi_resp_bits_data,
  output [1:0] io_dmi_resp_bits_resp,
  output io_ctrl_ndreset,
  output io_ctrl_dmactive,
  input io_ctrl_dmactiveAck,
  output io_innerCtrl_mem_resumereq_0,
  output [9:0] io_innerCtrl_mem_hartsel_0,
  output io_innerCtrl_mem_ackhavereset_0,
  output io_innerCtrl_mem_hrmask_0_0,
  input io_innerCtrl_ridx,
  output io_innerCtrl_widx,
  input io_innerCtrl_safe_ridx_valid,
  output io_innerCtrl_safe_widx_valid,
  output io_innerCtrl_safe_source_reset_n,
  input io_innerCtrl_safe_sink_reset_n,
  input io_hgDebugInt_0) ; 
   wire _io_innerCtrl_source_io_enq_ready ;  
   wire _dmactiveAck_dmactiveAckSync_io_q ;  
   wire _asource_auto_in_a_ready ;  
   wire _asource_auto_in_d_valid ;  
   wire [2:0] _asource_auto_in_d_bits_opcode ;  
   wire [1:0] _asource_auto_in_d_bits_param ;  
   wire [1:0] _asource_auto_in_d_bits_size ;  
   wire _asource_auto_in_d_bits_source ;  
   wire _asource_auto_in_d_bits_sink ;  
   wire _asource_auto_in_d_bits_denied ;  
   wire [31:0] _asource_auto_in_d_bits_data ;  
   wire _asource_auto_in_d_bits_corrupt ;  
   wire _dmiBypass_auto_node_out_out_a_valid ;  
   wire [2:0] _dmiBypass_auto_node_out_out_a_bits_opcode ;  
   wire [8:0] _dmiBypass_auto_node_out_out_a_bits_address ;  
   wire [31:0] _dmiBypass_auto_node_out_out_a_bits_data ;  
   wire _dmiBypass_auto_node_out_out_d_ready ;  
   wire _dmiBypass_auto_node_in_in_a_ready ;  
   wire _dmiBypass_auto_node_in_in_d_valid ;  
   wire [2:0] _dmiBypass_auto_node_in_in_d_bits_opcode ;  
   wire [1:0] _dmiBypass_auto_node_in_in_d_bits_param ;  
   wire [1:0] _dmiBypass_auto_node_in_in_d_bits_size ;  
   wire _dmiBypass_auto_node_in_in_d_bits_sink ;  
   wire _dmiBypass_auto_node_in_in_d_bits_denied ;  
   wire [31:0] _dmiBypass_auto_node_in_in_d_bits_data ;  
   wire _dmiBypass_auto_node_in_in_d_bits_corrupt ;  
   wire _dmOuter_auto_dmi_in_a_ready ;  
   wire _dmOuter_auto_dmi_in_d_valid ;  
   wire [2:0] _dmOuter_auto_dmi_in_d_bits_opcode ;  
   wire [31:0] _dmOuter_auto_dmi_in_d_bits_data ;  
   wire _dmOuter_auto_int_out_0 ;  
   wire _dmOuter_io_ctrl_dmactive ;  
   wire _dmOuter_io_innerCtrl_valid ;  
   wire _dmOuter_io_innerCtrl_bits_resumereq ;  
   wire [9:0] _dmOuter_io_innerCtrl_bits_hartsel ;  
   wire _dmOuter_io_innerCtrl_bits_ackhavereset ;  
   wire _dmOuter_io_innerCtrl_bits_hrmask_0 ;  
   wire _dmi2tl_auto_out_a_valid ;  
   wire [2:0] _dmi2tl_auto_out_a_bits_opcode ;  
   wire [8:0] _dmi2tl_auto_out_a_bits_address ;  
   wire [31:0] _dmi2tl_auto_out_a_bits_data ;  
   wire _dmi2tl_auto_out_d_ready ;  
   wire _dmiXbar_auto_in_a_ready ;  
   wire _dmiXbar_auto_in_d_valid ;  
   wire _dmiXbar_auto_in_d_bits_denied ;  
   wire [31:0] _dmiXbar_auto_in_d_bits_data ;  
   wire _dmiXbar_auto_in_d_bits_corrupt ;  
   wire _dmiXbar_auto_out_1_a_valid ;  
   wire [2:0] _dmiXbar_auto_out_1_a_bits_opcode ;  
   wire [6:0] _dmiXbar_auto_out_1_a_bits_address ;  
   wire [31:0] _dmiXbar_auto_out_1_a_bits_data ;  
   wire _dmiXbar_auto_out_1_d_ready ;  
   wire _dmiXbar_auto_out_0_a_valid ;  
   wire [2:0] _dmiXbar_auto_out_0_a_bits_opcode ;  
   wire [8:0] _dmiXbar_auto_out_0_a_bits_address ;  
   wire [31:0] _dmiXbar_auto_out_0_a_bits_data ;  
   wire _dmiXbar_auto_out_0_d_ready ;  
  TLXbar_10 dmiXbar(.clock(io_dmi_clock),.reset(io_dmi_reset),.auto_in_a_ready(_dmiXbar_auto_in_a_ready),.auto_in_a_valid(_dmi2tl_auto_out_a_valid),.auto_in_a_bits_opcode(_dmi2tl_auto_out_a_bits_opcode),.auto_in_a_bits_address(_dmi2tl_auto_out_a_bits_address),.auto_in_a_bits_data(_dmi2tl_auto_out_a_bits_data),.auto_in_d_ready(_dmi2tl_auto_out_d_ready),.auto_in_d_valid(_dmiXbar_auto_in_d_valid),.auto_in_d_bits_denied(_dmiXbar_auto_in_d_bits_denied),.auto_in_d_bits_data(_dmiXbar_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_dmiXbar_auto_in_d_bits_corrupt),.auto_out_1_a_ready(_dmOuter_auto_dmi_in_a_ready),.auto_out_1_a_valid(_dmiXbar_auto_out_1_a_valid),.auto_out_1_a_bits_opcode(_dmiXbar_auto_out_1_a_bits_opcode),.auto_out_1_a_bits_address(_dmiXbar_auto_out_1_a_bits_address),.auto_out_1_a_bits_data(_dmiXbar_auto_out_1_a_bits_data),.auto_out_1_d_ready(_dmiXbar_auto_out_1_d_ready),.auto_out_1_d_valid(_dmOuter_auto_dmi_in_d_valid),.auto_out_1_d_bits_opcode(_dmOuter_auto_dmi_in_d_bits_opcode),.auto_out_1_d_bits_data(_dmOuter_auto_dmi_in_d_bits_data),.auto_out_0_a_ready(_dmiBypass_auto_node_in_in_a_ready),.auto_out_0_a_valid(_dmiXbar_auto_out_0_a_valid),.auto_out_0_a_bits_opcode(_dmiXbar_auto_out_0_a_bits_opcode),.auto_out_0_a_bits_address(_dmiXbar_auto_out_0_a_bits_address),.auto_out_0_a_bits_data(_dmiXbar_auto_out_0_a_bits_data),.auto_out_0_d_ready(_dmiXbar_auto_out_0_d_ready),.auto_out_0_d_valid(_dmiBypass_auto_node_in_in_d_valid),.auto_out_0_d_bits_opcode(_dmiBypass_auto_node_in_in_d_bits_opcode),.auto_out_0_d_bits_param(_dmiBypass_auto_node_in_in_d_bits_param),.auto_out_0_d_bits_size(_dmiBypass_auto_node_in_in_d_bits_size),.auto_out_0_d_bits_sink(_dmiBypass_auto_node_in_in_d_bits_sink),.auto_out_0_d_bits_denied(_dmiBypass_auto_node_in_in_d_bits_denied),.auto_out_0_d_bits_data(_dmiBypass_auto_node_in_in_d_bits_data),.auto_out_0_d_bits_corrupt(_dmiBypass_auto_node_in_in_d_bits_corrupt)); 
  DMIToTL dmi2tl(.auto_out_a_ready(_dmiXbar_auto_in_a_ready),.auto_out_a_valid(_dmi2tl_auto_out_a_valid),.auto_out_a_bits_opcode(_dmi2tl_auto_out_a_bits_opcode),.auto_out_a_bits_address(_dmi2tl_auto_out_a_bits_address),.auto_out_a_bits_data(_dmi2tl_auto_out_a_bits_data),.auto_out_d_ready(_dmi2tl_auto_out_d_ready),.auto_out_d_valid(_dmiXbar_auto_in_d_valid),.auto_out_d_bits_denied(_dmiXbar_auto_in_d_bits_denied),.auto_out_d_bits_data(_dmiXbar_auto_in_d_bits_data),.auto_out_d_bits_corrupt(_dmiXbar_auto_in_d_bits_corrupt),.io_dmi_req_ready(io_dmi_req_ready),.io_dmi_req_valid(io_dmi_req_valid),.io_dmi_req_bits_addr(io_dmi_req_bits_addr),.io_dmi_req_bits_data(io_dmi_req_bits_data),.io_dmi_req_bits_op(io_dmi_req_bits_op),.io_dmi_resp_ready(io_dmi_resp_ready),.io_dmi_resp_valid(io_dmi_resp_valid),.io_dmi_resp_bits_data(io_dmi_resp_bits_data),.io_dmi_resp_bits_resp(io_dmi_resp_bits_resp)); 
  TLDebugModuleOuter dmOuter(.clock(io_dmi_clock),.reset(io_dmi_reset),.auto_dmi_in_a_ready(_dmOuter_auto_dmi_in_a_ready),.auto_dmi_in_a_valid(_dmiXbar_auto_out_1_a_valid),.auto_dmi_in_a_bits_opcode(_dmiXbar_auto_out_1_a_bits_opcode),.auto_dmi_in_a_bits_address(_dmiXbar_auto_out_1_a_bits_address),.auto_dmi_in_a_bits_data(_dmiXbar_auto_out_1_a_bits_data),.auto_dmi_in_d_ready(_dmiXbar_auto_out_1_d_ready),.auto_dmi_in_d_valid(_dmOuter_auto_dmi_in_d_valid),.auto_dmi_in_d_bits_opcode(_dmOuter_auto_dmi_in_d_bits_opcode),.auto_dmi_in_d_bits_data(_dmOuter_auto_dmi_in_d_bits_data),.auto_int_out_0(_dmOuter_auto_int_out_0),.io_ctrl_ndreset(io_ctrl_ndreset),.io_ctrl_dmactive(_dmOuter_io_ctrl_dmactive),.io_ctrl_dmactiveAck(_dmactiveAck_dmactiveAckSync_io_q),.io_innerCtrl_ready(_io_innerCtrl_source_io_enq_ready),.io_innerCtrl_valid(_dmOuter_io_innerCtrl_valid),.io_innerCtrl_bits_resumereq(_dmOuter_io_innerCtrl_bits_resumereq),.io_innerCtrl_bits_hartsel(_dmOuter_io_innerCtrl_bits_hartsel),.io_innerCtrl_bits_ackhavereset(_dmOuter_io_innerCtrl_bits_ackhavereset),.io_innerCtrl_bits_hrmask_0(_dmOuter_io_innerCtrl_bits_hrmask_0),.io_hgDebugInt_0(io_hgDebugInt_0)); 
  IntSyncCrossingSource_4 intsource(.auto_in_0(_dmOuter_auto_int_out_0),.auto_out_sync_0(auto_intsource_out_sync_0)); 
  TLBusBypass dmiBypass(.clock(io_dmi_clock),.reset(io_dmi_reset),.auto_node_out_out_a_ready(_asource_auto_in_a_ready),.auto_node_out_out_a_valid(_dmiBypass_auto_node_out_out_a_valid),.auto_node_out_out_a_bits_opcode(_dmiBypass_auto_node_out_out_a_bits_opcode),.auto_node_out_out_a_bits_address(_dmiBypass_auto_node_out_out_a_bits_address),.auto_node_out_out_a_bits_data(_dmiBypass_auto_node_out_out_a_bits_data),.auto_node_out_out_d_ready(_dmiBypass_auto_node_out_out_d_ready),.auto_node_out_out_d_valid(_asource_auto_in_d_valid),.auto_node_out_out_d_bits_opcode(_asource_auto_in_d_bits_opcode),.auto_node_out_out_d_bits_param(_asource_auto_in_d_bits_param),.auto_node_out_out_d_bits_size(_asource_auto_in_d_bits_size),.auto_node_out_out_d_bits_source(_asource_auto_in_d_bits_source),.auto_node_out_out_d_bits_sink(_asource_auto_in_d_bits_sink),.auto_node_out_out_d_bits_denied(_asource_auto_in_d_bits_denied),.auto_node_out_out_d_bits_data(_asource_auto_in_d_bits_data),.auto_node_out_out_d_bits_corrupt(_asource_auto_in_d_bits_corrupt),.auto_node_in_in_a_ready(_dmiBypass_auto_node_in_in_a_ready),.auto_node_in_in_a_valid(_dmiXbar_auto_out_0_a_valid),.auto_node_in_in_a_bits_opcode(_dmiXbar_auto_out_0_a_bits_opcode),.auto_node_in_in_a_bits_address(_dmiXbar_auto_out_0_a_bits_address),.auto_node_in_in_a_bits_data(_dmiXbar_auto_out_0_a_bits_data),.auto_node_in_in_d_ready(_dmiXbar_auto_out_0_d_ready),.auto_node_in_in_d_valid(_dmiBypass_auto_node_in_in_d_valid),.auto_node_in_in_d_bits_opcode(_dmiBypass_auto_node_in_in_d_bits_opcode),.auto_node_in_in_d_bits_param(_dmiBypass_auto_node_in_in_d_bits_param),.auto_node_in_in_d_bits_size(_dmiBypass_auto_node_in_in_d_bits_size),.auto_node_in_in_d_bits_sink(_dmiBypass_auto_node_in_in_d_bits_sink),.auto_node_in_in_d_bits_denied(_dmiBypass_auto_node_in_in_d_bits_denied),.auto_node_in_in_d_bits_data(_dmiBypass_auto_node_in_in_d_bits_data),.auto_node_in_in_d_bits_corrupt(_dmiBypass_auto_node_in_in_d_bits_corrupt),.io_bypass(~_dmOuter_io_ctrl_dmactive|~_dmactiveAck_dmactiveAckSync_io_q)); 
  TLAsyncCrossingSource asource(.clock(io_dmi_clock),.reset(io_dmi_reset),.auto_in_a_ready(_asource_auto_in_a_ready),.auto_in_a_valid(_dmiBypass_auto_node_out_out_a_valid),.auto_in_a_bits_opcode(_dmiBypass_auto_node_out_out_a_bits_opcode),.auto_in_a_bits_address(_dmiBypass_auto_node_out_out_a_bits_address),.auto_in_a_bits_data(_dmiBypass_auto_node_out_out_a_bits_data),.auto_in_d_ready(_dmiBypass_auto_node_out_out_d_ready),.auto_in_d_valid(_asource_auto_in_d_valid),.auto_in_d_bits_opcode(_asource_auto_in_d_bits_opcode),.auto_in_d_bits_param(_asource_auto_in_d_bits_param),.auto_in_d_bits_size(_asource_auto_in_d_bits_size),.auto_in_d_bits_source(_asource_auto_in_d_bits_source),.auto_in_d_bits_sink(_asource_auto_in_d_bits_sink),.auto_in_d_bits_denied(_asource_auto_in_d_bits_denied),.auto_in_d_bits_data(_asource_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_asource_auto_in_d_bits_corrupt),.auto_out_a_mem_0_opcode(auto_asource_out_a_mem_0_opcode),.auto_out_a_mem_0_address(auto_asource_out_a_mem_0_address),.auto_out_a_mem_0_data(auto_asource_out_a_mem_0_data),.auto_out_a_ridx(auto_asource_out_a_ridx),.auto_out_a_widx(auto_asource_out_a_widx),.auto_out_a_safe_ridx_valid(auto_asource_out_a_safe_ridx_valid),.auto_out_a_safe_widx_valid(auto_asource_out_a_safe_widx_valid),.auto_out_a_safe_source_reset_n(auto_asource_out_a_safe_source_reset_n),.auto_out_a_safe_sink_reset_n(auto_asource_out_a_safe_sink_reset_n),.auto_out_d_mem_0_opcode(auto_asource_out_d_mem_0_opcode),.auto_out_d_mem_0_size(auto_asource_out_d_mem_0_size),.auto_out_d_mem_0_source(auto_asource_out_d_mem_0_source),.auto_out_d_mem_0_data(auto_asource_out_d_mem_0_data),.auto_out_d_ridx(auto_asource_out_d_ridx),.auto_out_d_widx(auto_asource_out_d_widx),.auto_out_d_safe_ridx_valid(auto_asource_out_d_safe_ridx_valid),.auto_out_d_safe_widx_valid(auto_asource_out_d_safe_widx_valid),.auto_out_d_safe_source_reset_n(auto_asource_out_d_safe_source_reset_n),.auto_out_d_safe_sink_reset_n(auto_asource_out_d_safe_sink_reset_n)); 
  AsyncResetSynchronizerShiftReg_w1_d3_i0 dmactiveAck_dmactiveAckSync(.clock(io_dmi_clock),.reset(io_dmi_reset),.io_d(io_ctrl_dmactiveAck),.io_q(_dmactiveAck_dmactiveAckSync_io_q)); 
  AsyncQueueSource_1 io_innerCtrl_source(.clock(io_dmi_clock),.reset(io_dmi_reset),.io_enq_ready(_io_innerCtrl_source_io_enq_ready),.io_enq_valid(_dmOuter_io_innerCtrl_valid),.io_enq_bits_resumereq(_dmOuter_io_innerCtrl_bits_resumereq),.io_enq_bits_hartsel(_dmOuter_io_innerCtrl_bits_hartsel),.io_enq_bits_ackhavereset(_dmOuter_io_innerCtrl_bits_ackhavereset),.io_enq_bits_hrmask_0(_dmOuter_io_innerCtrl_bits_hrmask_0),.io_async_mem_resumereq_0(io_innerCtrl_mem_resumereq_0),.io_async_mem_hartsel_0(io_innerCtrl_mem_hartsel_0),.io_async_mem_ackhavereset_0(io_innerCtrl_mem_ackhavereset_0),.io_async_mem_hrmask_0_0(io_innerCtrl_mem_hrmask_0_0),.io_async_ridx(io_innerCtrl_ridx),.io_async_widx(io_innerCtrl_widx),.io_async_safe_ridx_valid(io_innerCtrl_safe_ridx_valid),.io_async_safe_widx_valid(io_innerCtrl_safe_widx_valid),.io_async_safe_source_reset_n(io_innerCtrl_safe_source_reset_n),.io_async_safe_sink_reset_n(io_innerCtrl_safe_sink_reset_n)); 
  assign io_ctrl_dmactive=_dmOuter_io_ctrl_dmactive; 
endmodule
 
module TLMonitor_33 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [1:0] io_in_a_bits_size,
  input io_in_a_bits_source,
  input [8:0] io_in_a_bits_address,
  input [3:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_size,
  input io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [1:0] size ;  
   reg source ;  
   reg [8:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] size_1 ;  
   reg source_1 ;  
   reg inflight ;  
   reg [3:0] inflight_opcodes ;  
   reg [3:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire [3:0] _GEN={1'h0,io_in_d_bits_source,2'h0} ;  
   wire [3:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire _GEN_0=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg inflight_1 ;  
   reg [3:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire [4:0] _is_aligned_mask_T_1=5'h3<<io_in_a_bits_size ;  
   wire [1:0] _GEN_1=io_in_a_bits_address[1:0]&~(_is_aligned_mask_T_1[1:0]) ;  
   wire mask_acc=io_in_a_bits_size[1]|io_in_a_bits_size[0]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_1=io_in_a_bits_size[1]|io_in_a_bits_size[0]&io_in_a_bits_address[1] ;  
   wire [3:0] mask={mask_acc_1|io_in_a_bits_address[1]&io_in_a_bits_address[0],mask_acc_1|io_in_a_bits_address[1]&~(io_in_a_bits_address[0]),mask_acc|~(io_in_a_bits_address[1])&io_in_a_bits_address[0],mask_acc|~(io_in_a_bits_address[1])&~(io_in_a_bits_address[0])} ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_3=io_in_a_bits_param>3'h2 ;  
   wire _GEN_4=io_in_a_bits_mask!=4'hF ;  
   wire _GEN_5=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_6=io_in_a_bits_size==2'h2&~io_in_a_bits_source ;  
   wire _GEN_7=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire [4:0] _GEN_8=io_in_a_bits_address[6:2]^5'h11 ;  
   wire _GEN_9=io_in_a_bits_size!=2'h3&(io_in_a_bits_address[8:6]==3'h0|{io_in_a_bits_address[8:7],_GEN_8[4:2],_GEN_8[0]}==6'h0|{io_in_a_bits_address[8:7],io_in_a_bits_address[6:3]^4'hB}==6'h0|{io_in_a_bits_address[8:7],~(io_in_a_bits_address[6:5])}==4'h0|{io_in_a_bits_address[8],~(io_in_a_bits_address[7])}==2'h0|io_in_a_bits_address[8]) ;  
   wire _GEN_10=io_in_a_bits_mask!=mask ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_15=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_16=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_18=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_19=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_20=io_in_d_valid&d_first_counter&~reset ;  
   wire _GEN_21=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_22=_GEN_21&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&~a_first_counter_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_23=_GEN_22&same_cycle_resp&~reset ;  
   wire _GEN_24=_GEN_22&~same_cycle_resp&~reset ;  
   wire [3:0] _GEN_25={2'h0,io_in_d_bits_size} ;  
   wire _GEN_26=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
   wire [3:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
   wire [3:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~(io_in_a_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~(io_in_a_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_5&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&~(_GEN_6&_GEN_9))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~(io_in_d_bits_size[1]))
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&io_in_d_bits_source)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&inflight>>io_in_a_bits_source)
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~reset&~(inflight>>io_in_d_bits_source|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_23&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&_GEN_25!={1'h0,_a_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~a_first_counter_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&~(inflight_1>>io_in_d_bits_source))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_26&_GEN_25!={1'h0,_c_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(~inflight_1|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Debug.scala:1855:19)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [30:0] _GEN_27={28'h0,io_in_d_bits_source,2'h0} ;  
   wire [30:0] _d_opcodes_clr_T_5=31'hF<<_GEN_27 ;  
   wire [18:0] _a_opcodes_set_T_1={15'h0,_GEN_0 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{16'h0,io_in_a_bits_source,2'h0} ;  
   wire [30:0] _d_sizes_clr_T_5=31'hF<<_GEN_27 ;  
   wire [17:0] _a_sizes_set_T_1={15'h0,_GEN_0 ? {io_in_a_bits_size,1'h1}:3'h0}<<{15'h0,io_in_a_bits_source,2'h0} ;  
   wire [30:0] _d_sizes_clr_T_11=31'hF<<_GEN_27 ;  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_28=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire _GEN_29=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=1'h0;
              inflight_opcodes <=4'h0;
              inflight_sizes <=4'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=1'h0;
              inflight_sizes_1 <=4'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|_GEN_0&~io_in_a_bits_source)&~(_GEN_28&~io_in_d_bits_source);
              inflight_opcodes <=(inflight_opcodes|(_GEN_0 ? _a_opcodes_set_T_1[3:0]:4'h0))&~(_GEN_28 ? _d_opcodes_clr_T_5[3:0]:4'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_0 ? _a_sizes_set_T_1[3:0]:4'h0))&~(_GEN_28 ? _d_sizes_clr_T_5[3:0]:4'h0);
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_29&~io_in_d_bits_source);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_29 ? _d_sizes_clr_T_11[3:0]:4'h0);
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module TLMonitor_34 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [1:0] io_in_a_bits_size,
  input [8:0] io_in_a_bits_source,
  input [11:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [2:0] io_in_d_bits_opcode,
  input [1:0] io_in_d_bits_size,
  input [8:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_1_out ;  
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [1:0] size ;  
   reg [8:0] source ;  
   reg [11:0] address ;  
   reg d_first_counter ;  
   reg [2:0] opcode_1 ;  
   reg [1:0] size_1 ;  
   reg [8:0] source_1 ;  
   reg [303:0] inflight ;  
   reg [1215:0] inflight_opcodes ;  
   reg [1215:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire [1215:0] _GEN={1205'h0,io_in_d_bits_source,2'h0} ;  
   wire [1215:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire _GEN_0=a_first_done&~a_first_counter_1 ;  
   wire d_release_ack=io_in_d_bits_opcode==3'h6 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   reg [303:0] inflight_1 ;  
   reg [1215:0] inflight_sizes_1 ;  
   reg d_first_counter_2 ;  
   reg [31:0] watchdog_1 ;  
   wire [5:0] _is_aligned_mask_T_1=6'h7<<io_in_a_bits_size ;  
   wire [2:0] _GEN_1=io_in_a_bits_address[2:0]&~(_is_aligned_mask_T_1[2:0]) ;  
   wire mask_size=io_in_a_bits_size==2'h2 ;  
   wire mask_acc=(&io_in_a_bits_size)|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=(&io_in_a_bits_size)|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_3=io_in_a_bits_source>9'h12F ;  
   wire _GEN_4=io_in_a_bits_param>3'h2 ;  
   wire _GEN_5=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_6=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_7=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_8=io_in_a_bits_mask!=mask ;  
   wire _GEN_9=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_14=io_in_d_valid&io_in_d_bits_opcode==3'h6&~reset ;  
   wire _GEN_15=io_in_d_bits_source>9'h12F ;  
   wire _GEN_16=io_in_d_bits_size!=2'h3 ;  
   wire _GEN_17=io_in_d_valid&io_in_d_bits_opcode==3'h4&~reset ;  
   wire _GEN_18=io_in_d_valid&io_in_d_bits_opcode==3'h5&~reset ;  
   wire _GEN_19=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_20=io_in_d_valid&d_first_counter&~reset ;  
   wire _GEN_21=io_in_d_valid&~d_first_counter_1 ;  
   wire _GEN_22=_GEN_21&~d_release_ack ;  
   wire same_cycle_resp=io_in_a_valid&~a_first_counter_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire [303:0] _GEN_23={295'h0,io_in_d_bits_source} ;  
   wire _GEN_24=_GEN_22&same_cycle_resp&~reset ;  
   wire _GEN_25=_GEN_22&~same_cycle_resp&~reset ;  
   wire [3:0] _GEN_26={2'h0,io_in_d_bits_size} ;  
   wire _GEN_27=io_in_d_valid&~d_first_counter_2&d_release_ack&~reset ;  
   wire [303:0] _GEN_28=inflight>>io_in_a_bits_source ;  
   wire [303:0] _GEN_29=inflight>>_GEN_23 ;  
   wire [1215:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
   wire [303:0] _GEN_30=inflight_1>>_GEN_23 ;  
   wire [1215:0] _c_size_lookup_T_1=inflight_sizes_1>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_9&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&(&io_in_d_bits_opcode))
            begin 
              if (1)$display("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&_GEN_16)
            begin 
              if (1)$display("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h0&~reset&_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h1&~reset&_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&io_in_d_bits_opcode==3'h2&~reset&_GEN_15)
            begin 
              if (1)$display("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_d_bits_opcode!=opcode_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_20&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&_GEN_28[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_22&~reset&~(_GEN_29[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&~(io_in_d_bits_opcode==casez_tmp|io_in_d_bits_opcode==casez_tmp_0))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_24&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&~(io_in_d_bits_opcode==casez_tmp_1|io_in_d_bits_opcode==casez_tmp_2))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_25&_GEN_26!={1'h0,_a_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_21&~a_first_counter_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~d_release_ack&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==304'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&~(_GEN_30[0]))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_27&_GEN_26!={1'h0,_c_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight_1==304'h0|_plusarg_reader_1_out==32'h0|watchdog_1<_plusarg_reader_1_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/debug/Periphery.scala:87:15)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [511:0] _GEN_31={503'h0,io_in_d_bits_source} ;  
   wire [4110:0] _GEN_32={4100'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _d_clr_T=512'h1<<_GEN_31 ;  
   wire [511:0] _a_set_T=512'h1<<io_in_a_bits_source ;  
   wire [4110:0] _d_opcodes_clr_T_5=4111'hF<<_GEN_32 ;  
   wire [4098:0] _a_opcodes_set_T_1={4095'h0,_GEN_0 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{4088'h0,io_in_a_bits_source,2'h0} ;  
   wire [4110:0] _d_sizes_clr_T_5=4111'hF<<_GEN_32 ;  
   wire [4097:0] _a_sizes_set_T_1={4095'h0,_GEN_0 ? {io_in_a_bits_size,1'h1}:3'h0}<<{4087'h0,io_in_a_bits_source,2'h0} ;  
   wire [511:0] _d_clr_T_1=512'h1<<_GEN_31 ;  
   wire [4110:0] _d_sizes_clr_T_11=4111'hF<<_GEN_32 ;  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_33=d_first_done&~d_first_counter_1&~d_release_ack ;  
   wire _GEN_34=d_first_done&~d_first_counter_2&d_release_ack ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=304'h0;
              inflight_opcodes <=1216'h0;
              inflight_sizes <=1216'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
              inflight_1 <=304'h0;
              inflight_sizes_1 <=1216'h0;
              d_first_counter_2 <=1'h0;
              watchdog_1 <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|(_GEN_0 ? _a_set_T[303:0]:304'h0))&~(_GEN_33 ? _d_clr_T[303:0]:304'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_0 ? _a_opcodes_set_T_1[1215:0]:1216'h0))&~(_GEN_33 ? _d_opcodes_clr_T_5[1215:0]:1216'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_0 ? _a_sizes_set_T_1[1215:0]:1216'h0))&~(_GEN_33 ? _d_sizes_clr_T_5[1215:0]:1216'h0);
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
              inflight_1 <=inflight_1&~(_GEN_34 ? _d_clr_T_1[303:0]:304'h0);
              inflight_sizes_1 <=inflight_sizes_1&~(_GEN_34 ? _d_sizes_clr_T_11[1215:0]:1216'h0);
              d_first_counter_2 <=(~d_first_done|d_first_counter_2-1'h1)&d_first_counter_2;
              if (d_first_done)
                 watchdog_1 <=32'h0;
               else 
                 watchdog_1 <=watchdog_1+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              opcode_1 <=io_in_d_bits_opcode;
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module TLDebugModuleInner (
  input clock,
  input reset,
  output auto_tl_in_a_ready,
  input auto_tl_in_a_valid,
  input [2:0] auto_tl_in_a_bits_opcode,
  input [2:0] auto_tl_in_a_bits_param,
  input [1:0] auto_tl_in_a_bits_size,
  input [8:0] auto_tl_in_a_bits_source,
  input [11:0] auto_tl_in_a_bits_address,
  input [7:0] auto_tl_in_a_bits_mask,
  input [63:0] auto_tl_in_a_bits_data,
  input auto_tl_in_a_bits_corrupt,
  input auto_tl_in_d_ready,
  output auto_tl_in_d_valid,
  output [2:0] auto_tl_in_d_bits_opcode,
  output [1:0] auto_tl_in_d_bits_size,
  output [8:0] auto_tl_in_d_bits_source,
  output [63:0] auto_tl_in_d_bits_data,
  output auto_dmi_in_a_ready,
  input auto_dmi_in_a_valid,
  input [2:0] auto_dmi_in_a_bits_opcode,
  input [2:0] auto_dmi_in_a_bits_param,
  input [1:0] auto_dmi_in_a_bits_size,
  input auto_dmi_in_a_bits_source,
  input [8:0] auto_dmi_in_a_bits_address,
  input [3:0] auto_dmi_in_a_bits_mask,
  input [31:0] auto_dmi_in_a_bits_data,
  input auto_dmi_in_a_bits_corrupt,
  input auto_dmi_in_d_ready,
  output auto_dmi_in_d_valid,
  output [2:0] auto_dmi_in_d_bits_opcode,
  output [1:0] auto_dmi_in_d_bits_size,
  output auto_dmi_in_d_bits_source,
  output [31:0] auto_dmi_in_d_bits_data,
  input io_dmactive,
  input io_innerCtrl_valid,
  input io_innerCtrl_bits_resumereq,
  input [9:0] io_innerCtrl_bits_hartsel,
  input io_innerCtrl_bits_ackhavereset,
  input io_innerCtrl_bits_hrmask_0,
  output io_hgDebugInt_0,
  input io_hartIsInReset_0) ; 
   wire abstractCommandBusy ;  
   wire out_woready_1_345 ;  
   wire out_woready_1_528 ;  
   wire out_woready_31 ;  
   wire out_woready_7 ;  
   wire out_woready_54 ;  
   wire out_woready_93 ;  
   wire out_woready_23 ;  
   wire out_woready_35 ;  
   wire out_woready_9 ;  
   wire out_woready_97 ;  
   wire out_woready_15 ;  
   wire out_woready_46 ;  
   wire out_woready_42 ;  
   wire out_woready_99 ;  
   wire out_woready_19 ;  
   wire out_woready_82 ;  
   wire out_woready_50 ;  
   wire out_woready_78 ;  
   wire out_woready_38 ;  
   wire out_woready_3 ;  
   wire out_woready_27 ;  
   wire _out_wofireMux_T_2 ;  
   wire out_roready_31 ;  
   wire out_roready_7 ;  
   wire out_roready_54 ;  
   wire out_roready_93 ;  
   wire out_roready_23 ;  
   wire out_roready_35 ;  
   wire out_roready_9 ;  
   wire out_roready_97 ;  
   wire out_roready_15 ;  
   wire out_roready_46 ;  
   wire out_roready_42 ;  
   wire out_roready_99 ;  
   wire out_roready_19 ;  
   wire out_roready_82 ;  
   wire out_roready_50 ;  
   wire out_roready_78 ;  
   wire out_roready_3 ;  
   wire out_roready_27 ;  
   wire out_backSel_7 ;  
   wire out_backSel_6 ;  
   wire _hartIsInResetSync_0_debug_hartReset_0_io_q ;  
   reg haltedBitRegs ;  
   reg resumeReqRegs ;  
   reg haveResetBitRegs ;  
   wire hamaskWrSel_0=io_innerCtrl_bits_hartsel==10'h0 ;  
   reg hrmaskReg_0 ;  
   reg hrDebugIntReg_0 ;  
   wire resumereq=io_innerCtrl_valid&io_innerCtrl_bits_resumereq ;  
   reg [2:0] ABSTRACTCSReg_cmderr ;  
   reg [15:0] ABSTRACTAUTOReg_autoexecprogbuf ;  
   reg [11:0] ABSTRACTAUTOReg_autoexecdata ;  
   reg [7:0] COMMANDReg_cmdtype ;  
   reg [23:0] COMMANDReg_control ;  
   reg [7:0] abstractDataMem_0 ;  
   reg [7:0] abstractDataMem_1 ;  
   reg [7:0] abstractDataMem_2 ;  
   reg [7:0] abstractDataMem_3 ;  
   reg [7:0] abstractDataMem_4 ;  
   reg [7:0] abstractDataMem_5 ;  
   reg [7:0] abstractDataMem_6 ;  
   reg [7:0] abstractDataMem_7 ;  
   reg [7:0] programBufferMem_0 ;  
   reg [7:0] programBufferMem_1 ;  
   reg [7:0] programBufferMem_2 ;  
   reg [7:0] programBufferMem_3 ;  
   reg [7:0] programBufferMem_4 ;  
   reg [7:0] programBufferMem_5 ;  
   reg [7:0] programBufferMem_6 ;  
   reg [7:0] programBufferMem_7 ;  
   reg [7:0] programBufferMem_8 ;  
   reg [7:0] programBufferMem_9 ;  
   reg [7:0] programBufferMem_10 ;  
   reg [7:0] programBufferMem_11 ;  
   reg [7:0] programBufferMem_12 ;  
   reg [7:0] programBufferMem_13 ;  
   reg [7:0] programBufferMem_14 ;  
   reg [7:0] programBufferMem_15 ;  
   reg [7:0] programBufferMem_16 ;  
   reg [7:0] programBufferMem_17 ;  
   reg [7:0] programBufferMem_18 ;  
   reg [7:0] programBufferMem_19 ;  
   reg [7:0] programBufferMem_20 ;  
   reg [7:0] programBufferMem_21 ;  
   reg [7:0] programBufferMem_22 ;  
   reg [7:0] programBufferMem_23 ;  
   reg [7:0] programBufferMem_24 ;  
   reg [7:0] programBufferMem_25 ;  
   reg [7:0] programBufferMem_26 ;  
   reg [7:0] programBufferMem_27 ;  
   reg [7:0] programBufferMem_28 ;  
   reg [7:0] programBufferMem_29 ;  
   reg [7:0] programBufferMem_30 ;  
   reg [7:0] programBufferMem_31 ;  
   reg [7:0] programBufferMem_32 ;  
   reg [7:0] programBufferMem_33 ;  
   reg [7:0] programBufferMem_34 ;  
   reg [7:0] programBufferMem_35 ;  
   reg [7:0] programBufferMem_36 ;  
   reg [7:0] programBufferMem_37 ;  
   reg [7:0] programBufferMem_38 ;  
   reg [7:0] programBufferMem_39 ;  
   reg [7:0] programBufferMem_40 ;  
   reg [7:0] programBufferMem_41 ;  
   reg [7:0] programBufferMem_42 ;  
   reg [7:0] programBufferMem_43 ;  
   reg [7:0] programBufferMem_44 ;  
   reg [7:0] programBufferMem_45 ;  
   reg [7:0] programBufferMem_46 ;  
   reg [7:0] programBufferMem_47 ;  
   reg [7:0] programBufferMem_48 ;  
   reg [7:0] programBufferMem_49 ;  
   reg [7:0] programBufferMem_50 ;  
   reg [7:0] programBufferMem_51 ;  
   reg [7:0] programBufferMem_52 ;  
   reg [7:0] programBufferMem_53 ;  
   reg [7:0] programBufferMem_54 ;  
   reg [7:0] programBufferMem_55 ;  
   reg [7:0] programBufferMem_56 ;  
   reg [7:0] programBufferMem_57 ;  
   reg [7:0] programBufferMem_58 ;  
   reg [7:0] programBufferMem_59 ;  
   reg [7:0] programBufferMem_60 ;  
   reg [7:0] programBufferMem_61 ;  
   reg [7:0] programBufferMem_62 ;  
   reg [7:0] programBufferMem_63 ;  
   wire in_bits_read=auto_dmi_in_a_bits_opcode==3'h4 ;  
   wire [1:0] _GEN={auto_dmi_in_a_bits_address[8],auto_dmi_in_a_bits_address[6]} ;  
   wire _out_T_45=_GEN==2'h0 ;  
   wire _out_T_47=_GEN==2'h1 ;  
   wire [7:0] _out_backMask_T_9={8{auto_dmi_in_a_bits_mask[2]}} ;  
   wire [7:0] _out_backMask_T_11={8{auto_dmi_in_a_bits_mask[3]}} ;  
   wire dmiAbstractDataWrEnMaybe_4=out_woready_3&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiAbstractDataWrEnMaybe_5=out_woready_3&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiAbstractDataWrEnMaybe_6=out_woready_3&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiAbstractDataWrEnMaybe_7=out_woready_3&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_56=out_woready_7&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_57=out_woready_7&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_58=out_woready_7&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_59=out_woready_7&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_36=out_woready_9&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_37=out_woready_9&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_38=out_woready_9&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_39=out_woready_9&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_28=out_woready_15&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_29=out_woready_15&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_30=out_woready_15&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_31=out_woready_15&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_12=out_woready_19&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_13=out_woready_19&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_14=out_woready_19&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_15=out_woready_19&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_44=out_woready_23&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_45=out_woready_23&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_46=out_woready_23&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_47=out_woready_23&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiAbstractDataWrEnMaybe_0=out_woready_27&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiAbstractDataWrEnMaybe_1=out_woready_27&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiAbstractDataWrEnMaybe_2=out_woready_27&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiAbstractDataWrEnMaybe_3=out_woready_27&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_60=out_woready_31&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_61=out_woready_31&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_62=out_woready_31&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_63=out_woready_31&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_40=out_woready_35&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_41=out_woready_35&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_42=out_woready_35&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_43=out_woready_35&auto_dmi_in_a_bits_mask[3] ;  
   wire autoexecdataWrEnMaybe=out_woready_38&auto_dmi_in_a_bits_mask[0] ;  
   wire autoexecprogbufWrEnMaybe=out_woready_38&(&{_out_backMask_T_11,_out_backMask_T_9}) ;  
   wire dmiProgramBufferWrEnMaybe_20=out_woready_42&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_21=out_woready_42&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_22=out_woready_42&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_23=out_woready_42&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_24=out_woready_46&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_25=out_woready_46&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_26=out_woready_46&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_27=out_woready_46&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_4=out_woready_50&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_5=out_woready_50&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_6=out_woready_50&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_7=out_woready_50&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_52=out_woready_54&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_53=out_woready_54&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_54=out_woready_54&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_55=out_woready_54&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_0=out_woready_78&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_1=out_woready_78&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_2=out_woready_78&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_3=out_woready_78&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_8=out_woready_82&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_9=out_woready_82&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_10=out_woready_82&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_11=out_woready_82&auto_dmi_in_a_bits_mask[3] ;  
   wire ABSTRACTCSWrEnMaybe=_out_wofireMux_T_2&out_backSel_6&_out_T_47&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_48=out_woready_93&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_49=out_woready_93&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_50=out_woready_93&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_51=out_woready_93&auto_dmi_in_a_bits_mask[3] ;  
   wire dmiProgramBufferWrEnMaybe_32=out_woready_97&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_33=out_woready_97&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_34=out_woready_97&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_35=out_woready_97&auto_dmi_in_a_bits_mask[3] ;  
   wire COMMANDWrEnMaybe=_out_wofireMux_T_2&out_backSel_7&_out_T_47&(&{_out_backMask_T_11,_out_backMask_T_9,{8{auto_dmi_in_a_bits_mask[1]}},{8{auto_dmi_in_a_bits_mask[0]}}}) ;  
   wire [31:0] COMMANDWrDataVal=COMMANDWrEnMaybe ? auto_dmi_in_a_bits_data:32'h0 ;  
   wire dmiProgramBufferWrEnMaybe_16=out_woready_99&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferWrEnMaybe_17=out_woready_99&auto_dmi_in_a_bits_mask[1] ;  
   wire dmiProgramBufferWrEnMaybe_18=out_woready_99&auto_dmi_in_a_bits_mask[2] ;  
   wire dmiProgramBufferWrEnMaybe_19=out_woready_99&auto_dmi_in_a_bits_mask[3] ;  
   wire [4:0] out_oindex={auto_dmi_in_a_bits_address[7],auto_dmi_in_a_bits_address[5:2]} ;  
   wire [4:0] _GEN_0={auto_dmi_in_a_bits_address[7],auto_dmi_in_a_bits_address[5:2]} ;  
   wire out_backSel_4=_GEN_0==5'h4 ;  
   wire out_backSel_5=_GEN_0==5'h5 ;  
  assign out_backSel_6=_GEN_0==5'h6; 
  assign out_backSel_7=_GEN_0==5'h7; 
   wire out_backSel_16=_GEN_0==5'h10 ;  
   wire out_backSel_17=_GEN_0==5'h11 ;  
   wire out_backSel_18=_GEN_0==5'h12 ;  
   wire out_backSel_19=_GEN_0==5'h13 ;  
   wire out_backSel_20=_GEN_0==5'h14 ;  
   wire out_backSel_21=_GEN_0==5'h15 ;  
   wire out_backSel_22=_GEN_0==5'h16 ;  
   wire out_backSel_23=_GEN_0==5'h17 ;  
   wire out_backSel_24=_GEN_0==5'h18 ;  
   wire out_backSel_25=_GEN_0==5'h19 ;  
   wire out_backSel_26=_GEN_0==5'h1A ;  
   wire out_backSel_27=_GEN_0==5'h1B ;  
   wire out_backSel_28=_GEN_0==5'h1C ;  
   wire out_backSel_29=_GEN_0==5'h1D ;  
   wire out_backSel_30=_GEN_0==5'h1E ;  
   wire _out_wofireMux_T=auto_dmi_in_a_valid&auto_dmi_in_d_ready ;  
   wire _out_rofireMux_T_1=_out_wofireMux_T&in_bits_read ;  
  assign out_roready_27=_out_rofireMux_T_1&out_backSel_4&_out_T_45; 
  assign out_roready_3=_out_rofireMux_T_1&out_backSel_5&_out_T_45; 
  assign out_roready_78=_out_rofireMux_T_1&out_backSel_16&_out_T_45; 
  assign out_roready_50=_out_rofireMux_T_1&out_backSel_17&_out_T_45; 
  assign out_roready_82=_out_rofireMux_T_1&out_backSel_18&_out_T_45; 
  assign out_roready_19=_out_rofireMux_T_1&out_backSel_19&_out_T_45; 
  assign out_roready_99=_out_rofireMux_T_1&out_backSel_20&_out_T_45; 
  assign out_roready_42=_out_rofireMux_T_1&out_backSel_21&_out_T_45; 
  assign out_roready_46=_out_rofireMux_T_1&out_backSel_22&_out_T_45; 
  assign out_roready_15=_out_rofireMux_T_1&out_backSel_23&_out_T_45; 
  assign out_roready_97=_out_rofireMux_T_1&out_backSel_24&_out_T_45; 
  assign out_roready_9=_out_rofireMux_T_1&out_backSel_25&_out_T_45; 
  assign out_roready_35=_out_rofireMux_T_1&out_backSel_26&_out_T_45; 
  assign out_roready_23=_out_rofireMux_T_1&out_backSel_27&_out_T_45; 
  assign out_roready_93=_out_rofireMux_T_1&out_backSel_28&_out_T_45; 
  assign out_roready_54=_out_rofireMux_T_1&out_backSel_29&_out_T_45; 
  assign out_roready_7=_out_rofireMux_T_1&out_backSel_30&_out_T_45; 
  assign out_roready_31=_out_rofireMux_T_1&(&_GEN_0)&_out_T_45; 
  assign _out_wofireMux_T_2=_out_wofireMux_T&~in_bits_read; 
  assign out_woready_27=_out_wofireMux_T_2&out_backSel_4&_out_T_45; 
  assign out_woready_3=_out_wofireMux_T_2&out_backSel_5&_out_T_45; 
  assign out_woready_38=_out_wofireMux_T_2&_GEN_0==5'h8&_out_T_47; 
  assign out_woready_78=_out_wofireMux_T_2&out_backSel_16&_out_T_45; 
  assign out_woready_50=_out_wofireMux_T_2&out_backSel_17&_out_T_45; 
  assign out_woready_82=_out_wofireMux_T_2&out_backSel_18&_out_T_45; 
  assign out_woready_19=_out_wofireMux_T_2&out_backSel_19&_out_T_45; 
  assign out_woready_99=_out_wofireMux_T_2&out_backSel_20&_out_T_45; 
  assign out_woready_42=_out_wofireMux_T_2&out_backSel_21&_out_T_45; 
  assign out_woready_46=_out_wofireMux_T_2&out_backSel_22&_out_T_45; 
  assign out_woready_15=_out_wofireMux_T_2&out_backSel_23&_out_T_45; 
  assign out_woready_97=_out_wofireMux_T_2&out_backSel_24&_out_T_45; 
  assign out_woready_9=_out_wofireMux_T_2&out_backSel_25&_out_T_45; 
  assign out_woready_35=_out_wofireMux_T_2&out_backSel_26&_out_T_45; 
  assign out_woready_23=_out_wofireMux_T_2&out_backSel_27&_out_T_45; 
  assign out_woready_93=_out_wofireMux_T_2&out_backSel_28&_out_T_45; 
  assign out_woready_54=_out_wofireMux_T_2&out_backSel_29&_out_T_45; 
  assign out_woready_7=_out_wofireMux_T_2&out_backSel_30&_out_T_45; 
  assign out_woready_31=_out_wofireMux_T_2&(&_GEN_0)&_out_T_45; 
   reg casez_tmp ;  
  always @(*)
       begin 
         casez (out_oindex)
          5 'b00000:
             casez_tmp =_GEN==2'h2;
          5 'b00001:
             casez_tmp =_out_T_47;
          5 'b00010:
             casez_tmp =1'h1;
          5 'b00011:
             casez_tmp =_out_T_47;
          5 'b00100:
             casez_tmp =_out_T_45;
          5 'b00101:
             casez_tmp =_out_T_45;
          5 'b00110:
             casez_tmp =_out_T_47;
          5 'b00111:
             casez_tmp =_out_T_47;
          5 'b01000:
             casez_tmp =_out_T_47;
          5 'b01001:
             casez_tmp =1'h1;
          5 'b01010:
             casez_tmp =1'h1;
          5 'b01011:
             casez_tmp =1'h1;
          5 'b01100:
             casez_tmp =1'h1;
          5 'b01101:
             casez_tmp =1'h1;
          5 'b01110:
             casez_tmp =1'h1;
          5 'b01111:
             casez_tmp =1'h1;
          5 'b10000:
             casez_tmp =_out_T_45;
          5 'b10001:
             casez_tmp =_out_T_45;
          5 'b10010:
             casez_tmp =_out_T_45;
          5 'b10011:
             casez_tmp =_out_T_45;
          5 'b10100:
             casez_tmp =_out_T_45;
          5 'b10101:
             casez_tmp =_out_T_45;
          5 'b10110:
             casez_tmp =_out_T_45;
          5 'b10111:
             casez_tmp =_out_T_45;
          5 'b11000:
             casez_tmp =_out_T_45;
          5 'b11001:
             casez_tmp =_out_T_45;
          5 'b11010:
             casez_tmp =_out_T_45;
          5 'b11011:
             casez_tmp =_out_T_45;
          5 'b11100:
             casez_tmp =_out_T_45;
          5 'b11101:
             casez_tmp =_out_T_45;
          5 'b11110:
             casez_tmp =_out_T_45;
          default :
             casez_tmp =_out_T_45;
         endcase 
       end
  
   reg [31:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (out_oindex)
          5 'b00000:
             casez_tmp_0 ={31'h0,haltedBitRegs};
          5 'b00001:
             casez_tmp_0 ={12'h0,{2{haveResetBitRegs}},{2{resumereq ? ~resumeReqRegs&~hamaskWrSel_0:~resumeReqRegs}},4'h0,~haltedBitRegs,~haltedBitRegs,{2{haltedBitRegs}},8'hA2};
          5 'b00010:
             casez_tmp_0 =32'h0;
          5 'b00011:
             casez_tmp_0 ={31'h0,haltedBitRegs};
          5 'b00100:
             casez_tmp_0 ={abstractDataMem_3,abstractDataMem_2,abstractDataMem_1,abstractDataMem_0};
          5 'b00101:
             casez_tmp_0 ={abstractDataMem_7,abstractDataMem_6,abstractDataMem_5,abstractDataMem_4};
          5 'b00110:
             casez_tmp_0 ={19'h8000,abstractCommandBusy,1'h0,ABSTRACTCSReg_cmderr,8'h2};
          5 'b00111:
             casez_tmp_0 ={COMMANDReg_cmdtype,COMMANDReg_control};
          5 'b01000:
             casez_tmp_0 ={ABSTRACTAUTOReg_autoexecprogbuf,14'h0,ABSTRACTAUTOReg_autoexecdata[1:0]};
          5 'b01001:
             casez_tmp_0 =32'h0;
          5 'b01010:
             casez_tmp_0 =32'h0;
          5 'b01011:
             casez_tmp_0 =32'h0;
          5 'b01100:
             casez_tmp_0 =32'h0;
          5 'b01101:
             casez_tmp_0 =32'h0;
          5 'b01110:
             casez_tmp_0 =32'h0;
          5 'b01111:
             casez_tmp_0 =32'h0;
          5 'b10000:
             casez_tmp_0 ={programBufferMem_3,programBufferMem_2,programBufferMem_1,programBufferMem_0};
          5 'b10001:
             casez_tmp_0 ={programBufferMem_7,programBufferMem_6,programBufferMem_5,programBufferMem_4};
          5 'b10010:
             casez_tmp_0 ={programBufferMem_11,programBufferMem_10,programBufferMem_9,programBufferMem_8};
          5 'b10011:
             casez_tmp_0 ={programBufferMem_15,programBufferMem_14,programBufferMem_13,programBufferMem_12};
          5 'b10100:
             casez_tmp_0 ={programBufferMem_19,programBufferMem_18,programBufferMem_17,programBufferMem_16};
          5 'b10101:
             casez_tmp_0 ={programBufferMem_23,programBufferMem_22,programBufferMem_21,programBufferMem_20};
          5 'b10110:
             casez_tmp_0 ={programBufferMem_27,programBufferMem_26,programBufferMem_25,programBufferMem_24};
          5 'b10111:
             casez_tmp_0 ={programBufferMem_31,programBufferMem_30,programBufferMem_29,programBufferMem_28};
          5 'b11000:
             casez_tmp_0 ={programBufferMem_35,programBufferMem_34,programBufferMem_33,programBufferMem_32};
          5 'b11001:
             casez_tmp_0 ={programBufferMem_39,programBufferMem_38,programBufferMem_37,programBufferMem_36};
          5 'b11010:
             casez_tmp_0 ={programBufferMem_43,programBufferMem_42,programBufferMem_41,programBufferMem_40};
          5 'b11011:
             casez_tmp_0 ={programBufferMem_47,programBufferMem_46,programBufferMem_45,programBufferMem_44};
          5 'b11100:
             casez_tmp_0 ={programBufferMem_51,programBufferMem_50,programBufferMem_49,programBufferMem_48};
          5 'b11101:
             casez_tmp_0 ={programBufferMem_55,programBufferMem_54,programBufferMem_53,programBufferMem_52};
          5 'b11110:
             casez_tmp_0 ={programBufferMem_59,programBufferMem_58,programBufferMem_57,programBufferMem_56};
          default :
             casez_tmp_0 ={programBufferMem_63,programBufferMem_62,programBufferMem_61,programBufferMem_60};
         endcase 
       end
  
   wire [2:0] dmiNodeIn_d_bits_opcode={2'h0,in_bits_read} ;  
   reg goReg ;  
   reg [31:0] abstractGeneratedMem_0 ;  
   reg [31:0] abstractGeneratedMem_1 ;  
   wire in_1_bits_read=auto_tl_in_a_bits_opcode==3'h4 ;  
   wire [9:0] _out_womask_T_631={{2{auto_tl_in_a_bits_mask[1]}},{8{auto_tl_in_a_bits_mask[0]}}} ;  
   wire hartResumingWrEn=out_woready_1_345&(&_out_womask_T_631) ;  
   wire [9:0] _out_womask_T_632={{2{auto_tl_in_a_bits_mask[5]}},{8{auto_tl_in_a_bits_mask[4]}}} ;  
   wire hartExceptionWrEn=out_woready_1_345&(&_out_womask_T_632) ;  
   wire hartHaltedWrEn=out_woready_1_528&(&_out_womask_T_631) ;  
   wire hartGoingWrEn=out_woready_1_528&(&_out_womask_T_632) ;  
   wire _out_wofireMux_T_134=auto_tl_in_a_valid&auto_tl_in_d_ready&~in_1_bits_read ;  
  assign out_woready_1_528=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h20&~(auto_tl_in_a_bits_address[11]); 
  assign out_woready_1_345=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h21&~(auto_tl_in_a_bits_address[11]); 
   wire out_woready_1_922=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h68&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_510=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h69&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_191=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h6A&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_1074=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h6B&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_722=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h6C&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_442=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h6D&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_111=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h6E&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_1146=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h6F&~(auto_tl_in_a_bits_address[11]) ;  
   wire out_woready_1_818=_out_wofireMux_T_134&auto_tl_in_a_bits_address[10:3]==8'h70&~(auto_tl_in_a_bits_address[11]) ;  
   reg casez_tmp_1 ;  
  always @(*)
       begin 
         casez (auto_tl_in_a_bits_address[10:3])
          8 'b00000000:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00000001:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00000010:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00000011:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00000100:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00000101:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00000110:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00000111:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00001000:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00001001:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00001010:
             casez_tmp_1 =auto_tl_in_a_bits_address[11];
          8 'b00001011:
             casez_tmp_1 =1'h1;
          8 'b00001100:
             casez_tmp_1 =1'h1;
          8 'b00001101:
             casez_tmp_1 =1'h1;
          8 'b00001110:
             casez_tmp_1 =1'h1;
          8 'b00001111:
             casez_tmp_1 =1'h1;
          8 'b00010000:
             casez_tmp_1 =1'h1;
          8 'b00010001:
             casez_tmp_1 =1'h1;
          8 'b00010010:
             casez_tmp_1 =1'h1;
          8 'b00010011:
             casez_tmp_1 =1'h1;
          8 'b00010100:
             casez_tmp_1 =1'h1;
          8 'b00010101:
             casez_tmp_1 =1'h1;
          8 'b00010110:
             casez_tmp_1 =1'h1;
          8 'b00010111:
             casez_tmp_1 =1'h1;
          8 'b00011000:
             casez_tmp_1 =1'h1;
          8 'b00011001:
             casez_tmp_1 =1'h1;
          8 'b00011010:
             casez_tmp_1 =1'h1;
          8 'b00011011:
             casez_tmp_1 =1'h1;
          8 'b00011100:
             casez_tmp_1 =1'h1;
          8 'b00011101:
             casez_tmp_1 =1'h1;
          8 'b00011110:
             casez_tmp_1 =1'h1;
          8 'b00011111:
             casez_tmp_1 =1'h1;
          8 'b00100000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b00100001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b00100010:
             casez_tmp_1 =1'h1;
          8 'b00100011:
             casez_tmp_1 =1'h1;
          8 'b00100100:
             casez_tmp_1 =1'h1;
          8 'b00100101:
             casez_tmp_1 =1'h1;
          8 'b00100110:
             casez_tmp_1 =1'h1;
          8 'b00100111:
             casez_tmp_1 =1'h1;
          8 'b00101000:
             casez_tmp_1 =1'h1;
          8 'b00101001:
             casez_tmp_1 =1'h1;
          8 'b00101010:
             casez_tmp_1 =1'h1;
          8 'b00101011:
             casez_tmp_1 =1'h1;
          8 'b00101100:
             casez_tmp_1 =1'h1;
          8 'b00101101:
             casez_tmp_1 =1'h1;
          8 'b00101110:
             casez_tmp_1 =1'h1;
          8 'b00101111:
             casez_tmp_1 =1'h1;
          8 'b00110000:
             casez_tmp_1 =1'h1;
          8 'b00110001:
             casez_tmp_1 =1'h1;
          8 'b00110010:
             casez_tmp_1 =1'h1;
          8 'b00110011:
             casez_tmp_1 =1'h1;
          8 'b00110100:
             casez_tmp_1 =1'h1;
          8 'b00110101:
             casez_tmp_1 =1'h1;
          8 'b00110110:
             casez_tmp_1 =1'h1;
          8 'b00110111:
             casez_tmp_1 =1'h1;
          8 'b00111000:
             casez_tmp_1 =1'h1;
          8 'b00111001:
             casez_tmp_1 =1'h1;
          8 'b00111010:
             casez_tmp_1 =1'h1;
          8 'b00111011:
             casez_tmp_1 =1'h1;
          8 'b00111100:
             casez_tmp_1 =1'h1;
          8 'b00111101:
             casez_tmp_1 =1'h1;
          8 'b00111110:
             casez_tmp_1 =1'h1;
          8 'b00111111:
             casez_tmp_1 =1'h1;
          8 'b01000000:
             casez_tmp_1 =1'h1;
          8 'b01000001:
             casez_tmp_1 =1'h1;
          8 'b01000010:
             casez_tmp_1 =1'h1;
          8 'b01000011:
             casez_tmp_1 =1'h1;
          8 'b01000100:
             casez_tmp_1 =1'h1;
          8 'b01000101:
             casez_tmp_1 =1'h1;
          8 'b01000110:
             casez_tmp_1 =1'h1;
          8 'b01000111:
             casez_tmp_1 =1'h1;
          8 'b01001000:
             casez_tmp_1 =1'h1;
          8 'b01001001:
             casez_tmp_1 =1'h1;
          8 'b01001010:
             casez_tmp_1 =1'h1;
          8 'b01001011:
             casez_tmp_1 =1'h1;
          8 'b01001100:
             casez_tmp_1 =1'h1;
          8 'b01001101:
             casez_tmp_1 =1'h1;
          8 'b01001110:
             casez_tmp_1 =1'h1;
          8 'b01001111:
             casez_tmp_1 =1'h1;
          8 'b01010000:
             casez_tmp_1 =1'h1;
          8 'b01010001:
             casez_tmp_1 =1'h1;
          8 'b01010010:
             casez_tmp_1 =1'h1;
          8 'b01010011:
             casez_tmp_1 =1'h1;
          8 'b01010100:
             casez_tmp_1 =1'h1;
          8 'b01010101:
             casez_tmp_1 =1'h1;
          8 'b01010110:
             casez_tmp_1 =1'h1;
          8 'b01010111:
             casez_tmp_1 =1'h1;
          8 'b01011000:
             casez_tmp_1 =1'h1;
          8 'b01011001:
             casez_tmp_1 =1'h1;
          8 'b01011010:
             casez_tmp_1 =1'h1;
          8 'b01011011:
             casez_tmp_1 =1'h1;
          8 'b01011100:
             casez_tmp_1 =1'h1;
          8 'b01011101:
             casez_tmp_1 =1'h1;
          8 'b01011110:
             casez_tmp_1 =1'h1;
          8 'b01011111:
             casez_tmp_1 =1'h1;
          8 'b01100000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01100001:
             casez_tmp_1 =1'h1;
          8 'b01100010:
             casez_tmp_1 =1'h1;
          8 'b01100011:
             casez_tmp_1 =1'h1;
          8 'b01100100:
             casez_tmp_1 =1'h1;
          8 'b01100101:
             casez_tmp_1 =1'h1;
          8 'b01100110:
             casez_tmp_1 =1'h1;
          8 'b01100111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01101111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01110000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b01110001:
             casez_tmp_1 =1'h1;
          8 'b01110010:
             casez_tmp_1 =1'h1;
          8 'b01110011:
             casez_tmp_1 =1'h1;
          8 'b01110100:
             casez_tmp_1 =1'h1;
          8 'b01110101:
             casez_tmp_1 =1'h1;
          8 'b01110110:
             casez_tmp_1 =1'h1;
          8 'b01110111:
             casez_tmp_1 =1'h1;
          8 'b01111000:
             casez_tmp_1 =1'h1;
          8 'b01111001:
             casez_tmp_1 =1'h1;
          8 'b01111010:
             casez_tmp_1 =1'h1;
          8 'b01111011:
             casez_tmp_1 =1'h1;
          8 'b01111100:
             casez_tmp_1 =1'h1;
          8 'b01111101:
             casez_tmp_1 =1'h1;
          8 'b01111110:
             casez_tmp_1 =1'h1;
          8 'b01111111:
             casez_tmp_1 =1'h1;
          8 'b10000000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10000001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10000010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10000011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10000100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10000101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10000110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10000111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10001111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10010111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10011111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10100111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10101111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10110111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b10111111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11000111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11001111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11010111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11011111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11100111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11101111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11110111:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11111000:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11111001:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11111010:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11111011:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11111100:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11111101:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          8 'b11111110:
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
          default :
             casez_tmp_1 =~(auto_tl_in_a_bits_address[11]);
         endcase 
       end
  
   reg [63:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (auto_tl_in_a_bits_address[10:3])
          8 'b00000000:
             casez_tmp_2 =64'h380006F00C0006F;
          8 'b00000001:
             casez_tmp_2 =64'hFF0000F0440006F;
          8 'b00000010:
             casez_tmp_2 =64'hF14024737B241073;
          8 'b00000011:
             casez_tmp_2 =64'h4004440310802023;
          8 'b00000100:
             casez_tmp_2 =64'hFE0408E300347413;
          8 'b00000101:
             casez_tmp_2 =64'h4086300147413;
          8 'b00000110:
             casez_tmp_2 =64'h100022237B202473;
          8 'b00000111:
             casez_tmp_2 =64'hF140247330000067;
          8 'b00001000:
             casez_tmp_2 =64'h7B20247310802423;
          8 'b00001001:
             casez_tmp_2 =64'h100026237B200073;
          8 'b00001010:
             casez_tmp_2 =64'h100073;
          8 'b00001011:
             casez_tmp_2 =64'h0;
          8 'b00001100:
             casez_tmp_2 =64'h0;
          8 'b00001101:
             casez_tmp_2 =64'h0;
          8 'b00001110:
             casez_tmp_2 =64'h0;
          8 'b00001111:
             casez_tmp_2 =64'h0;
          8 'b00010000:
             casez_tmp_2 =64'h0;
          8 'b00010001:
             casez_tmp_2 =64'h0;
          8 'b00010010:
             casez_tmp_2 =64'h0;
          8 'b00010011:
             casez_tmp_2 =64'h0;
          8 'b00010100:
             casez_tmp_2 =64'h0;
          8 'b00010101:
             casez_tmp_2 =64'h0;
          8 'b00010110:
             casez_tmp_2 =64'h0;
          8 'b00010111:
             casez_tmp_2 =64'h0;
          8 'b00011000:
             casez_tmp_2 =64'h0;
          8 'b00011001:
             casez_tmp_2 =64'h0;
          8 'b00011010:
             casez_tmp_2 =64'h0;
          8 'b00011011:
             casez_tmp_2 =64'h0;
          8 'b00011100:
             casez_tmp_2 =64'h0;
          8 'b00011101:
             casez_tmp_2 =64'h0;
          8 'b00011110:
             casez_tmp_2 =64'h0;
          8 'b00011111:
             casez_tmp_2 =64'h0;
          8 'b00100000:
             casez_tmp_2 =64'h0;
          8 'b00100001:
             casez_tmp_2 =64'h0;
          8 'b00100010:
             casez_tmp_2 =64'h0;
          8 'b00100011:
             casez_tmp_2 =64'h0;
          8 'b00100100:
             casez_tmp_2 =64'h0;
          8 'b00100101:
             casez_tmp_2 =64'h0;
          8 'b00100110:
             casez_tmp_2 =64'h0;
          8 'b00100111:
             casez_tmp_2 =64'h0;
          8 'b00101000:
             casez_tmp_2 =64'h0;
          8 'b00101001:
             casez_tmp_2 =64'h0;
          8 'b00101010:
             casez_tmp_2 =64'h0;
          8 'b00101011:
             casez_tmp_2 =64'h0;
          8 'b00101100:
             casez_tmp_2 =64'h0;
          8 'b00101101:
             casez_tmp_2 =64'h0;
          8 'b00101110:
             casez_tmp_2 =64'h0;
          8 'b00101111:
             casez_tmp_2 =64'h0;
          8 'b00110000:
             casez_tmp_2 =64'h0;
          8 'b00110001:
             casez_tmp_2 =64'h0;
          8 'b00110010:
             casez_tmp_2 =64'h0;
          8 'b00110011:
             casez_tmp_2 =64'h0;
          8 'b00110100:
             casez_tmp_2 =64'h0;
          8 'b00110101:
             casez_tmp_2 =64'h0;
          8 'b00110110:
             casez_tmp_2 =64'h0;
          8 'b00110111:
             casez_tmp_2 =64'h0;
          8 'b00111000:
             casez_tmp_2 =64'h0;
          8 'b00111001:
             casez_tmp_2 =64'h0;
          8 'b00111010:
             casez_tmp_2 =64'h0;
          8 'b00111011:
             casez_tmp_2 =64'h0;
          8 'b00111100:
             casez_tmp_2 =64'h0;
          8 'b00111101:
             casez_tmp_2 =64'h0;
          8 'b00111110:
             casez_tmp_2 =64'h0;
          8 'b00111111:
             casez_tmp_2 =64'h0;
          8 'b01000000:
             casez_tmp_2 =64'h0;
          8 'b01000001:
             casez_tmp_2 =64'h0;
          8 'b01000010:
             casez_tmp_2 =64'h0;
          8 'b01000011:
             casez_tmp_2 =64'h0;
          8 'b01000100:
             casez_tmp_2 =64'h0;
          8 'b01000101:
             casez_tmp_2 =64'h0;
          8 'b01000110:
             casez_tmp_2 =64'h0;
          8 'b01000111:
             casez_tmp_2 =64'h0;
          8 'b01001000:
             casez_tmp_2 =64'h0;
          8 'b01001001:
             casez_tmp_2 =64'h0;
          8 'b01001010:
             casez_tmp_2 =64'h0;
          8 'b01001011:
             casez_tmp_2 =64'h0;
          8 'b01001100:
             casez_tmp_2 =64'h0;
          8 'b01001101:
             casez_tmp_2 =64'h0;
          8 'b01001110:
             casez_tmp_2 =64'h0;
          8 'b01001111:
             casez_tmp_2 =64'h0;
          8 'b01010000:
             casez_tmp_2 =64'h0;
          8 'b01010001:
             casez_tmp_2 =64'h0;
          8 'b01010010:
             casez_tmp_2 =64'h0;
          8 'b01010011:
             casez_tmp_2 =64'h0;
          8 'b01010100:
             casez_tmp_2 =64'h0;
          8 'b01010101:
             casez_tmp_2 =64'h0;
          8 'b01010110:
             casez_tmp_2 =64'h0;
          8 'b01010111:
             casez_tmp_2 =64'h0;
          8 'b01011000:
             casez_tmp_2 =64'h0;
          8 'b01011001:
             casez_tmp_2 =64'h0;
          8 'b01011010:
             casez_tmp_2 =64'h0;
          8 'b01011011:
             casez_tmp_2 =64'h0;
          8 'b01011100:
             casez_tmp_2 =64'h0;
          8 'b01011101:
             casez_tmp_2 =64'h0;
          8 'b01011110:
             casez_tmp_2 =64'h0;
          8 'b01011111:
             casez_tmp_2 =64'h0;
          8 'b01100000:
             casez_tmp_2 =64'h380006F;
          8 'b01100001:
             casez_tmp_2 =64'h0;
          8 'b01100010:
             casez_tmp_2 =64'h0;
          8 'b01100011:
             casez_tmp_2 =64'h0;
          8 'b01100100:
             casez_tmp_2 =64'h0;
          8 'b01100101:
             casez_tmp_2 =64'h0;
          8 'b01100110:
             casez_tmp_2 =64'h0;
          8 'b01100111:
             casez_tmp_2 ={abstractGeneratedMem_1,abstractGeneratedMem_0};
          8 'b01101000:
             casez_tmp_2 ={programBufferMem_7,programBufferMem_6,programBufferMem_5,programBufferMem_4,programBufferMem_3,programBufferMem_2,programBufferMem_1,programBufferMem_0};
          8 'b01101001:
             casez_tmp_2 ={programBufferMem_15,programBufferMem_14,programBufferMem_13,programBufferMem_12,programBufferMem_11,programBufferMem_10,programBufferMem_9,programBufferMem_8};
          8 'b01101010:
             casez_tmp_2 ={programBufferMem_23,programBufferMem_22,programBufferMem_21,programBufferMem_20,programBufferMem_19,programBufferMem_18,programBufferMem_17,programBufferMem_16};
          8 'b01101011:
             casez_tmp_2 ={programBufferMem_31,programBufferMem_30,programBufferMem_29,programBufferMem_28,programBufferMem_27,programBufferMem_26,programBufferMem_25,programBufferMem_24};
          8 'b01101100:
             casez_tmp_2 ={programBufferMem_39,programBufferMem_38,programBufferMem_37,programBufferMem_36,programBufferMem_35,programBufferMem_34,programBufferMem_33,programBufferMem_32};
          8 'b01101101:
             casez_tmp_2 ={programBufferMem_47,programBufferMem_46,programBufferMem_45,programBufferMem_44,programBufferMem_43,programBufferMem_42,programBufferMem_41,programBufferMem_40};
          8 'b01101110:
             casez_tmp_2 ={programBufferMem_55,programBufferMem_54,programBufferMem_53,programBufferMem_52,programBufferMem_51,programBufferMem_50,programBufferMem_49,programBufferMem_48};
          8 'b01101111:
             casez_tmp_2 ={programBufferMem_63,programBufferMem_62,programBufferMem_61,programBufferMem_60,programBufferMem_59,programBufferMem_58,programBufferMem_57,programBufferMem_56};
          8 'b01110000:
             casez_tmp_2 ={abstractDataMem_7,abstractDataMem_6,abstractDataMem_5,abstractDataMem_4,abstractDataMem_3,abstractDataMem_2,abstractDataMem_1,abstractDataMem_0};
          8 'b01110001:
             casez_tmp_2 =64'h0;
          8 'b01110010:
             casez_tmp_2 =64'h0;
          8 'b01110011:
             casez_tmp_2 =64'h0;
          8 'b01110100:
             casez_tmp_2 =64'h0;
          8 'b01110101:
             casez_tmp_2 =64'h0;
          8 'b01110110:
             casez_tmp_2 =64'h0;
          8 'b01110111:
             casez_tmp_2 =64'h0;
          8 'b01111000:
             casez_tmp_2 =64'h0;
          8 'b01111001:
             casez_tmp_2 =64'h0;
          8 'b01111010:
             casez_tmp_2 =64'h0;
          8 'b01111011:
             casez_tmp_2 =64'h0;
          8 'b01111100:
             casez_tmp_2 =64'h0;
          8 'b01111101:
             casez_tmp_2 =64'h0;
          8 'b01111110:
             casez_tmp_2 =64'h0;
          8 'b01111111:
             casez_tmp_2 =64'h0;
          8 'b10000000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10000001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10000010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10000011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10000100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10000101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10000110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10000111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10001111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10010111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10011111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10100111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10101111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10110111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b10111111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11000111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11001111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11010111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11011111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11100111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11101111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11110111:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11111000:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11111001:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11111010:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11111011:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11111100:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11111101:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          8 'b11111110:
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
          default :
             casez_tmp_2 ={6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg,6'h0,resumeReqRegs,goReg};
         endcase 
       end
  
   wire [2:0] tlNodeIn_d_bits_opcode={2'h0,in_1_bits_read} ;  
   reg [1:0] ctrlStateReg ;  
  assign abstractCommandBusy=|ctrlStateReg; 
   wire commandRegIsAccessRegister=COMMANDReg_cmdtype==8'h0 ;  
   wire _GEN_1=~(COMMANDReg_control[17])|(|(COMMANDReg_control[15:12]))&COMMANDReg_control[15:0]<16'h1020&(COMMANDReg_control[22:20]==3'h2|COMMANDReg_control[22:20]==3'h3) ;  
   wire commandRegIsUnsupported=~commandRegIsAccessRegister|~_GEN_1 ;  
   wire commandRegBadHaltResume=commandRegIsAccessRegister&_GEN_1&~haltedBitRegs ;  
   wire _GEN_2=ctrlStateReg==2'h1 ;  
   wire _GEN_3=commandRegIsUnsupported|commandRegBadHaltResume ;  
   wire goAbstract=(|ctrlStateReg)&_GEN_2&~_GEN_3 ;  
   wire _GEN_4=ctrlStateReg==2'h2 ;  
   wire _GEN_5=(|ctrlStateReg)&~_GEN_2 ;  
  always @( posedge clock)
       begin 
         if (io_dmactive&~goAbstract&hartGoingWrEn&~reset&(|(auto_tl_in_a_bits_data[41:32])))
            begin 
              if (1)$display("Assertion failed: Unexpected 'GOING' hart.\n    at Debug.scala:1499 assert(hartGoingId === 0.U, \"Unexpected 'GOING' hart.\")//Chisel3 #540 %%%%x, expected %%%%x\", hartGoingId, 0.U)\n");
              if (1)$display("");
            end 
         if (_GEN_5&_GEN_4&hartExceptionWrEn&~reset&(|(auto_tl_in_a_bits_data[41:32])))
            begin 
              if (1)$display("Assertion failed: Unexpected 'EXCEPTION' hart\n    at Debug.scala:1820 assert(hartExceptionId === 0.U, \"Unexpected 'EXCEPTION' hart\")//Chisel3 #540, %%%%x, expected %%%%x\", hartExceptionId, 0.U)\n");
              if (1)$display("");
            end 
         if (_GEN_5&~_GEN_4&(&ctrlStateReg)&~reset)
            begin 
              if (1)$display("Assertion failed: Should not be in custom state unless we need it.\n    at Debug.scala:1825 assert(needCustom.B, \"Should not be in custom state unless we need it.\")\n");
              if (1)$display("");
            end 
         if (~reset&~(~io_dmactive|~hartExceptionWrEn|_GEN_4))
            begin 
              if (1)$display("Assertion failed: Unexpected EXCEPTION write: should only get it in Debug Module EXEC state\n    at Debug.scala:1838 assert ((!io.dmactive || !hartExceptionWrEn || ctrlStateReg === CtrlState(Exec)),\n");
              if (1)$display("");
            end 
       end
  
   wire dmiAbstractDataAccessVec_0=dmiAbstractDataWrEnMaybe_0|out_roready_27&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiAbstractDataAccessVec_4=dmiAbstractDataWrEnMaybe_4|out_roready_3&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_0=dmiProgramBufferWrEnMaybe_0|out_roready_78&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_4=dmiProgramBufferWrEnMaybe_4|out_roready_50&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_8=dmiProgramBufferWrEnMaybe_8|out_roready_82&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_12=dmiProgramBufferWrEnMaybe_12|out_roready_19&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_16=dmiProgramBufferWrEnMaybe_16|out_roready_99&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_20=dmiProgramBufferWrEnMaybe_20|out_roready_42&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_24=dmiProgramBufferWrEnMaybe_24|out_roready_46&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_28=dmiProgramBufferWrEnMaybe_28|out_roready_15&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_32=dmiProgramBufferWrEnMaybe_32|out_roready_97&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_36=dmiProgramBufferWrEnMaybe_36|out_roready_9&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_40=dmiProgramBufferWrEnMaybe_40|out_roready_35&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_44=dmiProgramBufferWrEnMaybe_44|out_roready_23&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_48=dmiProgramBufferWrEnMaybe_48|out_roready_93&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_52=dmiProgramBufferWrEnMaybe_52|out_roready_54&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_56=dmiProgramBufferWrEnMaybe_56|out_roready_7&auto_dmi_in_a_bits_mask[0] ;  
   wire dmiProgramBufferAccessVec_60=dmiProgramBufferWrEnMaybe_60|out_roready_31&auto_dmi_in_a_bits_mask[0] ;  
   wire autoexec=dmiAbstractDataAccessVec_0&ABSTRACTAUTOReg_autoexecdata[0]|dmiAbstractDataAccessVec_4&ABSTRACTAUTOReg_autoexecdata[1]|dmiProgramBufferAccessVec_0&ABSTRACTAUTOReg_autoexecprogbuf[0]|dmiProgramBufferAccessVec_4&ABSTRACTAUTOReg_autoexecprogbuf[1]|dmiProgramBufferAccessVec_8&ABSTRACTAUTOReg_autoexecprogbuf[2]|dmiProgramBufferAccessVec_12&ABSTRACTAUTOReg_autoexecprogbuf[3]|dmiProgramBufferAccessVec_16&ABSTRACTAUTOReg_autoexecprogbuf[4]|dmiProgramBufferAccessVec_20&ABSTRACTAUTOReg_autoexecprogbuf[5]|dmiProgramBufferAccessVec_24&ABSTRACTAUTOReg_autoexecprogbuf[6]|dmiProgramBufferAccessVec_28&ABSTRACTAUTOReg_autoexecprogbuf[7]|dmiProgramBufferAccessVec_32&ABSTRACTAUTOReg_autoexecprogbuf[8]|dmiProgramBufferAccessVec_36&ABSTRACTAUTOReg_autoexecprogbuf[9]|dmiProgramBufferAccessVec_40&ABSTRACTAUTOReg_autoexecprogbuf[10]|dmiProgramBufferAccessVec_44&ABSTRACTAUTOReg_autoexecprogbuf[11]|dmiProgramBufferAccessVec_48&ABSTRACTAUTOReg_autoexecprogbuf[12]|dmiProgramBufferAccessVec_52&ABSTRACTAUTOReg_autoexecprogbuf[13]|dmiProgramBufferAccessVec_56&ABSTRACTAUTOReg_autoexecprogbuf[14]|dmiProgramBufferAccessVec_60&ABSTRACTAUTOReg_autoexecprogbuf[15] ;  
   wire COMMANDWrEn=COMMANDWrEnMaybe&~(|ctrlStateReg) ;  
   wire _regAccessRegisterCommand_T_1=ABSTRACTCSReg_cmderr==3'h0 ;  
   wire _GEN_6=COMMANDWrEn&~(|(COMMANDWrDataVal[31:24]))&_regAccessRegisterCommand_T_1|autoexec&commandRegIsAccessRegister&_regAccessRegisterCommand_T_1 ;  
  always @( posedge clock)
       begin 
         haltedBitRegs <=io_dmactive&(hartHaltedWrEn|~hartResumingWrEn&haltedBitRegs)&~_hartIsInResetSync_0_debug_hartReset_0_io_q;
         resumeReqRegs <=io_dmactive&(resumereq ? (resumeReqRegs|hamaskWrSel_0)&~_hartIsInResetSync_0_debug_hartReset_0_io_q:~hartResumingWrEn&resumeReqRegs&~_hartIsInResetSync_0_debug_hartReset_0_io_q);
         haveResetBitRegs <=io_dmactive&(io_innerCtrl_valid&io_innerCtrl_bits_ackhavereset ? haveResetBitRegs&~hamaskWrSel_0|_hartIsInResetSync_0_debug_hartReset_0_io_q:haveResetBitRegs|_hartIsInResetSync_0_debug_hartReset_0_io_q);
         if (io_dmactive)
            begin 
              if (ABSTRACTCSWrEnMaybe&(|ctrlStateReg)|autoexecdataWrEnMaybe&(|ctrlStateReg)|autoexecprogbufWrEnMaybe&(|ctrlStateReg)|COMMANDWrEnMaybe&(|ctrlStateReg)|(dmiAbstractDataAccessVec_0|dmiAbstractDataWrEnMaybe_1|out_roready_27&auto_dmi_in_a_bits_mask[1]|dmiAbstractDataWrEnMaybe_2|out_roready_27&auto_dmi_in_a_bits_mask[2]|dmiAbstractDataWrEnMaybe_3|out_roready_27&auto_dmi_in_a_bits_mask[3]|dmiAbstractDataAccessVec_4|dmiAbstractDataWrEnMaybe_5|out_roready_3&auto_dmi_in_a_bits_mask[1]|dmiAbstractDataWrEnMaybe_6|out_roready_3&auto_dmi_in_a_bits_mask[2]|dmiAbstractDataWrEnMaybe_7|out_roready_3&auto_dmi_in_a_bits_mask[3])&(|ctrlStateReg)|(dmiProgramBufferAccessVec_0|dmiProgramBufferWrEnMaybe_1|out_roready_78&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_2|out_roready_78&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_3|out_roready_78&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_4|dmiProgramBufferWrEnMaybe_5|out_roready_50&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_6|out_roready_50&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_7|out_roready_50&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_8|dmiProgramBufferWrEnMaybe_9|out_roready_82&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_10|out_roready_82&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_11|out_roready_82&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_12|dmiProgramBufferWrEnMaybe_13|out_roready_19&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_14|out_roready_19&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_15|out_roready_19&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_16|dmiProgramBufferWrEnMaybe_17|out_roready_99&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_18|out_roready_99&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_19|out_roready_99&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_20|dmiProgramBufferWrEnMaybe_21|out_roready_42&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_22|out_roready_42&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_23|out_roready_42&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_24|dmiProgramBufferWrEnMaybe_25|out_roready_46&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_26|out_roready_46&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_27|out_roready_46&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_28|dmiProgramBufferWrEnMaybe_29|out_roready_15&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_30|out_roready_15&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_31|out_roready_15&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_32|dmiProgramBufferWrEnMaybe_33|out_roready_97&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_34|out_roready_97&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_35|out_roready_97&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_36|dmiProgramBufferWrEnMaybe_37|out_roready_9&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_38|out_roready_9&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_39|out_roready_9&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_40|dmiProgramBufferWrEnMaybe_41|out_roready_35&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_42|out_roready_35&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_43|out_roready_35&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_44|dmiProgramBufferWrEnMaybe_45|out_roready_23&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_46|out_roready_23&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_47|out_roready_23&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_48|dmiProgramBufferWrEnMaybe_49|out_roready_93&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_50|out_roready_93&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_51|out_roready_93&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_52|dmiProgramBufferWrEnMaybe_53|out_roready_54&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_54|out_roready_54&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_55|out_roready_54&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_56|dmiProgramBufferWrEnMaybe_57|out_roready_7&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_58|out_roready_7&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_59|out_roready_7&auto_dmi_in_a_bits_mask[3]|dmiProgramBufferAccessVec_60|dmiProgramBufferWrEnMaybe_61|out_roready_31&auto_dmi_in_a_bits_mask[1]|dmiProgramBufferWrEnMaybe_62|out_roready_31&auto_dmi_in_a_bits_mask[2]|dmiProgramBufferWrEnMaybe_63|out_roready_31&auto_dmi_in_a_bits_mask[3])&(|ctrlStateReg))
                 ABSTRACTCSReg_cmderr <=3'h1;
               else 
                 if (~(~(|ctrlStateReg)|_GEN_2)&_GEN_4&hartExceptionWrEn)
                    ABSTRACTCSReg_cmderr <=3'h3;
                  else 
                    if ((|ctrlStateReg) ? _GEN_2&commandRegIsUnsupported:~_GEN_6&(COMMANDWrEn&(|(COMMANDWrDataVal[31:24]))|autoexec&commandRegIsUnsupported))
                       ABSTRACTCSReg_cmderr <=3'h2;
                     else 
                       if ((|ctrlStateReg)&_GEN_2&~commandRegIsUnsupported&commandRegBadHaltResume)
                          ABSTRACTCSReg_cmderr <=3'h4;
                        else 
                          ABSTRACTCSReg_cmderr <=({3{~(ABSTRACTCSWrEnMaybe&~(|ctrlStateReg))}}|~(auto_dmi_in_a_bits_data[10:8]))&ABSTRACTCSReg_cmderr;
              if (autoexecprogbufWrEnMaybe&~(|ctrlStateReg))
                 ABSTRACTAUTOReg_autoexecprogbuf <=auto_dmi_in_a_bits_data[31:16];
              if (autoexecdataWrEnMaybe&~(|ctrlStateReg))
                 ABSTRACTAUTOReg_autoexecdata <={10'h0,auto_dmi_in_a_bits_data[1:0]};
              if (COMMANDWrEn)
                 begin 
                   COMMANDReg_cmdtype <=COMMANDWrDataVal[31:24];
                   COMMANDReg_control <=COMMANDWrDataVal[23:0];
                 end 
              if (out_woready_1_818&auto_tl_in_a_bits_mask[0])
                 abstractDataMem_0 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiAbstractDataWrEnMaybe_0&~(|ctrlStateReg))
                    abstractDataMem_0 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_818&auto_tl_in_a_bits_mask[1])
                 abstractDataMem_1 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiAbstractDataWrEnMaybe_1&~(|ctrlStateReg))
                    abstractDataMem_1 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_818&auto_tl_in_a_bits_mask[2])
                 abstractDataMem_2 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiAbstractDataWrEnMaybe_2&~(|ctrlStateReg))
                    abstractDataMem_2 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_818&auto_tl_in_a_bits_mask[3])
                 abstractDataMem_3 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiAbstractDataWrEnMaybe_3&~(|ctrlStateReg))
                    abstractDataMem_3 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_818&auto_tl_in_a_bits_mask[4])
                 abstractDataMem_4 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiAbstractDataWrEnMaybe_4&~(|ctrlStateReg))
                    abstractDataMem_4 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_818&auto_tl_in_a_bits_mask[5])
                 abstractDataMem_5 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiAbstractDataWrEnMaybe_5&~(|ctrlStateReg))
                    abstractDataMem_5 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_818&auto_tl_in_a_bits_mask[6])
                 abstractDataMem_6 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiAbstractDataWrEnMaybe_6&~(|ctrlStateReg))
                    abstractDataMem_6 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_818&auto_tl_in_a_bits_mask[7])
                 abstractDataMem_7 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiAbstractDataWrEnMaybe_7&~(|ctrlStateReg))
                    abstractDataMem_7 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[0])
                 programBufferMem_0 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_0&~(|ctrlStateReg))
                    programBufferMem_0 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[1])
                 programBufferMem_1 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_1&~(|ctrlStateReg))
                    programBufferMem_1 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[2])
                 programBufferMem_2 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_2&~(|ctrlStateReg))
                    programBufferMem_2 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[3])
                 programBufferMem_3 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_3&~(|ctrlStateReg))
                    programBufferMem_3 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[4])
                 programBufferMem_4 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_4&~(|ctrlStateReg))
                    programBufferMem_4 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[5])
                 programBufferMem_5 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_5&~(|ctrlStateReg))
                    programBufferMem_5 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[6])
                 programBufferMem_6 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_6&~(|ctrlStateReg))
                    programBufferMem_6 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_922&auto_tl_in_a_bits_mask[7])
                 programBufferMem_7 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_7&~(|ctrlStateReg))
                    programBufferMem_7 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[0])
                 programBufferMem_8 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_8&~(|ctrlStateReg))
                    programBufferMem_8 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[1])
                 programBufferMem_9 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_9&~(|ctrlStateReg))
                    programBufferMem_9 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[2])
                 programBufferMem_10 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_10&~(|ctrlStateReg))
                    programBufferMem_10 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[3])
                 programBufferMem_11 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_11&~(|ctrlStateReg))
                    programBufferMem_11 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[4])
                 programBufferMem_12 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_12&~(|ctrlStateReg))
                    programBufferMem_12 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[5])
                 programBufferMem_13 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_13&~(|ctrlStateReg))
                    programBufferMem_13 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[6])
                 programBufferMem_14 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_14&~(|ctrlStateReg))
                    programBufferMem_14 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_510&auto_tl_in_a_bits_mask[7])
                 programBufferMem_15 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_15&~(|ctrlStateReg))
                    programBufferMem_15 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[0])
                 programBufferMem_16 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_16&~(|ctrlStateReg))
                    programBufferMem_16 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[1])
                 programBufferMem_17 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_17&~(|ctrlStateReg))
                    programBufferMem_17 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[2])
                 programBufferMem_18 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_18&~(|ctrlStateReg))
                    programBufferMem_18 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[3])
                 programBufferMem_19 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_19&~(|ctrlStateReg))
                    programBufferMem_19 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[4])
                 programBufferMem_20 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_20&~(|ctrlStateReg))
                    programBufferMem_20 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[5])
                 programBufferMem_21 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_21&~(|ctrlStateReg))
                    programBufferMem_21 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[6])
                 programBufferMem_22 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_22&~(|ctrlStateReg))
                    programBufferMem_22 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_191&auto_tl_in_a_bits_mask[7])
                 programBufferMem_23 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_23&~(|ctrlStateReg))
                    programBufferMem_23 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[0])
                 programBufferMem_24 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_24&~(|ctrlStateReg))
                    programBufferMem_24 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[1])
                 programBufferMem_25 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_25&~(|ctrlStateReg))
                    programBufferMem_25 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[2])
                 programBufferMem_26 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_26&~(|ctrlStateReg))
                    programBufferMem_26 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[3])
                 programBufferMem_27 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_27&~(|ctrlStateReg))
                    programBufferMem_27 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[4])
                 programBufferMem_28 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_28&~(|ctrlStateReg))
                    programBufferMem_28 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[5])
                 programBufferMem_29 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_29&~(|ctrlStateReg))
                    programBufferMem_29 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[6])
                 programBufferMem_30 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_30&~(|ctrlStateReg))
                    programBufferMem_30 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_1074&auto_tl_in_a_bits_mask[7])
                 programBufferMem_31 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_31&~(|ctrlStateReg))
                    programBufferMem_31 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[0])
                 programBufferMem_32 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_32&~(|ctrlStateReg))
                    programBufferMem_32 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[1])
                 programBufferMem_33 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_33&~(|ctrlStateReg))
                    programBufferMem_33 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[2])
                 programBufferMem_34 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_34&~(|ctrlStateReg))
                    programBufferMem_34 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[3])
                 programBufferMem_35 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_35&~(|ctrlStateReg))
                    programBufferMem_35 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[4])
                 programBufferMem_36 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_36&~(|ctrlStateReg))
                    programBufferMem_36 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[5])
                 programBufferMem_37 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_37&~(|ctrlStateReg))
                    programBufferMem_37 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[6])
                 programBufferMem_38 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_38&~(|ctrlStateReg))
                    programBufferMem_38 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_722&auto_tl_in_a_bits_mask[7])
                 programBufferMem_39 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_39&~(|ctrlStateReg))
                    programBufferMem_39 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[0])
                 programBufferMem_40 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_40&~(|ctrlStateReg))
                    programBufferMem_40 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[1])
                 programBufferMem_41 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_41&~(|ctrlStateReg))
                    programBufferMem_41 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[2])
                 programBufferMem_42 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_42&~(|ctrlStateReg))
                    programBufferMem_42 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[3])
                 programBufferMem_43 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_43&~(|ctrlStateReg))
                    programBufferMem_43 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[4])
                 programBufferMem_44 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_44&~(|ctrlStateReg))
                    programBufferMem_44 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[5])
                 programBufferMem_45 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_45&~(|ctrlStateReg))
                    programBufferMem_45 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[6])
                 programBufferMem_46 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_46&~(|ctrlStateReg))
                    programBufferMem_46 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_442&auto_tl_in_a_bits_mask[7])
                 programBufferMem_47 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_47&~(|ctrlStateReg))
                    programBufferMem_47 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[0])
                 programBufferMem_48 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_48&~(|ctrlStateReg))
                    programBufferMem_48 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[1])
                 programBufferMem_49 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_49&~(|ctrlStateReg))
                    programBufferMem_49 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[2])
                 programBufferMem_50 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_50&~(|ctrlStateReg))
                    programBufferMem_50 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[3])
                 programBufferMem_51 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_51&~(|ctrlStateReg))
                    programBufferMem_51 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[4])
                 programBufferMem_52 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_52&~(|ctrlStateReg))
                    programBufferMem_52 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[5])
                 programBufferMem_53 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_53&~(|ctrlStateReg))
                    programBufferMem_53 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[6])
                 programBufferMem_54 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_54&~(|ctrlStateReg))
                    programBufferMem_54 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_111&auto_tl_in_a_bits_mask[7])
                 programBufferMem_55 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_55&~(|ctrlStateReg))
                    programBufferMem_55 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[0])
                 programBufferMem_56 <=auto_tl_in_a_bits_data[7:0];
               else 
                 if (dmiProgramBufferWrEnMaybe_56&~(|ctrlStateReg))
                    programBufferMem_56 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[1])
                 programBufferMem_57 <=auto_tl_in_a_bits_data[15:8];
               else 
                 if (dmiProgramBufferWrEnMaybe_57&~(|ctrlStateReg))
                    programBufferMem_57 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[2])
                 programBufferMem_58 <=auto_tl_in_a_bits_data[23:16];
               else 
                 if (dmiProgramBufferWrEnMaybe_58&~(|ctrlStateReg))
                    programBufferMem_58 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[3])
                 programBufferMem_59 <=auto_tl_in_a_bits_data[31:24];
               else 
                 if (dmiProgramBufferWrEnMaybe_59&~(|ctrlStateReg))
                    programBufferMem_59 <=auto_dmi_in_a_bits_data[31:24];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[4])
                 programBufferMem_60 <=auto_tl_in_a_bits_data[39:32];
               else 
                 if (dmiProgramBufferWrEnMaybe_60&~(|ctrlStateReg))
                    programBufferMem_60 <=auto_dmi_in_a_bits_data[7:0];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[5])
                 programBufferMem_61 <=auto_tl_in_a_bits_data[47:40];
               else 
                 if (dmiProgramBufferWrEnMaybe_61&~(|ctrlStateReg))
                    programBufferMem_61 <=auto_dmi_in_a_bits_data[15:8];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[6])
                 programBufferMem_62 <=auto_tl_in_a_bits_data[55:48];
               else 
                 if (dmiProgramBufferWrEnMaybe_62&~(|ctrlStateReg))
                    programBufferMem_62 <=auto_dmi_in_a_bits_data[23:16];
              if (out_woready_1_1146&auto_tl_in_a_bits_mask[7])
                 programBufferMem_63 <=auto_tl_in_a_bits_data[63:56];
               else 
                 if (dmiProgramBufferWrEnMaybe_63&~(|ctrlStateReg))
                    programBufferMem_63 <=auto_dmi_in_a_bits_data[31:24];
              if (|ctrlStateReg)
                 begin 
                   if (_GEN_2)
                      ctrlStateReg <={~_GEN_3,1'h0};
                    else 
                      if (_GEN_4&(hartExceptionWrEn|~goReg&hartHaltedWrEn))
                         ctrlStateReg <=2'h0;
                 end 
               else 
                 if (_GEN_6)
                    ctrlStateReg <=2'h1;
            end 
          else 
            begin 
              ABSTRACTCSReg_cmderr <=3'h0;
              ABSTRACTAUTOReg_autoexecprogbuf <=16'h0;
              ABSTRACTAUTOReg_autoexecdata <=12'h0;
              COMMANDReg_cmdtype <=8'h0;
              COMMANDReg_control <=24'h0;
              abstractDataMem_0 <=8'h0;
              abstractDataMem_1 <=8'h0;
              abstractDataMem_2 <=8'h0;
              abstractDataMem_3 <=8'h0;
              abstractDataMem_4 <=8'h0;
              abstractDataMem_5 <=8'h0;
              abstractDataMem_6 <=8'h0;
              abstractDataMem_7 <=8'h0;
              programBufferMem_0 <=8'h0;
              programBufferMem_1 <=8'h0;
              programBufferMem_2 <=8'h0;
              programBufferMem_3 <=8'h0;
              programBufferMem_4 <=8'h0;
              programBufferMem_5 <=8'h0;
              programBufferMem_6 <=8'h0;
              programBufferMem_7 <=8'h0;
              programBufferMem_8 <=8'h0;
              programBufferMem_9 <=8'h0;
              programBufferMem_10 <=8'h0;
              programBufferMem_11 <=8'h0;
              programBufferMem_12 <=8'h0;
              programBufferMem_13 <=8'h0;
              programBufferMem_14 <=8'h0;
              programBufferMem_15 <=8'h0;
              programBufferMem_16 <=8'h0;
              programBufferMem_17 <=8'h0;
              programBufferMem_18 <=8'h0;
              programBufferMem_19 <=8'h0;
              programBufferMem_20 <=8'h0;
              programBufferMem_21 <=8'h0;
              programBufferMem_22 <=8'h0;
              programBufferMem_23 <=8'h0;
              programBufferMem_24 <=8'h0;
              programBufferMem_25 <=8'h0;
              programBufferMem_26 <=8'h0;
              programBufferMem_27 <=8'h0;
              programBufferMem_28 <=8'h0;
              programBufferMem_29 <=8'h0;
              programBufferMem_30 <=8'h0;
              programBufferMem_31 <=8'h0;
              programBufferMem_32 <=8'h0;
              programBufferMem_33 <=8'h0;
              programBufferMem_34 <=8'h0;
              programBufferMem_35 <=8'h0;
              programBufferMem_36 <=8'h0;
              programBufferMem_37 <=8'h0;
              programBufferMem_38 <=8'h0;
              programBufferMem_39 <=8'h0;
              programBufferMem_40 <=8'h0;
              programBufferMem_41 <=8'h0;
              programBufferMem_42 <=8'h0;
              programBufferMem_43 <=8'h0;
              programBufferMem_44 <=8'h0;
              programBufferMem_45 <=8'h0;
              programBufferMem_46 <=8'h0;
              programBufferMem_47 <=8'h0;
              programBufferMem_48 <=8'h0;
              programBufferMem_49 <=8'h0;
              programBufferMem_50 <=8'h0;
              programBufferMem_51 <=8'h0;
              programBufferMem_52 <=8'h0;
              programBufferMem_53 <=8'h0;
              programBufferMem_54 <=8'h0;
              programBufferMem_55 <=8'h0;
              programBufferMem_56 <=8'h0;
              programBufferMem_57 <=8'h0;
              programBufferMem_58 <=8'h0;
              programBufferMem_59 <=8'h0;
              programBufferMem_60 <=8'h0;
              programBufferMem_61 <=8'h0;
              programBufferMem_62 <=8'h0;
              programBufferMem_63 <=8'h0;
              ctrlStateReg <=2'h0;
            end 
         goReg <=io_dmactive&(goAbstract|~hartGoingWrEn&goReg);
         if (goAbstract)
            begin 
              abstractGeneratedMem_0 <=COMMANDReg_control[17] ? (COMMANDReg_control[16] ? {17'h7000,COMMANDReg_control[22:20],COMMANDReg_control[4:0],7'h3}:{7'h1C,COMMANDReg_control[4:0],5'h0,COMMANDReg_control[22:20],12'h23}):32'h13;
              abstractGeneratedMem_1 <=COMMANDReg_control[18] ? 32'h13:32'h100073;
            end 
         if (reset)
            hrmaskReg_0 <=1'h0;
          else 
            hrmaskReg_0 <=io_dmactive&(io_innerCtrl_valid ? io_innerCtrl_bits_hrmask_0:hrmaskReg_0);
       end
  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            hrDebugIntReg_0 <=1'h0;
          else 
            hrDebugIntReg_0 <=io_dmactive&hrmaskReg_0&(_hartIsInResetSync_0_debug_hartReset_0_io_q|hrDebugIntReg_0&~haltedBitRegs);
       end
  
  TLMonitor_33 monitor(.clock(clock),.reset(reset),.io_in_a_ready(auto_dmi_in_d_ready),.io_in_a_valid(auto_dmi_in_a_valid),.io_in_a_bits_opcode(auto_dmi_in_a_bits_opcode),.io_in_a_bits_param(auto_dmi_in_a_bits_param),.io_in_a_bits_size(auto_dmi_in_a_bits_size),.io_in_a_bits_source(auto_dmi_in_a_bits_source),.io_in_a_bits_address(auto_dmi_in_a_bits_address),.io_in_a_bits_mask(auto_dmi_in_a_bits_mask),.io_in_a_bits_corrupt(auto_dmi_in_a_bits_corrupt),.io_in_d_ready(auto_dmi_in_d_ready),.io_in_d_valid(auto_dmi_in_a_valid),.io_in_d_bits_opcode(dmiNodeIn_d_bits_opcode),.io_in_d_bits_size(auto_dmi_in_a_bits_size),.io_in_d_bits_source(auto_dmi_in_a_bits_source)); 
  TLMonitor_34 monitor_1(.clock(clock),.reset(reset),.io_in_a_ready(auto_tl_in_d_ready),.io_in_a_valid(auto_tl_in_a_valid),.io_in_a_bits_opcode(auto_tl_in_a_bits_opcode),.io_in_a_bits_param(auto_tl_in_a_bits_param),.io_in_a_bits_size(auto_tl_in_a_bits_size),.io_in_a_bits_source(auto_tl_in_a_bits_source),.io_in_a_bits_address(auto_tl_in_a_bits_address),.io_in_a_bits_mask(auto_tl_in_a_bits_mask),.io_in_a_bits_corrupt(auto_tl_in_a_bits_corrupt),.io_in_d_ready(auto_tl_in_d_ready),.io_in_d_valid(auto_tl_in_a_valid),.io_in_d_bits_opcode(tlNodeIn_d_bits_opcode),.io_in_d_bits_size(auto_tl_in_a_bits_size),.io_in_d_bits_source(auto_tl_in_a_bits_source)); 
  AsyncResetSynchronizerShiftReg_w1_d3_i0 hartIsInResetSync_0_debug_hartReset_0(.clock(clock),.reset(reset),.io_d(io_hartIsInReset_0),.io_q(_hartIsInResetSync_0_debug_hartReset_0_io_q)); 
  assign auto_tl_in_a_ready=auto_tl_in_d_ready; 
  assign auto_tl_in_d_valid=auto_tl_in_a_valid; 
  assign auto_tl_in_d_bits_opcode=tlNodeIn_d_bits_opcode; 
  assign auto_tl_in_d_bits_size=auto_tl_in_a_bits_size; 
  assign auto_tl_in_d_bits_source=auto_tl_in_a_bits_source; 
  assign auto_tl_in_d_bits_data=casez_tmp_1 ? casez_tmp_2:64'h0; 
  assign auto_dmi_in_a_ready=auto_dmi_in_d_ready; 
  assign auto_dmi_in_d_valid=auto_dmi_in_a_valid; 
  assign auto_dmi_in_d_bits_opcode=dmiNodeIn_d_bits_opcode; 
  assign auto_dmi_in_d_bits_size=auto_dmi_in_a_bits_size; 
  assign auto_dmi_in_d_bits_source=auto_dmi_in_a_bits_source; 
  assign auto_dmi_in_d_bits_data=casez_tmp ? casez_tmp_0:32'h0; 
  assign io_hgDebugInt_0=hrDebugIntReg_0; 
endmodule
 
module ClockCrossingReg_w55 (
  input clock,
  input [54:0] io_d,
  output [54:0] io_q,
  input io_en) ; 
   reg [54:0] cdc_reg ;  
  always @( posedge clock)
       begin 
         if (io_en)
            cdc_reg <=io_d;
       end
  
  assign io_q=cdc_reg; 
endmodule
 
module AsyncQueueSink_1 (
  input clock,
  input reset,
  input io_deq_ready,
  output io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [2:0] io_deq_bits_param,
  output [1:0] io_deq_bits_size,
  output io_deq_bits_source,
  output [8:0] io_deq_bits_address,
  output [3:0] io_deq_bits_mask,
  output [31:0] io_deq_bits_data,
  output io_deq_bits_corrupt,
  input [2:0] io_async_mem_0_opcode,
  input [8:0] io_async_mem_0_address,
  input [31:0] io_async_mem_0_data,
  output io_async_ridx,
  input io_async_widx,
  output io_async_safe_ridx_valid,
  input io_async_safe_widx_valid,
  input io_async_safe_source_reset_n,
  output io_async_safe_sink_reset_n) ; 
   wire io_deq_valid_0 ;  
   wire _source_valid_io_out ;  
   wire _source_extend_io_out ;  
   wire _sink_valid_0_io_out ;  
   wire [54:0] _io_deq_bits_deq_bits_reg_io_q ;  
   wire _widx_widx_gray_io_q ;  
   reg ridx_ridx_bin ;  
   wire ridx=_source_valid_io_out&ridx_ridx_bin+(io_deq_ready&io_deq_valid_0) ;  
   wire valid=_source_valid_io_out&ridx!=_widx_widx_gray_io_q ;  
   reg valid_reg ;  
  assign io_deq_valid_0=valid_reg&_source_valid_io_out; 
   reg ridx_gray ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              ridx_ridx_bin <=1'h0;
              valid_reg <=1'h0;
              ridx_gray <=1'h0;
            end 
          else 
            begin 
              ridx_ridx_bin <=ridx;
              valid_reg <=valid;
              ridx_gray <=ridx;
            end 
       end
  
  AsyncResetSynchronizerShiftReg_w1_d3_i0 widx_widx_gray(.clock(clock),.reset(reset),.io_d(io_async_widx),.io_q(_widx_widx_gray_io_q)); 
  ClockCrossingReg_w55 io_deq_bits_deq_bits_reg(.clock(clock),.io_d({io_async_mem_0_opcode,6'h4,io_async_mem_0_address,4'hF,io_async_mem_0_data,1'h0}),.io_q(_io_deq_bits_deq_bits_reg_io_q),.io_en(valid)); 
  AsyncValidSync sink_valid_0(.io_in(1'h1),.io_out(_sink_valid_0_io_out),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync sink_valid_1(.io_in(_sink_valid_0_io_out),.io_out(io_async_safe_ridx_valid),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync source_extend(.io_in(io_async_safe_widx_valid),.io_out(_source_extend_io_out),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync source_valid(.io_in(_source_extend_io_out),.io_out(_source_valid_io_out),.clock(clock),.reset(reset)); 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_opcode=_io_deq_bits_deq_bits_reg_io_q[54:52]; 
  assign io_deq_bits_param=_io_deq_bits_deq_bits_reg_io_q[51:49]; 
  assign io_deq_bits_size=_io_deq_bits_deq_bits_reg_io_q[48:47]; 
  assign io_deq_bits_source=_io_deq_bits_deq_bits_reg_io_q[46]; 
  assign io_deq_bits_address=_io_deq_bits_deq_bits_reg_io_q[45:37]; 
  assign io_deq_bits_mask=_io_deq_bits_deq_bits_reg_io_q[36:33]; 
  assign io_deq_bits_data=_io_deq_bits_deq_bits_reg_io_q[32:1]; 
  assign io_deq_bits_corrupt=_io_deq_bits_deq_bits_reg_io_q[0]; 
  assign io_async_ridx=ridx_gray; 
  assign io_async_safe_sink_reset_n=~reset; 
endmodule
 
module AsyncQueueSource_2 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [2:0] io_enq_bits_opcode,
  input [1:0] io_enq_bits_size,
  input io_enq_bits_source,
  input [31:0] io_enq_bits_data,
  output [2:0] io_async_mem_0_opcode,
  output [1:0] io_async_mem_0_size,
  output io_async_mem_0_source,
  output [31:0] io_async_mem_0_data,
  input io_async_ridx,
  output io_async_widx,
  input io_async_safe_ridx_valid,
  output io_async_safe_widx_valid,
  output io_async_safe_source_reset_n,
  input io_async_safe_sink_reset_n) ; 
   wire io_enq_ready_0 ;  
   wire _sink_valid_io_out ;  
   wire _sink_extend_io_out ;  
   wire _source_valid_0_io_out ;  
   wire _ridx_ridx_gray_io_q ;  
   reg [2:0] mem_0_opcode ;  
   reg [1:0] mem_0_size ;  
   reg mem_0_source ;  
   reg [31:0] mem_0_data ;  
   wire _widx_T_1=io_enq_ready_0&io_enq_valid ;  
   reg widx_widx_bin ;  
   reg ready_reg ;  
  assign io_enq_ready_0=ready_reg&_sink_valid_io_out; 
   reg widx_gray ;  
  always @( posedge clock)
       begin 
         if (_widx_T_1)
            begin 
              mem_0_opcode <=io_enq_bits_opcode;
              mem_0_size <=io_enq_bits_size;
              mem_0_source <=io_enq_bits_source;
              mem_0_data <=io_enq_bits_data;
            end 
       end
  
   wire widx=_sink_valid_io_out&widx_widx_bin+_widx_T_1 ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              widx_widx_bin <=1'h0;
              ready_reg <=1'h0;
              widx_gray <=1'h0;
            end 
          else 
            begin 
              widx_widx_bin <=widx;
              ready_reg <=_sink_valid_io_out&widx!=~_ridx_ridx_gray_io_q;
              widx_gray <=widx;
            end 
       end
  
  AsyncResetSynchronizerShiftReg_w1_d3_i0 ridx_ridx_gray(.clock(clock),.reset(reset),.io_d(io_async_ridx),.io_q(_ridx_ridx_gray_io_q)); 
  AsyncValidSync source_valid_0(.io_in(1'h1),.io_out(_source_valid_0_io_out),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync source_valid_1(.io_in(_source_valid_0_io_out),.io_out(io_async_safe_widx_valid),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync sink_extend(.io_in(io_async_safe_ridx_valid),.io_out(_sink_extend_io_out),.clock(clock),.reset(reset|~io_async_safe_sink_reset_n)); 
  AsyncValidSync sink_valid(.io_in(_sink_extend_io_out),.io_out(_sink_valid_io_out),.clock(clock),.reset(reset)); 
  assign io_enq_ready=io_enq_ready_0; 
  assign io_async_mem_0_opcode=mem_0_opcode; 
  assign io_async_mem_0_size=mem_0_size; 
  assign io_async_mem_0_source=mem_0_source; 
  assign io_async_mem_0_data=mem_0_data; 
  assign io_async_widx=widx_gray; 
  assign io_async_safe_source_reset_n=~reset; 
endmodule
 
module TLAsyncCrossingSink (
  input clock,
  input reset,
  input [2:0] auto_in_a_mem_0_opcode,
  input [8:0] auto_in_a_mem_0_address,
  input [31:0] auto_in_a_mem_0_data,
  output auto_in_a_ridx,
  input auto_in_a_widx,
  output auto_in_a_safe_ridx_valid,
  input auto_in_a_safe_widx_valid,
  input auto_in_a_safe_source_reset_n,
  output auto_in_a_safe_sink_reset_n,
  output [2:0] auto_in_d_mem_0_opcode,
  output [1:0] auto_in_d_mem_0_size,
  output auto_in_d_mem_0_source,
  output [31:0] auto_in_d_mem_0_data,
  input auto_in_d_ridx,
  output auto_in_d_widx,
  input auto_in_d_safe_ridx_valid,
  output auto_in_d_safe_widx_valid,
  output auto_in_d_safe_source_reset_n,
  input auto_in_d_safe_sink_reset_n,
  input auto_out_a_ready,
  output auto_out_a_valid,
  output [2:0] auto_out_a_bits_opcode,
  output [2:0] auto_out_a_bits_param,
  output [1:0] auto_out_a_bits_size,
  output auto_out_a_bits_source,
  output [8:0] auto_out_a_bits_address,
  output [3:0] auto_out_a_bits_mask,
  output [31:0] auto_out_a_bits_data,
  output auto_out_a_bits_corrupt,
  output auto_out_d_ready,
  input auto_out_d_valid,
  input [2:0] auto_out_d_bits_opcode,
  input [1:0] auto_out_d_bits_size,
  input auto_out_d_bits_source,
  input [31:0] auto_out_d_bits_data) ; 
  AsyncQueueSink_1 nodeOut_a_sink(.clock(clock),.reset(reset),.io_deq_ready(auto_out_a_ready),.io_deq_valid(auto_out_a_valid),.io_deq_bits_opcode(auto_out_a_bits_opcode),.io_deq_bits_param(auto_out_a_bits_param),.io_deq_bits_size(auto_out_a_bits_size),.io_deq_bits_source(auto_out_a_bits_source),.io_deq_bits_address(auto_out_a_bits_address),.io_deq_bits_mask(auto_out_a_bits_mask),.io_deq_bits_data(auto_out_a_bits_data),.io_deq_bits_corrupt(auto_out_a_bits_corrupt),.io_async_mem_0_opcode(auto_in_a_mem_0_opcode),.io_async_mem_0_address(auto_in_a_mem_0_address),.io_async_mem_0_data(auto_in_a_mem_0_data),.io_async_ridx(auto_in_a_ridx),.io_async_widx(auto_in_a_widx),.io_async_safe_ridx_valid(auto_in_a_safe_ridx_valid),.io_async_safe_widx_valid(auto_in_a_safe_widx_valid),.io_async_safe_source_reset_n(auto_in_a_safe_source_reset_n),.io_async_safe_sink_reset_n(auto_in_a_safe_sink_reset_n)); 
  AsyncQueueSource_2 nodeIn_d_source(.clock(clock),.reset(reset),.io_enq_ready(auto_out_d_ready),.io_enq_valid(auto_out_d_valid),.io_enq_bits_opcode(auto_out_d_bits_opcode),.io_enq_bits_size(auto_out_d_bits_size),.io_enq_bits_source(auto_out_d_bits_source),.io_enq_bits_data(auto_out_d_bits_data),.io_async_mem_0_opcode(auto_in_d_mem_0_opcode),.io_async_mem_0_size(auto_in_d_mem_0_size),.io_async_mem_0_source(auto_in_d_mem_0_source),.io_async_mem_0_data(auto_in_d_mem_0_data),.io_async_ridx(auto_in_d_ridx),.io_async_widx(auto_in_d_widx),.io_async_safe_ridx_valid(auto_in_d_safe_ridx_valid),.io_async_safe_widx_valid(auto_in_d_safe_widx_valid),.io_async_safe_source_reset_n(auto_in_d_safe_source_reset_n),.io_async_safe_sink_reset_n(auto_in_d_safe_sink_reset_n)); 
endmodule
 
module ClockCrossingReg_w15 (
  input clock,
  input [14:0] io_d,
  output [14:0] io_q,
  input io_en) ; 
   reg [14:0] cdc_reg ;  
  always @( posedge clock)
       begin 
         if (io_en)
            cdc_reg <=io_d;
       end
  
  assign io_q=cdc_reg; 
endmodule
 
module AsyncQueueSink_2 (
  input clock,
  input reset,
  output io_deq_valid,
  output io_deq_bits_resumereq,
  output [9:0] io_deq_bits_hartsel,
  output io_deq_bits_ackhavereset,
  output io_deq_bits_hrmask_0,
  input io_async_mem_resumereq_0,
  input [9:0] io_async_mem_hartsel_0,
  input io_async_mem_ackhavereset_0,
  input io_async_mem_hrmask_0_0,
  output io_async_ridx,
  input io_async_widx,
  output io_async_safe_ridx_valid,
  input io_async_safe_widx_valid,
  input io_async_safe_source_reset_n,
  output io_async_safe_sink_reset_n) ; 
   wire io_deq_valid_0 ;  
   wire _source_valid_io_out ;  
   wire _source_extend_io_out ;  
   wire _sink_valid_0_io_out ;  
   wire [14:0] _io_deq_bits_deq_bits_reg_io_q ;  
   wire _widx_widx_gray_io_q ;  
   reg ridx_ridx_bin ;  
   wire ridx=_source_valid_io_out&ridx_ridx_bin+io_deq_valid_0 ;  
   wire valid=_source_valid_io_out&ridx!=_widx_widx_gray_io_q ;  
   reg valid_reg ;  
  assign io_deq_valid_0=valid_reg&_source_valid_io_out; 
   reg ridx_gray ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            begin 
              ridx_ridx_bin <=1'h0;
              valid_reg <=1'h0;
              ridx_gray <=1'h0;
            end 
          else 
            begin 
              ridx_ridx_bin <=ridx;
              valid_reg <=valid;
              ridx_gray <=ridx;
            end 
       end
  
  AsyncResetSynchronizerShiftReg_w1_d3_i0 widx_widx_gray(.clock(clock),.reset(reset),.io_d(io_async_widx),.io_q(_widx_widx_gray_io_q)); 
  ClockCrossingReg_w15 io_deq_bits_deq_bits_reg(.clock(clock),.io_d({io_async_mem_resumereq_0,io_async_mem_hartsel_0,io_async_mem_ackhavereset_0,2'h0,io_async_mem_hrmask_0_0}),.io_q(_io_deq_bits_deq_bits_reg_io_q),.io_en(valid)); 
  AsyncValidSync sink_valid_0(.io_in(1'h1),.io_out(_sink_valid_0_io_out),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync sink_valid_1(.io_in(_sink_valid_0_io_out),.io_out(io_async_safe_ridx_valid),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync source_extend(.io_in(io_async_safe_widx_valid),.io_out(_source_extend_io_out),.clock(clock),.reset(reset|~io_async_safe_source_reset_n)); 
  AsyncValidSync source_valid(.io_in(_source_extend_io_out),.io_out(_source_valid_io_out),.clock(clock),.reset(reset)); 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_resumereq=_io_deq_bits_deq_bits_reg_io_q[14]; 
  assign io_deq_bits_hartsel=_io_deq_bits_deq_bits_reg_io_q[13:4]; 
  assign io_deq_bits_ackhavereset=_io_deq_bits_deq_bits_reg_io_q[3]; 
  assign io_deq_bits_hrmask_0=_io_deq_bits_deq_bits_reg_io_q[0]; 
  assign io_async_ridx=ridx_gray; 
  assign io_async_safe_sink_reset_n=~reset; 
endmodule
 
module TLDebugModuleInnerAsync (
  input [2:0] auto_dmiXing_in_a_mem_0_opcode,
  input [8:0] auto_dmiXing_in_a_mem_0_address,
  input [31:0] auto_dmiXing_in_a_mem_0_data,
  output auto_dmiXing_in_a_ridx,
  input auto_dmiXing_in_a_widx,
  output auto_dmiXing_in_a_safe_ridx_valid,
  input auto_dmiXing_in_a_safe_widx_valid,
  input auto_dmiXing_in_a_safe_source_reset_n,
  output auto_dmiXing_in_a_safe_sink_reset_n,
  output [2:0] auto_dmiXing_in_d_mem_0_opcode,
  output [1:0] auto_dmiXing_in_d_mem_0_size,
  output auto_dmiXing_in_d_mem_0_source,
  output [31:0] auto_dmiXing_in_d_mem_0_data,
  input auto_dmiXing_in_d_ridx,
  output auto_dmiXing_in_d_widx,
  input auto_dmiXing_in_d_safe_ridx_valid,
  output auto_dmiXing_in_d_safe_widx_valid,
  output auto_dmiXing_in_d_safe_source_reset_n,
  input auto_dmiXing_in_d_safe_sink_reset_n,
  output auto_dmInner_tl_in_a_ready,
  input auto_dmInner_tl_in_a_valid,
  input [2:0] auto_dmInner_tl_in_a_bits_opcode,
  input [2:0] auto_dmInner_tl_in_a_bits_param,
  input [1:0] auto_dmInner_tl_in_a_bits_size,
  input [8:0] auto_dmInner_tl_in_a_bits_source,
  input [11:0] auto_dmInner_tl_in_a_bits_address,
  input [7:0] auto_dmInner_tl_in_a_bits_mask,
  input [63:0] auto_dmInner_tl_in_a_bits_data,
  input auto_dmInner_tl_in_a_bits_corrupt,
  input auto_dmInner_tl_in_d_ready,
  output auto_dmInner_tl_in_d_valid,
  output [2:0] auto_dmInner_tl_in_d_bits_opcode,
  output [1:0] auto_dmInner_tl_in_d_bits_size,
  output [8:0] auto_dmInner_tl_in_d_bits_source,
  output [63:0] auto_dmInner_tl_in_d_bits_data,
  input io_debug_clock,
  input io_debug_reset,
  input io_dmactive,
  input io_innerCtrl_mem_resumereq_0,
  input [9:0] io_innerCtrl_mem_hartsel_0,
  input io_innerCtrl_mem_ackhavereset_0,
  input io_innerCtrl_mem_hrmask_0_0,
  output io_innerCtrl_ridx,
  input io_innerCtrl_widx,
  output io_innerCtrl_safe_ridx_valid,
  input io_innerCtrl_safe_widx_valid,
  input io_innerCtrl_safe_source_reset_n,
  output io_innerCtrl_safe_sink_reset_n,
  output io_hgDebugInt_0,
  input io_hartIsInReset_0) ; 
   wire _dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_valid ;  
   wire _dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_resumereq ;  
   wire [9:0] _dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hartsel ;  
   wire _dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_ackhavereset ;  
   wire _dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hrmask_0 ;  
   wire _dmactive_synced_dmactive_synced_dmactiveSync_io_q ;  
   wire _dmiXing_auto_out_a_valid ;  
   wire [2:0] _dmiXing_auto_out_a_bits_opcode ;  
   wire [2:0] _dmiXing_auto_out_a_bits_param ;  
   wire [1:0] _dmiXing_auto_out_a_bits_size ;  
   wire _dmiXing_auto_out_a_bits_source ;  
   wire [8:0] _dmiXing_auto_out_a_bits_address ;  
   wire [3:0] _dmiXing_auto_out_a_bits_mask ;  
   wire [31:0] _dmiXing_auto_out_a_bits_data ;  
   wire _dmiXing_auto_out_a_bits_corrupt ;  
   wire _dmiXing_auto_out_d_ready ;  
   wire _dmInner_auto_dmi_in_a_ready ;  
   wire _dmInner_auto_dmi_in_d_valid ;  
   wire [2:0] _dmInner_auto_dmi_in_d_bits_opcode ;  
   wire [1:0] _dmInner_auto_dmi_in_d_bits_size ;  
   wire _dmInner_auto_dmi_in_d_bits_source ;  
   wire [31:0] _dmInner_auto_dmi_in_d_bits_data ;  
  TLDebugModuleInner dmInner(.clock(io_debug_clock),.reset(io_debug_reset),.auto_tl_in_a_ready(auto_dmInner_tl_in_a_ready),.auto_tl_in_a_valid(auto_dmInner_tl_in_a_valid),.auto_tl_in_a_bits_opcode(auto_dmInner_tl_in_a_bits_opcode),.auto_tl_in_a_bits_param(auto_dmInner_tl_in_a_bits_param),.auto_tl_in_a_bits_size(auto_dmInner_tl_in_a_bits_size),.auto_tl_in_a_bits_source(auto_dmInner_tl_in_a_bits_source),.auto_tl_in_a_bits_address(auto_dmInner_tl_in_a_bits_address),.auto_tl_in_a_bits_mask(auto_dmInner_tl_in_a_bits_mask),.auto_tl_in_a_bits_data(auto_dmInner_tl_in_a_bits_data),.auto_tl_in_a_bits_corrupt(auto_dmInner_tl_in_a_bits_corrupt),.auto_tl_in_d_ready(auto_dmInner_tl_in_d_ready),.auto_tl_in_d_valid(auto_dmInner_tl_in_d_valid),.auto_tl_in_d_bits_opcode(auto_dmInner_tl_in_d_bits_opcode),.auto_tl_in_d_bits_size(auto_dmInner_tl_in_d_bits_size),.auto_tl_in_d_bits_source(auto_dmInner_tl_in_d_bits_source),.auto_tl_in_d_bits_data(auto_dmInner_tl_in_d_bits_data),.auto_dmi_in_a_ready(_dmInner_auto_dmi_in_a_ready),.auto_dmi_in_a_valid(_dmiXing_auto_out_a_valid),.auto_dmi_in_a_bits_opcode(_dmiXing_auto_out_a_bits_opcode),.auto_dmi_in_a_bits_param(_dmiXing_auto_out_a_bits_param),.auto_dmi_in_a_bits_size(_dmiXing_auto_out_a_bits_size),.auto_dmi_in_a_bits_source(_dmiXing_auto_out_a_bits_source),.auto_dmi_in_a_bits_address(_dmiXing_auto_out_a_bits_address),.auto_dmi_in_a_bits_mask(_dmiXing_auto_out_a_bits_mask),.auto_dmi_in_a_bits_data(_dmiXing_auto_out_a_bits_data),.auto_dmi_in_a_bits_corrupt(_dmiXing_auto_out_a_bits_corrupt),.auto_dmi_in_d_ready(_dmiXing_auto_out_d_ready),.auto_dmi_in_d_valid(_dmInner_auto_dmi_in_d_valid),.auto_dmi_in_d_bits_opcode(_dmInner_auto_dmi_in_d_bits_opcode),.auto_dmi_in_d_bits_size(_dmInner_auto_dmi_in_d_bits_size),.auto_dmi_in_d_bits_source(_dmInner_auto_dmi_in_d_bits_source),.auto_dmi_in_d_bits_data(_dmInner_auto_dmi_in_d_bits_data),.io_dmactive(_dmactive_synced_dmactive_synced_dmactiveSync_io_q),.io_innerCtrl_valid(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_valid),.io_innerCtrl_bits_resumereq(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_resumereq),.io_innerCtrl_bits_hartsel(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hartsel),.io_innerCtrl_bits_ackhavereset(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_ackhavereset),.io_innerCtrl_bits_hrmask_0(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hrmask_0),.io_hgDebugInt_0(io_hgDebugInt_0),.io_hartIsInReset_0(io_hartIsInReset_0)); 
  TLAsyncCrossingSink dmiXing(.clock(io_debug_clock),.reset(io_debug_reset),.auto_in_a_mem_0_opcode(auto_dmiXing_in_a_mem_0_opcode),.auto_in_a_mem_0_address(auto_dmiXing_in_a_mem_0_address),.auto_in_a_mem_0_data(auto_dmiXing_in_a_mem_0_data),.auto_in_a_ridx(auto_dmiXing_in_a_ridx),.auto_in_a_widx(auto_dmiXing_in_a_widx),.auto_in_a_safe_ridx_valid(auto_dmiXing_in_a_safe_ridx_valid),.auto_in_a_safe_widx_valid(auto_dmiXing_in_a_safe_widx_valid),.auto_in_a_safe_source_reset_n(auto_dmiXing_in_a_safe_source_reset_n),.auto_in_a_safe_sink_reset_n(auto_dmiXing_in_a_safe_sink_reset_n),.auto_in_d_mem_0_opcode(auto_dmiXing_in_d_mem_0_opcode),.auto_in_d_mem_0_size(auto_dmiXing_in_d_mem_0_size),.auto_in_d_mem_0_source(auto_dmiXing_in_d_mem_0_source),.auto_in_d_mem_0_data(auto_dmiXing_in_d_mem_0_data),.auto_in_d_ridx(auto_dmiXing_in_d_ridx),.auto_in_d_widx(auto_dmiXing_in_d_widx),.auto_in_d_safe_ridx_valid(auto_dmiXing_in_d_safe_ridx_valid),.auto_in_d_safe_widx_valid(auto_dmiXing_in_d_safe_widx_valid),.auto_in_d_safe_source_reset_n(auto_dmiXing_in_d_safe_source_reset_n),.auto_in_d_safe_sink_reset_n(auto_dmiXing_in_d_safe_sink_reset_n),.auto_out_a_ready(_dmInner_auto_dmi_in_a_ready),.auto_out_a_valid(_dmiXing_auto_out_a_valid),.auto_out_a_bits_opcode(_dmiXing_auto_out_a_bits_opcode),.auto_out_a_bits_param(_dmiXing_auto_out_a_bits_param),.auto_out_a_bits_size(_dmiXing_auto_out_a_bits_size),.auto_out_a_bits_source(_dmiXing_auto_out_a_bits_source),.auto_out_a_bits_address(_dmiXing_auto_out_a_bits_address),.auto_out_a_bits_mask(_dmiXing_auto_out_a_bits_mask),.auto_out_a_bits_data(_dmiXing_auto_out_a_bits_data),.auto_out_a_bits_corrupt(_dmiXing_auto_out_a_bits_corrupt),.auto_out_d_ready(_dmiXing_auto_out_d_ready),.auto_out_d_valid(_dmInner_auto_dmi_in_d_valid),.auto_out_d_bits_opcode(_dmInner_auto_dmi_in_d_bits_opcode),.auto_out_d_bits_size(_dmInner_auto_dmi_in_d_bits_size),.auto_out_d_bits_source(_dmInner_auto_dmi_in_d_bits_source),.auto_out_d_bits_data(_dmInner_auto_dmi_in_d_bits_data)); 
  AsyncResetSynchronizerShiftReg_w1_d3_i0 dmactive_synced_dmactive_synced_dmactiveSync(.clock(io_debug_clock),.reset(io_debug_reset),.io_d(io_dmactive),.io_q(_dmactive_synced_dmactive_synced_dmactiveSync_io_q)); 
  AsyncQueueSink_2 dmactive_synced_dmInner_io_innerCtrl_sink(.clock(io_debug_clock),.reset(io_debug_reset),.io_deq_valid(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_valid),.io_deq_bits_resumereq(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_resumereq),.io_deq_bits_hartsel(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hartsel),.io_deq_bits_ackhavereset(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_ackhavereset),.io_deq_bits_hrmask_0(_dmactive_synced_dmInner_io_innerCtrl_sink_io_deq_bits_hrmask_0),.io_async_mem_resumereq_0(io_innerCtrl_mem_resumereq_0),.io_async_mem_hartsel_0(io_innerCtrl_mem_hartsel_0),.io_async_mem_ackhavereset_0(io_innerCtrl_mem_ackhavereset_0),.io_async_mem_hrmask_0_0(io_innerCtrl_mem_hrmask_0_0),.io_async_ridx(io_innerCtrl_ridx),.io_async_widx(io_innerCtrl_widx),.io_async_safe_ridx_valid(io_innerCtrl_safe_ridx_valid),.io_async_safe_widx_valid(io_innerCtrl_safe_widx_valid),.io_async_safe_source_reset_n(io_innerCtrl_safe_source_reset_n),.io_async_safe_sink_reset_n(io_innerCtrl_safe_sink_reset_n)); 
endmodule
 
module TLDebugModule (
  output auto_dmInner_dmInner_tl_in_a_ready,
  input auto_dmInner_dmInner_tl_in_a_valid,
  input [2:0] auto_dmInner_dmInner_tl_in_a_bits_opcode,
  input [2:0] auto_dmInner_dmInner_tl_in_a_bits_param,
  input [1:0] auto_dmInner_dmInner_tl_in_a_bits_size,
  input [8:0] auto_dmInner_dmInner_tl_in_a_bits_source,
  input [11:0] auto_dmInner_dmInner_tl_in_a_bits_address,
  input [7:0] auto_dmInner_dmInner_tl_in_a_bits_mask,
  input [63:0] auto_dmInner_dmInner_tl_in_a_bits_data,
  input auto_dmInner_dmInner_tl_in_a_bits_corrupt,
  input auto_dmInner_dmInner_tl_in_d_ready,
  output auto_dmInner_dmInner_tl_in_d_valid,
  output [2:0] auto_dmInner_dmInner_tl_in_d_bits_opcode,
  output [1:0] auto_dmInner_dmInner_tl_in_d_bits_size,
  output [8:0] auto_dmInner_dmInner_tl_in_d_bits_source,
  output [63:0] auto_dmInner_dmInner_tl_in_d_bits_data,
  output auto_dmOuter_intsource_out_sync_0,
  input io_debug_clock,
  input io_debug_reset,
  output io_ctrl_ndreset,
  output io_ctrl_dmactive,
  input io_ctrl_dmactiveAck,
  output io_dmi_dmi_req_ready,
  input io_dmi_dmi_req_valid,
  input [6:0] io_dmi_dmi_req_bits_addr,
  input [31:0] io_dmi_dmi_req_bits_data,
  input [1:0] io_dmi_dmi_req_bits_op,
  input io_dmi_dmi_resp_ready,
  output io_dmi_dmi_resp_valid,
  output [31:0] io_dmi_dmi_resp_bits_data,
  output [1:0] io_dmi_dmi_resp_bits_resp,
  input io_dmi_dmiClock,
  input io_dmi_dmiReset,
  input io_hartIsInReset_0) ; 
   wire _dmInner_auto_dmiXing_in_a_ridx ;  
   wire _dmInner_auto_dmiXing_in_a_safe_ridx_valid ;  
   wire _dmInner_auto_dmiXing_in_a_safe_sink_reset_n ;  
   wire [2:0] _dmInner_auto_dmiXing_in_d_mem_0_opcode ;  
   wire [1:0] _dmInner_auto_dmiXing_in_d_mem_0_size ;  
   wire _dmInner_auto_dmiXing_in_d_mem_0_source ;  
   wire [31:0] _dmInner_auto_dmiXing_in_d_mem_0_data ;  
   wire _dmInner_auto_dmiXing_in_d_widx ;  
   wire _dmInner_auto_dmiXing_in_d_safe_widx_valid ;  
   wire _dmInner_auto_dmiXing_in_d_safe_source_reset_n ;  
   wire _dmInner_io_innerCtrl_ridx ;  
   wire _dmInner_io_innerCtrl_safe_ridx_valid ;  
   wire _dmInner_io_innerCtrl_safe_sink_reset_n ;  
   wire _dmInner_io_hgDebugInt_0 ;  
   wire [2:0] _dmOuter_auto_asource_out_a_mem_0_opcode ;  
   wire [8:0] _dmOuter_auto_asource_out_a_mem_0_address ;  
   wire [31:0] _dmOuter_auto_asource_out_a_mem_0_data ;  
   wire _dmOuter_auto_asource_out_a_widx ;  
   wire _dmOuter_auto_asource_out_a_safe_widx_valid ;  
   wire _dmOuter_auto_asource_out_a_safe_source_reset_n ;  
   wire _dmOuter_auto_asource_out_d_ridx ;  
   wire _dmOuter_auto_asource_out_d_safe_ridx_valid ;  
   wire _dmOuter_auto_asource_out_d_safe_sink_reset_n ;  
   wire _dmOuter_io_ctrl_dmactive ;  
   wire _dmOuter_io_innerCtrl_mem_resumereq_0 ;  
   wire [9:0] _dmOuter_io_innerCtrl_mem_hartsel_0 ;  
   wire _dmOuter_io_innerCtrl_mem_ackhavereset_0 ;  
   wire _dmOuter_io_innerCtrl_mem_hrmask_0_0 ;  
   wire _dmOuter_io_innerCtrl_widx ;  
   wire _dmOuter_io_innerCtrl_safe_widx_valid ;  
   wire _dmOuter_io_innerCtrl_safe_source_reset_n ;  
  TLDebugModuleOuterAsync dmOuter(.auto_asource_out_a_mem_0_opcode(_dmOuter_auto_asource_out_a_mem_0_opcode),.auto_asource_out_a_mem_0_address(_dmOuter_auto_asource_out_a_mem_0_address),.auto_asource_out_a_mem_0_data(_dmOuter_auto_asource_out_a_mem_0_data),.auto_asource_out_a_ridx(_dmInner_auto_dmiXing_in_a_ridx),.auto_asource_out_a_widx(_dmOuter_auto_asource_out_a_widx),.auto_asource_out_a_safe_ridx_valid(_dmInner_auto_dmiXing_in_a_safe_ridx_valid),.auto_asource_out_a_safe_widx_valid(_dmOuter_auto_asource_out_a_safe_widx_valid),.auto_asource_out_a_safe_source_reset_n(_dmOuter_auto_asource_out_a_safe_source_reset_n),.auto_asource_out_a_safe_sink_reset_n(_dmInner_auto_dmiXing_in_a_safe_sink_reset_n),.auto_asource_out_d_mem_0_opcode(_dmInner_auto_dmiXing_in_d_mem_0_opcode),.auto_asource_out_d_mem_0_size(_dmInner_auto_dmiXing_in_d_mem_0_size),.auto_asource_out_d_mem_0_source(_dmInner_auto_dmiXing_in_d_mem_0_source),.auto_asource_out_d_mem_0_data(_dmInner_auto_dmiXing_in_d_mem_0_data),.auto_asource_out_d_ridx(_dmOuter_auto_asource_out_d_ridx),.auto_asource_out_d_widx(_dmInner_auto_dmiXing_in_d_widx),.auto_asource_out_d_safe_ridx_valid(_dmOuter_auto_asource_out_d_safe_ridx_valid),.auto_asource_out_d_safe_widx_valid(_dmInner_auto_dmiXing_in_d_safe_widx_valid),.auto_asource_out_d_safe_source_reset_n(_dmInner_auto_dmiXing_in_d_safe_source_reset_n),.auto_asource_out_d_safe_sink_reset_n(_dmOuter_auto_asource_out_d_safe_sink_reset_n),.auto_intsource_out_sync_0(auto_dmOuter_intsource_out_sync_0),.io_dmi_clock(io_dmi_dmiClock),.io_dmi_reset(io_dmi_dmiReset),.io_dmi_req_ready(io_dmi_dmi_req_ready),.io_dmi_req_valid(io_dmi_dmi_req_valid),.io_dmi_req_bits_addr(io_dmi_dmi_req_bits_addr),.io_dmi_req_bits_data(io_dmi_dmi_req_bits_data),.io_dmi_req_bits_op(io_dmi_dmi_req_bits_op),.io_dmi_resp_ready(io_dmi_dmi_resp_ready),.io_dmi_resp_valid(io_dmi_dmi_resp_valid),.io_dmi_resp_bits_data(io_dmi_dmi_resp_bits_data),.io_dmi_resp_bits_resp(io_dmi_dmi_resp_bits_resp),.io_ctrl_ndreset(io_ctrl_ndreset),.io_ctrl_dmactive(_dmOuter_io_ctrl_dmactive),.io_ctrl_dmactiveAck(io_ctrl_dmactiveAck),.io_innerCtrl_mem_resumereq_0(_dmOuter_io_innerCtrl_mem_resumereq_0),.io_innerCtrl_mem_hartsel_0(_dmOuter_io_innerCtrl_mem_hartsel_0),.io_innerCtrl_mem_ackhavereset_0(_dmOuter_io_innerCtrl_mem_ackhavereset_0),.io_innerCtrl_mem_hrmask_0_0(_dmOuter_io_innerCtrl_mem_hrmask_0_0),.io_innerCtrl_ridx(_dmInner_io_innerCtrl_ridx),.io_innerCtrl_widx(_dmOuter_io_innerCtrl_widx),.io_innerCtrl_safe_ridx_valid(_dmInner_io_innerCtrl_safe_ridx_valid),.io_innerCtrl_safe_widx_valid(_dmOuter_io_innerCtrl_safe_widx_valid),.io_innerCtrl_safe_source_reset_n(_dmOuter_io_innerCtrl_safe_source_reset_n),.io_innerCtrl_safe_sink_reset_n(_dmInner_io_innerCtrl_safe_sink_reset_n),.io_hgDebugInt_0(_dmInner_io_hgDebugInt_0)); 
  TLDebugModuleInnerAsync dmInner(.auto_dmiXing_in_a_mem_0_opcode(_dmOuter_auto_asource_out_a_mem_0_opcode),.auto_dmiXing_in_a_mem_0_address(_dmOuter_auto_asource_out_a_mem_0_address),.auto_dmiXing_in_a_mem_0_data(_dmOuter_auto_asource_out_a_mem_0_data),.auto_dmiXing_in_a_ridx(_dmInner_auto_dmiXing_in_a_ridx),.auto_dmiXing_in_a_widx(_dmOuter_auto_asource_out_a_widx),.auto_dmiXing_in_a_safe_ridx_valid(_dmInner_auto_dmiXing_in_a_safe_ridx_valid),.auto_dmiXing_in_a_safe_widx_valid(_dmOuter_auto_asource_out_a_safe_widx_valid),.auto_dmiXing_in_a_safe_source_reset_n(_dmOuter_auto_asource_out_a_safe_source_reset_n),.auto_dmiXing_in_a_safe_sink_reset_n(_dmInner_auto_dmiXing_in_a_safe_sink_reset_n),.auto_dmiXing_in_d_mem_0_opcode(_dmInner_auto_dmiXing_in_d_mem_0_opcode),.auto_dmiXing_in_d_mem_0_size(_dmInner_auto_dmiXing_in_d_mem_0_size),.auto_dmiXing_in_d_mem_0_source(_dmInner_auto_dmiXing_in_d_mem_0_source),.auto_dmiXing_in_d_mem_0_data(_dmInner_auto_dmiXing_in_d_mem_0_data),.auto_dmiXing_in_d_ridx(_dmOuter_auto_asource_out_d_ridx),.auto_dmiXing_in_d_widx(_dmInner_auto_dmiXing_in_d_widx),.auto_dmiXing_in_d_safe_ridx_valid(_dmOuter_auto_asource_out_d_safe_ridx_valid),.auto_dmiXing_in_d_safe_widx_valid(_dmInner_auto_dmiXing_in_d_safe_widx_valid),.auto_dmiXing_in_d_safe_source_reset_n(_dmInner_auto_dmiXing_in_d_safe_source_reset_n),.auto_dmiXing_in_d_safe_sink_reset_n(_dmOuter_auto_asource_out_d_safe_sink_reset_n),.auto_dmInner_tl_in_a_ready(auto_dmInner_dmInner_tl_in_a_ready),.auto_dmInner_tl_in_a_valid(auto_dmInner_dmInner_tl_in_a_valid),.auto_dmInner_tl_in_a_bits_opcode(auto_dmInner_dmInner_tl_in_a_bits_opcode),.auto_dmInner_tl_in_a_bits_param(auto_dmInner_dmInner_tl_in_a_bits_param),.auto_dmInner_tl_in_a_bits_size(auto_dmInner_dmInner_tl_in_a_bits_size),.auto_dmInner_tl_in_a_bits_source(auto_dmInner_dmInner_tl_in_a_bits_source),.auto_dmInner_tl_in_a_bits_address(auto_dmInner_dmInner_tl_in_a_bits_address),.auto_dmInner_tl_in_a_bits_mask(auto_dmInner_dmInner_tl_in_a_bits_mask),.auto_dmInner_tl_in_a_bits_data(auto_dmInner_dmInner_tl_in_a_bits_data),.auto_dmInner_tl_in_a_bits_corrupt(auto_dmInner_dmInner_tl_in_a_bits_corrupt),.auto_dmInner_tl_in_d_ready(auto_dmInner_dmInner_tl_in_d_ready),.auto_dmInner_tl_in_d_valid(auto_dmInner_dmInner_tl_in_d_valid),.auto_dmInner_tl_in_d_bits_opcode(auto_dmInner_dmInner_tl_in_d_bits_opcode),.auto_dmInner_tl_in_d_bits_size(auto_dmInner_dmInner_tl_in_d_bits_size),.auto_dmInner_tl_in_d_bits_source(auto_dmInner_dmInner_tl_in_d_bits_source),.auto_dmInner_tl_in_d_bits_data(auto_dmInner_dmInner_tl_in_d_bits_data),.io_debug_clock(io_debug_clock),.io_debug_reset(io_debug_reset),.io_dmactive(_dmOuter_io_ctrl_dmactive),.io_innerCtrl_mem_resumereq_0(_dmOuter_io_innerCtrl_mem_resumereq_0),.io_innerCtrl_mem_hartsel_0(_dmOuter_io_innerCtrl_mem_hartsel_0),.io_innerCtrl_mem_ackhavereset_0(_dmOuter_io_innerCtrl_mem_ackhavereset_0),.io_innerCtrl_mem_hrmask_0_0(_dmOuter_io_innerCtrl_mem_hrmask_0_0),.io_innerCtrl_ridx(_dmInner_io_innerCtrl_ridx),.io_innerCtrl_widx(_dmOuter_io_innerCtrl_widx),.io_innerCtrl_safe_ridx_valid(_dmInner_io_innerCtrl_safe_ridx_valid),.io_innerCtrl_safe_widx_valid(_dmOuter_io_innerCtrl_safe_widx_valid),.io_innerCtrl_safe_source_reset_n(_dmOuter_io_innerCtrl_safe_source_reset_n),.io_innerCtrl_safe_sink_reset_n(_dmInner_io_innerCtrl_safe_sink_reset_n),.io_hgDebugInt_0(_dmInner_io_hgDebugInt_0),.io_hartIsInReset_0(io_hartIsInReset_0)); 
  assign io_ctrl_dmactive=_dmOuter_io_ctrl_dmactive; 
endmodule
 
module AsyncResetRegVec_w2_i0 (
  input clock,
  input reset,
  input [1:0] io_d,
  output [1:0] io_q) ; 
   reg [1:0] reg_0 ;  
  always @(  posedge clock or  posedge reset)
       begin 
         if (reset)
            reg_0 <=2'h0;
          else 
            reg_0 <=io_d;
       end
  
  assign io_q=reg_0; 
endmodule
 
module IntSyncCrossingSource_5 (
  input clock,
  input reset,
  input auto_in_0,
  input auto_in_1,
  output auto_out_sync_0,
  output auto_out_sync_1) ; 
   wire [1:0] _reg_io_q ;  
  AsyncResetRegVec_w2_i0 reg_0(.clock(clock),.reset(reset),.io_d({auto_in_1,auto_in_0}),.io_q(_reg_io_q)); 
  assign auto_out_sync_0=_reg_io_q[0]; 
  assign auto_out_sync_1=_reg_io_q[1]; 
endmodule
 
module TLMonitor_35 (
  input clock,
  input reset,
  input io_in_a_ready,
  input io_in_a_valid,
  input [2:0] io_in_a_bits_opcode,
  input [2:0] io_in_a_bits_param,
  input [1:0] io_in_a_bits_size,
  input [8:0] io_in_a_bits_source,
  input [16:0] io_in_a_bits_address,
  input [7:0] io_in_a_bits_mask,
  input io_in_a_bits_corrupt,
  input io_in_d_ready,
  input io_in_d_valid,
  input [1:0] io_in_d_bits_size,
  input [8:0] io_in_d_bits_source) ; 
   wire [31:0] _plusarg_reader_out ;  
   wire a_first_done=io_in_a_ready&io_in_a_valid ;  
   reg a_first_counter ;  
   reg [2:0] opcode ;  
   reg [2:0] param ;  
   reg [1:0] size ;  
   reg [8:0] source ;  
   reg [16:0] address ;  
   reg d_first_counter ;  
   reg [1:0] size_1 ;  
   reg [8:0] source_1 ;  
   reg [303:0] inflight ;  
   reg [1215:0] inflight_opcodes ;  
   reg [1215:0] inflight_sizes ;  
   reg a_first_counter_1 ;  
   reg d_first_counter_1 ;  
   wire [1215:0] _GEN={1205'h0,io_in_d_bits_source,2'h0} ;  
   wire [1215:0] _a_opcode_lookup_T_1=inflight_opcodes>>_GEN ;  
   wire _GEN_0=a_first_done&~a_first_counter_1 ;  
   reg [2:0] casez_tmp ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp =3'h0;
          3 'b001:
             casez_tmp =3'h0;
          3 'b010:
             casez_tmp =3'h1;
          3 'b011:
             casez_tmp =3'h1;
          3 'b100:
             casez_tmp =3'h1;
          3 'b101:
             casez_tmp =3'h2;
          3 'b110:
             casez_tmp =3'h4;
          default :
             casez_tmp =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_0 ;  
  always @(*)
       begin 
         casez (io_in_a_bits_opcode)
          3 'b000:
             casez_tmp_0 =3'h0;
          3 'b001:
             casez_tmp_0 =3'h0;
          3 'b010:
             casez_tmp_0 =3'h1;
          3 'b011:
             casez_tmp_0 =3'h1;
          3 'b100:
             casez_tmp_0 =3'h1;
          3 'b101:
             casez_tmp_0 =3'h2;
          3 'b110:
             casez_tmp_0 =3'h5;
          default :
             casez_tmp_0 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_1 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_1 =3'h0;
          3 'b001:
             casez_tmp_1 =3'h0;
          3 'b010:
             casez_tmp_1 =3'h1;
          3 'b011:
             casez_tmp_1 =3'h1;
          3 'b100:
             casez_tmp_1 =3'h1;
          3 'b101:
             casez_tmp_1 =3'h2;
          3 'b110:
             casez_tmp_1 =3'h4;
          default :
             casez_tmp_1 =3'h4;
         endcase 
       end
  
   reg [2:0] casez_tmp_2 ;  
  always @(*)
       begin 
         casez (_a_opcode_lookup_T_1[3:1])
          3 'b000:
             casez_tmp_2 =3'h0;
          3 'b001:
             casez_tmp_2 =3'h0;
          3 'b010:
             casez_tmp_2 =3'h1;
          3 'b011:
             casez_tmp_2 =3'h1;
          3 'b100:
             casez_tmp_2 =3'h1;
          3 'b101:
             casez_tmp_2 =3'h2;
          3 'b110:
             casez_tmp_2 =3'h5;
          default :
             casez_tmp_2 =3'h4;
         endcase 
       end
  
   reg [31:0] watchdog ;  
   wire [5:0] _is_aligned_mask_T_1=6'h7<<io_in_a_bits_size ;  
   wire [2:0] _GEN_1=io_in_a_bits_address[2:0]&~(_is_aligned_mask_T_1[2:0]) ;  
   wire mask_size=io_in_a_bits_size==2'h2 ;  
   wire mask_acc=(&io_in_a_bits_size)|mask_size&~(io_in_a_bits_address[2]) ;  
   wire mask_acc_1=(&io_in_a_bits_size)|mask_size&io_in_a_bits_address[2] ;  
   wire mask_size_1=io_in_a_bits_size==2'h1 ;  
   wire mask_eq_2=~(io_in_a_bits_address[2])&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_2=mask_acc|mask_size_1&mask_eq_2 ;  
   wire mask_eq_3=~(io_in_a_bits_address[2])&io_in_a_bits_address[1] ;  
   wire mask_acc_3=mask_acc|mask_size_1&mask_eq_3 ;  
   wire mask_eq_4=io_in_a_bits_address[2]&~(io_in_a_bits_address[1]) ;  
   wire mask_acc_4=mask_acc_1|mask_size_1&mask_eq_4 ;  
   wire mask_eq_5=io_in_a_bits_address[2]&io_in_a_bits_address[1] ;  
   wire mask_acc_5=mask_acc_1|mask_size_1&mask_eq_5 ;  
   wire [7:0] mask={mask_acc_5|mask_eq_5&io_in_a_bits_address[0],mask_acc_5|mask_eq_5&~(io_in_a_bits_address[0]),mask_acc_4|mask_eq_4&io_in_a_bits_address[0],mask_acc_4|mask_eq_4&~(io_in_a_bits_address[0]),mask_acc_3|mask_eq_3&io_in_a_bits_address[0],mask_acc_3|mask_eq_3&~(io_in_a_bits_address[0]),mask_acc_2|mask_eq_2&io_in_a_bits_address[0],mask_acc_2|mask_eq_2&~(io_in_a_bits_address[0])} ;  
   wire _GEN_2=io_in_a_valid&io_in_a_bits_opcode==3'h6&~reset ;  
   wire _GEN_3=io_in_a_bits_source>9'h12F ;  
   wire _GEN_4=io_in_a_bits_param>3'h2 ;  
   wire _GEN_5=io_in_a_bits_mask!=8'hFF ;  
   wire _GEN_6=io_in_a_valid&(&io_in_a_bits_opcode)&~reset ;  
   wire _GEN_7=io_in_a_valid&io_in_a_bits_opcode==3'h4&~reset ;  
   wire _GEN_8=_GEN_7&_GEN_3 ;  
   wire _GEN_9=io_in_a_bits_mask!=mask ;  
   wire _GEN_10=io_in_a_valid&io_in_a_bits_opcode==3'h0&~reset ;  
   wire _GEN_11=io_in_a_valid&io_in_a_bits_opcode==3'h1&~reset ;  
   wire _GEN_12=io_in_a_valid&io_in_a_bits_opcode==3'h2&~reset ;  
   wire _GEN_13=io_in_a_valid&io_in_a_bits_opcode==3'h3&~reset ;  
   wire _GEN_14=io_in_a_valid&io_in_a_bits_opcode==3'h5&~reset ;  
   wire _GEN_15=io_in_a_valid&a_first_counter&~reset ;  
   wire _GEN_16=io_in_d_valid&d_first_counter&~reset ;  
   wire _GEN_17=io_in_d_valid&~d_first_counter_1 ;  
   wire same_cycle_resp=io_in_a_valid&~a_first_counter_1&io_in_a_bits_source==io_in_d_bits_source ;  
   wire _GEN_18=_GEN_17&same_cycle_resp&~reset ;  
   wire _GEN_19=_GEN_17&~same_cycle_resp&~reset ;  
   wire [303:0] _GEN_20=inflight>>io_in_a_bits_source ;  
   wire [303:0] _GEN_21=inflight>>io_in_d_bits_source ;  
   wire [1215:0] _a_size_lookup_T_1=inflight_sizes>>_GEN ;  
  always @( posedge clock)
       begin 
         if (_GEN_2)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_2&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
              if (1)$display("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(&io_in_a_bits_size))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_4)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&~(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&_GEN_5)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_6&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&~(io_in_a_bits_address[16]))
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_8)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_7&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_10&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|io_in_a_bits_param))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_11&(|(io_in_a_bits_mask&~mask)))
            begin 
              if (1)$display("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&io_in_a_bits_param>3'h4)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_12&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&io_in_a_bits_param[2])
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_13&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14)
            begin 
              if (1)$display("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_3)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|_GEN_1))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&(|(io_in_a_bits_param[2:1])))
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&_GEN_9)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_14&io_in_a_bits_corrupt)
            begin 
              if (1)$display("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (io_in_d_valid&~reset&io_in_d_bits_source>9'h12F)
            begin 
              if (1)$display("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_opcode!=opcode)
            begin 
              if (1)$display("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_param!=param)
            begin 
              if (1)$display("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_size!=size)
            begin 
              if (1)$display("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_source!=source)
            begin 
              if (1)$display("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_15&io_in_a_bits_address!=address)
            begin 
              if (1)$display("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_d_bits_size!=size_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_16&io_in_d_bits_source!=source_1)
            begin 
              if (1)$display("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_0&~reset&_GEN_20[0])
            begin 
              if (1)$display("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~reset&~(_GEN_21[0]|same_cycle_resp))
            begin 
              if (1)$display("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&~(casez_tmp==3'h1|casez_tmp_0==3'h1))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_18&io_in_a_bits_size!=io_in_d_bits_size)
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&~(casez_tmp_1==3'h1|casez_tmp_2==3'h1))
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_19&{2'h0,io_in_d_bits_size}!={1'h0,_a_size_lookup_T_1[3:1]})
            begin 
              if (1)$display("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (_GEN_17&~a_first_counter_1&io_in_a_valid&io_in_a_bits_source==io_in_d_bits_source&~reset&~(~io_in_d_ready|io_in_a_ready))
            begin 
              if (1)$display("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
              if (1)$display("");
            end 
         if (~reset&~(inflight==304'h0|_plusarg_reader_out==32'h0|watchdog<_plusarg_reader_out))
            begin 
              if (1)$display("Assertion failed: TileLink timeout expired (connected at src/main/scala/devices/tilelink/BootROM.scala:86:18)\n    at Monitor.scala:42 assert(cond, message)\n");
              if (1)$display("");
            end 
       end
  
   wire [4110:0] _GEN_22={4100'h0,io_in_d_bits_source,2'h0} ;  
   wire [511:0] _d_clr_T=512'h1<<io_in_d_bits_source ;  
   wire [511:0] _a_set_T=512'h1<<io_in_a_bits_source ;  
   wire [4110:0] _d_opcodes_clr_T_5=4111'hF<<_GEN_22 ;  
   wire [4098:0] _a_opcodes_set_T_1={4095'h0,_GEN_0 ? {io_in_a_bits_opcode,1'h1}:4'h0}<<{4088'h0,io_in_a_bits_source,2'h0} ;  
   wire [4110:0] _d_sizes_clr_T_5=4111'hF<<_GEN_22 ;  
   wire [4097:0] _a_sizes_set_T_1={4095'h0,_GEN_0 ? {io_in_a_bits_size,1'h1}:3'h0}<<{4087'h0,io_in_a_bits_source,2'h0} ;  
   wire d_first_done=io_in_d_ready&io_in_d_valid ;  
   wire _GEN_23=d_first_done&~d_first_counter_1 ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              a_first_counter <=1'h0;
              d_first_counter <=1'h0;
              inflight <=304'h0;
              inflight_opcodes <=1216'h0;
              inflight_sizes <=1216'h0;
              a_first_counter_1 <=1'h0;
              d_first_counter_1 <=1'h0;
              watchdog <=32'h0;
            end 
          else 
            begin 
              a_first_counter <=(~a_first_done|a_first_counter-1'h1)&a_first_counter;
              d_first_counter <=(~d_first_done|d_first_counter-1'h1)&d_first_counter;
              inflight <=(inflight|(_GEN_0 ? _a_set_T[303:0]:304'h0))&~(_GEN_23 ? _d_clr_T[303:0]:304'h0);
              inflight_opcodes <=(inflight_opcodes|(_GEN_0 ? _a_opcodes_set_T_1[1215:0]:1216'h0))&~(_GEN_23 ? _d_opcodes_clr_T_5[1215:0]:1216'h0);
              inflight_sizes <=(inflight_sizes|(_GEN_0 ? _a_sizes_set_T_1[1215:0]:1216'h0))&~(_GEN_23 ? _d_sizes_clr_T_5[1215:0]:1216'h0);
              a_first_counter_1 <=(~a_first_done|a_first_counter_1-1'h1)&a_first_counter_1;
              d_first_counter_1 <=(~d_first_done|d_first_counter_1-1'h1)&d_first_counter_1;
              if (a_first_done|d_first_done)
                 watchdog <=32'h0;
               else 
                 watchdog <=watchdog+32'h1;
            end 
         if (a_first_done&~a_first_counter)
            begin 
              opcode <=io_in_a_bits_opcode;
              param <=io_in_a_bits_param;
              size <=io_in_a_bits_size;
              source <=io_in_a_bits_source;
              address <=io_in_a_bits_address;
            end 
         if (d_first_done&~d_first_counter)
            begin 
              size_1 <=io_in_d_bits_size;
              source_1 <=io_in_d_bits_source;
            end 
       end
  
endmodule
 
module TLROM (
  input clock,
  input reset,
  output auto_in_a_ready,
  input auto_in_a_valid,
  input [2:0] auto_in_a_bits_opcode,
  input [2:0] auto_in_a_bits_param,
  input [1:0] auto_in_a_bits_size,
  input [8:0] auto_in_a_bits_source,
  input [16:0] auto_in_a_bits_address,
  input [7:0] auto_in_a_bits_mask,
  input auto_in_a_bits_corrupt,
  input auto_in_d_ready,
  output auto_in_d_valid,
  output [1:0] auto_in_d_bits_size,
  output [8:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data) ; 
   reg [63:0] casez_tmp ;  
  always @(*)
       begin 
         casez (auto_in_a_bits_address[11:3])
          9 'b000000000:
             casez_tmp =64'h10041B7C105073;
          9 'b000000001:
             casez_tmp =64'hF140257301F41413;
          9 'b000000010:
             casez_tmp =64'h705859300000597;
          9 'b000000011:
             casez_tmp =64'h8402;
          9 'b000000100:
             casez_tmp =64'h0;
          9 'b000000101:
             casez_tmp =64'h0;
          9 'b000000110:
             casez_tmp =64'h0;
          9 'b000000111:
             casez_tmp =64'h0;
          9 'b000001000:
             casez_tmp =64'hF14025737C105073;
          9 'b000001001:
             casez_tmp =64'h385859300000597;
          9 'b000001010:
             casez_tmp =64'h1050007330405073;
          9 'b000001011:
             casez_tmp =64'hBFF5;
          9 'b000001100:
             casez_tmp =64'h0;
          9 'b000001101:
             casez_tmp =64'h0;
          9 'b000001110:
             casez_tmp =64'h0;
          9 'b000001111:
             casez_tmp =64'h0;
          9 'b000010000:
             casez_tmp =64'h2090000EDFE0DD0;
          9 'b000010001:
             casez_tmp =64'h2807000038000000;
          9 'b000010010:
             casez_tmp =64'h1100000028000000;
          9 'b000010011:
             casez_tmp =64'h10000000;
          9 'b000010100:
             casez_tmp =64'hF0060000DA010000;
          9 'b000010101:
             casez_tmp =64'h0;
          9 'b000010110:
             casez_tmp =64'h0;
          9 'b000010111:
             casez_tmp =64'h1000000;
          9 'b000011000:
             casez_tmp =64'h400000003000000;
          9 'b000011001:
             casez_tmp =64'h100000000000000;
          9 'b000011010:
             casez_tmp =64'h400000003000000;
          9 'b000011011:
             casez_tmp =64'h10000000F000000;
          9 'b000011100:
             casez_tmp =64'h2100000003000000;
          9 'b000011101:
             casez_tmp =64'h656572661B000000;
          9 'b000011110:
             casez_tmp =64'h6F722C7370696863;
          9 'b000011111:
             casez_tmp =64'h7069686374656B63;
          9 'b000100000:
             casez_tmp =64'h6E776F6E6B6E752D;
          9 'b000100001:
             casez_tmp =64'h7665642D;
          9 'b000100010:
             casez_tmp =64'h1D00000003000000;
          9 'b000100011:
             casez_tmp =64'h6565726626000000;
          9 'b000100100:
             casez_tmp =64'h6F722C7370696863;
          9 'b000100101:
             casez_tmp =64'h7069686374656B63;
          9 'b000100110:
             casez_tmp =64'h6E776F6E6B6E752D;
          9 'b000100111:
             casez_tmp =64'h100000000000000;
          9 'b000101000:
             casez_tmp =64'h73757063;
          9 'b000101001:
             casez_tmp =64'h400000003000000;
          9 'b000101010:
             casez_tmp =64'h100000000000000;
          9 'b000101011:
             casez_tmp =64'h400000003000000;
          9 'b000101100:
             casez_tmp =64'hF000000;
          9 'b000101101:
             casez_tmp =64'h400000003000000;
          9 'b000101110:
             casez_tmp =64'h40420F002C000000;
          9 'b000101111:
             casez_tmp =64'h4075706301000000;
          9 'b000110000:
             casez_tmp =64'h300000000000030;
          9 'b000110001:
             casez_tmp =64'h3F00000004000000;
          9 'b000110010:
             casez_tmp =64'h300000000000000;
          9 'b000110011:
             casez_tmp =64'h1B00000015000000;
          9 'b000110100:
             casez_tmp =64'h722C657669666973;
          9 'b000110101:
             casez_tmp =64'h72003074656B636F;
          9 'b000110110:
             casez_tmp =64'h76637369;
          9 'b000110111:
             casez_tmp =64'h400000003000000;
          9 'b000111000:
             casez_tmp =64'h400000004F000000;
          9 'b000111001:
             casez_tmp =64'h400000003000000;
          9 'b000111010:
             casez_tmp =64'h4000000062000000;
          9 'b000111011:
             casez_tmp =64'h400000003000000;
          9 'b000111100:
             casez_tmp =64'h1000006F000000;
          9 'b000111101:
             casez_tmp =64'h400000003000000;
          9 'b000111110:
             casez_tmp =64'h7570637C000000;
          9 'b000111111:
             casez_tmp =64'h400000003000000;
          9 'b001000000:
             casez_tmp =64'h100000088000000;
          9 'b001000001:
             casez_tmp =64'h400000003000000;
          9 'b001000010:
             casez_tmp =64'h40000000A7000000;
          9 'b001000011:
             casez_tmp =64'h400000003000000;
          9 'b001000100:
             casez_tmp =64'h40000000BA000000;
          9 'b001000101:
             casez_tmp =64'h400000003000000;
          9 'b001000110:
             casez_tmp =64'h100000C7000000;
          9 'b001000111:
             casez_tmp =64'h400000003000000;
          9 'b001001000:
             casez_tmp =64'h1000000D4000000;
          9 'b001001001:
             casez_tmp =64'h400000003000000;
          9 'b001001010:
             casez_tmp =64'hE5000000;
          9 'b001001011:
             casez_tmp =64'h2500000003000000;
          9 'b001001100:
             casez_tmp =64'h34367672E9000000;
          9 'b001001101:
             casez_tmp =64'h7363697A63616D69;
          9 'b001001110:
             casez_tmp =64'h636E6566697A5F72;
          9 'b001001111:
             casez_tmp =64'h6D7068697A5F6965;
          9 'b001010000:
             casez_tmp =64'h74656B636F72785F;
          9 'b001010001:
             casez_tmp =64'h300000000000000;
          9 'b001010010:
             casez_tmp =64'hF300000004000000;
          9 'b001010011:
             casez_tmp =64'h300000004000000;
          9 'b001010100:
             casez_tmp =64'h801000004000000;
          9 'b001010101:
             casez_tmp =64'h300000008000000;
          9 'b001010110:
             casez_tmp =64'h1901000005000000;
          9 'b001010111:
             casez_tmp =64'h79616B6F;
          9 'b001011000:
             casez_tmp =64'h400000003000000;
          9 'b001011001:
             casez_tmp =64'h40420F002C000000;
          9 'b001011010:
             casez_tmp =64'h65746E6901000000;
          9 'b001011011:
             casez_tmp =64'h6F632D7470757272;
          9 'b001011100:
             casez_tmp =64'h72656C6C6F72746E;
          9 'b001011101:
             casez_tmp =64'h300000000000000;
          9 'b001011110:
             casez_tmp =64'h2001000004000000;
          9 'b001011111:
             casez_tmp =64'h300000001000000;
          9 'b001100000:
             casez_tmp =64'h1B0000000F000000;
          9 'b001100001:
             casez_tmp =64'h70632C7663736972;
          9 'b001100010:
             casez_tmp =64'h63746E692D75;
          9 'b001100011:
             casez_tmp =64'h3000000;
          9 'b001100100:
             casez_tmp =64'h300000031010000;
          9 'b001100101:
             casez_tmp =64'h4601000004000000;
          9 'b001100110:
             casez_tmp =64'h200000002000000;
          9 'b001100111:
             casez_tmp =64'h200000002000000;
          9 'b001101000:
             casez_tmp =64'h6F6D656D01000000;
          9 'b001101001:
             casez_tmp =64'h3030303038407972;
          9 'b001101010:
             casez_tmp =64'h300000000303030;
          9 'b001101011:
             casez_tmp =64'h7C00000007000000;
          9 'b001101100:
             casez_tmp =64'h79726F6D656D;
          9 'b001101101:
             casez_tmp =64'h800000003000000;
          9 'b001101110:
             casez_tmp =64'h80E5000000;
          9 'b001101111:
             casez_tmp =64'h300000000000010;
          9 'b001110000:
             casez_tmp =64'h4601000004000000;
          9 'b001110001:
             casez_tmp =64'h200000001000000;
          9 'b001110010:
             casez_tmp =64'h636F7301000000;
          9 'b001110011:
             casez_tmp =64'h400000003000000;
          9 'b001110100:
             casez_tmp =64'h100000000000000;
          9 'b001110101:
             casez_tmp =64'h400000003000000;
          9 'b001110110:
             casez_tmp =64'h10000000F000000;
          9 'b001110111:
             casez_tmp =64'h2C00000003000000;
          9 'b001111000:
             casez_tmp =64'h656572661B000000;
          9 'b001111001:
             casez_tmp =64'h6F722C7370696863;
          9 'b001111010:
             casez_tmp =64'h7069686374656B63;
          9 'b001111011:
             casez_tmp =64'h6E776F6E6B6E752D;
          9 'b001111100:
             casez_tmp =64'h6D697300636F732D;
          9 'b001111101:
             casez_tmp =64'h7375622D656C70;
          9 'b001111110:
             casez_tmp =64'h3000000;
          9 'b001111111:
             casez_tmp =64'h10000004E010000;
          9 'b010000000:
             casez_tmp =64'h303240746E696C63;
          9 'b010000001:
             casez_tmp =64'h3030303030;
          9 'b010000010:
             casez_tmp =64'hD00000003000000;
          9 'b010000011:
             casez_tmp =64'h637369721B000000;
          9 'b010000100:
             casez_tmp =64'h30746E696C632C76;
          9 'b010000101:
             casez_tmp =64'h300000000000000;
          9 'b010000110:
             casez_tmp =64'h5501000010000000;
          9 'b010000111:
             casez_tmp =64'h300000002000000;
          9 'b010001000:
             casez_tmp =64'h700000002000000;
          9 'b010001001:
             casez_tmp =64'h800000003000000;
          9 'b010001010:
             casez_tmp =64'h2E5000000;
          9 'b010001011:
             casez_tmp =64'h300000000000100;
          9 'b010001100:
             casez_tmp =64'h6901000008000000;
          9 'b010001101:
             casez_tmp =64'h6C6F72746E6F63;
          9 'b010001110:
             casez_tmp =64'h100000002000000;
          9 'b010001111:
             casez_tmp =64'h6F632D6775626564;
          9 'b010010000:
             casez_tmp =64'h72656C6C6F72746E;
          9 'b010010001:
             casez_tmp =64'h300000000003040;
          9 'b010010010:
             casez_tmp =64'h1B00000021000000;
          9 'b010010011:
             casez_tmp =64'h642C657669666973;
          9 'b010010100:
             casez_tmp =64'h3331302D67756265;
          9 'b010010101:
             casez_tmp =64'h642C766373697200;
          9 'b010010110:
             casez_tmp =64'h3331302D67756265;
          9 'b010010111:
             casez_tmp =64'h300000000000000;
          9 'b010011000:
             casez_tmp =64'h7301000004000000;
          9 'b010011001:
             casez_tmp =64'h300000000696D64;
          9 'b010011010:
             casez_tmp =64'h5501000008000000;
          9 'b010011011:
             casez_tmp =64'hFFFF000002000000;
          9 'b010011100:
             casez_tmp =64'h800000003000000;
          9 'b010011101:
             casez_tmp =64'hE5000000;
          9 'b010011110:
             casez_tmp =64'h300000000100000;
          9 'b010011111:
             casez_tmp =64'h6901000008000000;
          9 'b010100000:
             casez_tmp =64'h6C6F72746E6F63;
          9 'b010100001:
             casez_tmp =64'h100000002000000;
          9 'b010100010:
             casez_tmp =64'h65642D726F727265;
          9 'b010100011:
             casez_tmp =64'h3030334065636976;
          9 'b010100100:
             casez_tmp =64'h300000000000030;
          9 'b010100101:
             casez_tmp =64'h1B0000000E000000;
          9 'b010100110:
             casez_tmp =64'h652C657669666973;
          9 'b010100111:
             casez_tmp =64'h30726F7272;
          9 'b010101000:
             casez_tmp =64'h800000003000000;
          9 'b010101001:
             casez_tmp =64'h300000E5000000;
          9 'b010101010:
             casez_tmp =64'h200000000100000;
          9 'b010101011:
             casez_tmp =64'h6574786501000000;
          9 'b010101100:
             casez_tmp =64'h746E692D6C616E72;
          9 'b010101101:
             casez_tmp =64'h73747075727265;
          9 'b010101110:
             casez_tmp =64'h400000003000000;
          9 'b010101111:
             casez_tmp =64'h300000080010000;
          9 'b010110000:
             casez_tmp =64'h800000003000000;
          9 'b010110001:
             casez_tmp =64'h100000091010000;
          9 'b010110010:
             casez_tmp =64'h200000002000000;
          9 'b010110011:
             casez_tmp =64'h65746E6901000000;
          9 'b010110100:
             casez_tmp =64'h6F632D7470757272;
          9 'b010110101:
             casez_tmp =64'h72656C6C6F72746E;
          9 'b010110110:
             casez_tmp =64'h3030303030306340;
          9 'b010110111:
             casez_tmp =64'h300000000000000;
          9 'b010111000:
             casez_tmp =64'h2001000004000000;
          9 'b010111001:
             casez_tmp =64'h300000001000000;
          9 'b010111010:
             casez_tmp =64'h1B0000000C000000;
          9 'b010111011:
             casez_tmp =64'h6C702C7663736972;
          9 'b010111100:
             casez_tmp =64'h300000000306369;
          9 'b010111101:
             casez_tmp =64'h3101000000000000;
          9 'b010111110:
             casez_tmp =64'h800000003000000;
          9 'b010111111:
             casez_tmp =64'h200000055010000;
          9 'b011000000:
             casez_tmp =64'h30000000B000000;
          9 'b011000001:
             casez_tmp =64'hE500000008000000;
          9 'b011000010:
             casez_tmp =64'h40000000C;
          9 'b011000011:
             casez_tmp =64'h800000003000000;
          9 'b011000100:
             casez_tmp =64'h746E6F6369010000;
          9 'b011000101:
             casez_tmp =64'h3000000006C6F72;
          9 'b011000110:
             casez_tmp =64'h9C01000004000000;
          9 'b011000111:
             casez_tmp =64'h300000003000000;
          9 'b011001000:
             casez_tmp =64'hAF01000004000000;
          9 'b011001001:
             casez_tmp =64'h300000002000000;
          9 'b011001010:
             casez_tmp =64'h4601000004000000;
          9 'b011001011:
             casez_tmp =64'h200000003000000;
          9 'b011001100:
             casez_tmp =64'h6F696D6D01000000;
          9 'b011001101:
             casez_tmp =64'h78612D74726F702D;
          9 'b011001110:
             casez_tmp =64'h3030303036403469;
          9 'b011001111:
             casez_tmp =64'h300000000303030;
          9 'b011010000:
             casez_tmp =64'h4000000;
          9 'b011010001:
             casez_tmp =64'h300000001000000;
          9 'b011010010:
             casez_tmp =64'hF00000004000000;
          9 'b011010011:
             casez_tmp =64'h300000001000000;
          9 'b011010100:
             casez_tmp =64'h1B0000000B000000;
          9 'b011010101:
             casez_tmp =64'h622D656C706D6973;
          9 'b011010110:
             casez_tmp =64'h300000000007375;
          9 'b011010111:
             casez_tmp =64'h4E0100000C000000;
          9 'b011011000:
             casez_tmp =64'h6000000060;
          9 'b011011001:
             casez_tmp =64'h200000000000020;
          9 'b011011010:
             casez_tmp =64'h406D6F7201000000;
          9 'b011011011:
             casez_tmp =64'h3030303031;
          9 'b011011100:
             casez_tmp =64'hC00000003000000;
          9 'b011011101:
             casez_tmp =64'h696669731B000000;
          9 'b011011110:
             casez_tmp =64'h306D6F722C6576;
          9 'b011011111:
             casez_tmp =64'h800000003000000;
          9 'b011100000:
             casez_tmp =64'h100E5000000;
          9 'b011100001:
             casez_tmp =64'h300000000000100;
          9 'b011100010:
             casez_tmp =64'h6901000004000000;
          9 'b011100011:
             casez_tmp =64'h2000000006D656D;
          9 'b011100100:
             casez_tmp =64'h7362757301000000;
          9 'b011100101:
             casez_tmp =64'h62705F6D65747379;
          9 'b011100110:
             casez_tmp =64'h6B636F6C635F7375;
          9 'b011100111:
             casez_tmp =64'h300000000000000;
          9 'b011101000:
             casez_tmp =64'hBA01000004000000;
          9 'b011101001:
             casez_tmp =64'h300000000000000;
          9 'b011101010:
             casez_tmp =64'h3F00000004000000;
          9 'b011101011:
             casez_tmp =64'h300000000E1F505;
          9 'b011101100:
             casez_tmp =64'hC701000015000000;
          9 'b011101101:
             casez_tmp =64'h6574737973627573;
          9 'b011101110:
             casez_tmp =64'h635F737562705F6D;
          9 'b011101111:
             casez_tmp =64'h6B636F6C;
          9 'b011110000:
             casez_tmp =64'hC00000003000000;
          9 'b011110001:
             casez_tmp =64'h657869661B000000;
          9 'b011110010:
             casez_tmp =64'h6B636F6C632D64;
          9 'b011110011:
             casez_tmp =64'h200000002000000;
          9 'b011110100:
             casez_tmp =64'h900000002000000;
          9 'b011110101:
             casez_tmp =64'h7373657264646123;
          9 'b011110110:
             casez_tmp =64'h2300736C6C65632D;
          9 'b011110111:
             casez_tmp =64'h6C65632D657A6973;
          9 'b011111000:
             casez_tmp =64'h61706D6F6300736C;
          9 'b011111001:
             casez_tmp =64'h6F6D00656C626974;
          9 'b011111010:
             casez_tmp =64'h656D6974006C6564;
          9 'b011111011:
             casez_tmp =64'h6572662D65736162;
          9 'b011111100:
             casez_tmp =64'h630079636E657571;
          9 'b011111101:
             casez_tmp =64'h6572662D6B636F6C;
          9 'b011111110:
             casez_tmp =64'h640079636E657571;
          9 'b011111111:
             casez_tmp =64'h622D65686361632D;
          9 'b100000000:
             casez_tmp =64'h7A69732D6B636F6C;
          9 'b100000001:
             casez_tmp =64'h686361632D640065;
          9 'b100000010:
             casez_tmp =64'h6400737465732D65;
          9 'b100000011:
             casez_tmp =64'h732D65686361632D;
          9 'b100000100:
             casez_tmp =64'h6976656400657A69;
          9 'b100000101:
             casez_tmp =64'h657079745F6563;
          9 'b100000110:
             casez_tmp =64'h6572617764726168;
          9 'b100000111:
             casez_tmp =64'h72622D636578652D;
          9 'b100001000:
             casez_tmp =64'h746E696F706B6165;
          9 'b100001001:
             casez_tmp =64'h6900746E756F632D;
          9 'b100001010:
             casez_tmp =64'h622D65686361632D;
          9 'b100001011:
             casez_tmp =64'h7A69732D6B636F6C;
          9 'b100001100:
             casez_tmp =64'h686361632D690065;
          9 'b100001101:
             casez_tmp =64'h6900737465732D65;
          9 'b100001110:
             casez_tmp =64'h732D65686361632D;
          9 'b100001111:
             casez_tmp =64'h7478656E00657A69;
          9 'b100010000:
             casez_tmp =64'h632D6C6576656C2D;
          9 'b100010001:
             casez_tmp =64'h6765720065686361;
          9 'b100010010:
             casez_tmp =64'h692C766373697200;
          9 'b100010011:
             casez_tmp =64'h7663736972006173;
          9 'b100010100:
             casez_tmp =64'h6E617267706D702C;
          9 'b100010101:
             casez_tmp =64'h79746972616C75;
          9 'b100010110:
             casez_tmp =64'h6D702C7663736972;
          9 'b100010111:
             casez_tmp =64'h736E6F6967657270;
          9 'b100011000:
             casez_tmp =64'h73757461747300;
          9 'b100011001:
             casez_tmp =64'h75727265746E6923;
          9 'b100011010:
             casez_tmp =64'h736C6C65632D7470;
          9 'b100011011:
             casez_tmp =64'h75727265746E6900;
          9 'b100011100:
             casez_tmp =64'h72746E6F632D7470;
          9 'b100011101:
             casez_tmp =64'h68700072656C6C6F;
          9 'b100011110:
             casez_tmp =64'h617200656C646E61;
          9 'b100011111:
             casez_tmp =64'h746E69007365676E;
          9 'b100100000:
             casez_tmp =64'h2D73747075727265;
          9 'b100100001:
             casez_tmp =64'h6465646E65747865;
          9 'b100100010:
             casez_tmp =64'h6D616E2D67657200;
          9 'b100100011:
             casez_tmp =64'h6775626564007365;
          9 'b100100100:
             casez_tmp =64'h6863617474612D;
          9 'b100100101:
             casez_tmp =64'h7075727265746E69;
          9 'b100100110:
             casez_tmp =64'h746E657261702D74;
          9 'b100100111:
             casez_tmp =64'h75727265746E6900;
          9 'b100101000:
             casez_tmp =64'h6373697200737470;
          9 'b100101001:
             casez_tmp =64'h72702D78616D2C76;
          9 'b100101010:
             casez_tmp =64'h7200797469726F69;
          9 'b100101011:
             casez_tmp =64'h65646E2C76637369;
          9 'b100101100:
             casez_tmp =64'h6B636F6C63230076;
          9 'b100101101:
             casez_tmp =64'h6300736C6C65632D;
          9 'b100101110:
             casez_tmp =64'h74756F2D6B636F6C;
          9 'b100101111:
             casez_tmp =64'h656D616E2D747570;
          9 'b100110000:
             casez_tmp =64'h73;
          9 'b100110001:
             casez_tmp =64'h0;
          9 'b100110010:
             casez_tmp =64'h0;
          9 'b100110011:
             casez_tmp =64'h0;
          9 'b100110100:
             casez_tmp =64'h0;
          9 'b100110101:
             casez_tmp =64'h0;
          9 'b100110110:
             casez_tmp =64'h0;
          9 'b100110111:
             casez_tmp =64'h0;
          9 'b100111000:
             casez_tmp =64'h0;
          9 'b100111001:
             casez_tmp =64'h0;
          9 'b100111010:
             casez_tmp =64'h0;
          9 'b100111011:
             casez_tmp =64'h0;
          9 'b100111100:
             casez_tmp =64'h0;
          9 'b100111101:
             casez_tmp =64'h0;
          9 'b100111110:
             casez_tmp =64'h0;
          9 'b100111111:
             casez_tmp =64'h0;
          9 'b101000000:
             casez_tmp =64'h0;
          9 'b101000001:
             casez_tmp =64'h0;
          9 'b101000010:
             casez_tmp =64'h0;
          9 'b101000011:
             casez_tmp =64'h0;
          9 'b101000100:
             casez_tmp =64'h0;
          9 'b101000101:
             casez_tmp =64'h0;
          9 'b101000110:
             casez_tmp =64'h0;
          9 'b101000111:
             casez_tmp =64'h0;
          9 'b101001000:
             casez_tmp =64'h0;
          9 'b101001001:
             casez_tmp =64'h0;
          9 'b101001010:
             casez_tmp =64'h0;
          9 'b101001011:
             casez_tmp =64'h0;
          9 'b101001100:
             casez_tmp =64'h0;
          9 'b101001101:
             casez_tmp =64'h0;
          9 'b101001110:
             casez_tmp =64'h0;
          9 'b101001111:
             casez_tmp =64'h0;
          9 'b101010000:
             casez_tmp =64'h0;
          9 'b101010001:
             casez_tmp =64'h0;
          9 'b101010010:
             casez_tmp =64'h0;
          9 'b101010011:
             casez_tmp =64'h0;
          9 'b101010100:
             casez_tmp =64'h0;
          9 'b101010101:
             casez_tmp =64'h0;
          9 'b101010110:
             casez_tmp =64'h0;
          9 'b101010111:
             casez_tmp =64'h0;
          9 'b101011000:
             casez_tmp =64'h0;
          9 'b101011001:
             casez_tmp =64'h0;
          9 'b101011010:
             casez_tmp =64'h0;
          9 'b101011011:
             casez_tmp =64'h0;
          9 'b101011100:
             casez_tmp =64'h0;
          9 'b101011101:
             casez_tmp =64'h0;
          9 'b101011110:
             casez_tmp =64'h0;
          9 'b101011111:
             casez_tmp =64'h0;
          9 'b101100000:
             casez_tmp =64'h0;
          9 'b101100001:
             casez_tmp =64'h0;
          9 'b101100010:
             casez_tmp =64'h0;
          9 'b101100011:
             casez_tmp =64'h0;
          9 'b101100100:
             casez_tmp =64'h0;
          9 'b101100101:
             casez_tmp =64'h0;
          9 'b101100110:
             casez_tmp =64'h0;
          9 'b101100111:
             casez_tmp =64'h0;
          9 'b101101000:
             casez_tmp =64'h0;
          9 'b101101001:
             casez_tmp =64'h0;
          9 'b101101010:
             casez_tmp =64'h0;
          9 'b101101011:
             casez_tmp =64'h0;
          9 'b101101100:
             casez_tmp =64'h0;
          9 'b101101101:
             casez_tmp =64'h0;
          9 'b101101110:
             casez_tmp =64'h0;
          9 'b101101111:
             casez_tmp =64'h0;
          9 'b101110000:
             casez_tmp =64'h0;
          9 'b101110001:
             casez_tmp =64'h0;
          9 'b101110010:
             casez_tmp =64'h0;
          9 'b101110011:
             casez_tmp =64'h0;
          9 'b101110100:
             casez_tmp =64'h0;
          9 'b101110101:
             casez_tmp =64'h0;
          9 'b101110110:
             casez_tmp =64'h0;
          9 'b101110111:
             casez_tmp =64'h0;
          9 'b101111000:
             casez_tmp =64'h0;
          9 'b101111001:
             casez_tmp =64'h0;
          9 'b101111010:
             casez_tmp =64'h0;
          9 'b101111011:
             casez_tmp =64'h0;
          9 'b101111100:
             casez_tmp =64'h0;
          9 'b101111101:
             casez_tmp =64'h0;
          9 'b101111110:
             casez_tmp =64'h0;
          9 'b101111111:
             casez_tmp =64'h0;
          9 'b110000000:
             casez_tmp =64'h0;
          9 'b110000001:
             casez_tmp =64'h0;
          9 'b110000010:
             casez_tmp =64'h0;
          9 'b110000011:
             casez_tmp =64'h0;
          9 'b110000100:
             casez_tmp =64'h0;
          9 'b110000101:
             casez_tmp =64'h0;
          9 'b110000110:
             casez_tmp =64'h0;
          9 'b110000111:
             casez_tmp =64'h0;
          9 'b110001000:
             casez_tmp =64'h0;
          9 'b110001001:
             casez_tmp =64'h0;
          9 'b110001010:
             casez_tmp =64'h0;
          9 'b110001011:
             casez_tmp =64'h0;
          9 'b110001100:
             casez_tmp =64'h0;
          9 'b110001101:
             casez_tmp =64'h0;
          9 'b110001110:
             casez_tmp =64'h0;
          9 'b110001111:
             casez_tmp =64'h0;
          9 'b110010000:
             casez_tmp =64'h0;
          9 'b110010001:
             casez_tmp =64'h0;
          9 'b110010010:
             casez_tmp =64'h0;
          9 'b110010011:
             casez_tmp =64'h0;
          9 'b110010100:
             casez_tmp =64'h0;
          9 'b110010101:
             casez_tmp =64'h0;
          9 'b110010110:
             casez_tmp =64'h0;
          9 'b110010111:
             casez_tmp =64'h0;
          9 'b110011000:
             casez_tmp =64'h0;
          9 'b110011001:
             casez_tmp =64'h0;
          9 'b110011010:
             casez_tmp =64'h0;
          9 'b110011011:
             casez_tmp =64'h0;
          9 'b110011100:
             casez_tmp =64'h0;
          9 'b110011101:
             casez_tmp =64'h0;
          9 'b110011110:
             casez_tmp =64'h0;
          9 'b110011111:
             casez_tmp =64'h0;
          9 'b110100000:
             casez_tmp =64'h0;
          9 'b110100001:
             casez_tmp =64'h0;
          9 'b110100010:
             casez_tmp =64'h0;
          9 'b110100011:
             casez_tmp =64'h0;
          9 'b110100100:
             casez_tmp =64'h0;
          9 'b110100101:
             casez_tmp =64'h0;
          9 'b110100110:
             casez_tmp =64'h0;
          9 'b110100111:
             casez_tmp =64'h0;
          9 'b110101000:
             casez_tmp =64'h0;
          9 'b110101001:
             casez_tmp =64'h0;
          9 'b110101010:
             casez_tmp =64'h0;
          9 'b110101011:
             casez_tmp =64'h0;
          9 'b110101100:
             casez_tmp =64'h0;
          9 'b110101101:
             casez_tmp =64'h0;
          9 'b110101110:
             casez_tmp =64'h0;
          9 'b110101111:
             casez_tmp =64'h0;
          9 'b110110000:
             casez_tmp =64'h0;
          9 'b110110001:
             casez_tmp =64'h0;
          9 'b110110010:
             casez_tmp =64'h0;
          9 'b110110011:
             casez_tmp =64'h0;
          9 'b110110100:
             casez_tmp =64'h0;
          9 'b110110101:
             casez_tmp =64'h0;
          9 'b110110110:
             casez_tmp =64'h0;
          9 'b110110111:
             casez_tmp =64'h0;
          9 'b110111000:
             casez_tmp =64'h0;
          9 'b110111001:
             casez_tmp =64'h0;
          9 'b110111010:
             casez_tmp =64'h0;
          9 'b110111011:
             casez_tmp =64'h0;
          9 'b110111100:
             casez_tmp =64'h0;
          9 'b110111101:
             casez_tmp =64'h0;
          9 'b110111110:
             casez_tmp =64'h0;
          9 'b110111111:
             casez_tmp =64'h0;
          9 'b111000000:
             casez_tmp =64'h0;
          9 'b111000001:
             casez_tmp =64'h0;
          9 'b111000010:
             casez_tmp =64'h0;
          9 'b111000011:
             casez_tmp =64'h0;
          9 'b111000100:
             casez_tmp =64'h0;
          9 'b111000101:
             casez_tmp =64'h0;
          9 'b111000110:
             casez_tmp =64'h0;
          9 'b111000111:
             casez_tmp =64'h0;
          9 'b111001000:
             casez_tmp =64'h0;
          9 'b111001001:
             casez_tmp =64'h0;
          9 'b111001010:
             casez_tmp =64'h0;
          9 'b111001011:
             casez_tmp =64'h0;
          9 'b111001100:
             casez_tmp =64'h0;
          9 'b111001101:
             casez_tmp =64'h0;
          9 'b111001110:
             casez_tmp =64'h0;
          9 'b111001111:
             casez_tmp =64'h0;
          9 'b111010000:
             casez_tmp =64'h0;
          9 'b111010001:
             casez_tmp =64'h0;
          9 'b111010010:
             casez_tmp =64'h0;
          9 'b111010011:
             casez_tmp =64'h0;
          9 'b111010100:
             casez_tmp =64'h0;
          9 'b111010101:
             casez_tmp =64'h0;
          9 'b111010110:
             casez_tmp =64'h0;
          9 'b111010111:
             casez_tmp =64'h0;
          9 'b111011000:
             casez_tmp =64'h0;
          9 'b111011001:
             casez_tmp =64'h0;
          9 'b111011010:
             casez_tmp =64'h0;
          9 'b111011011:
             casez_tmp =64'h0;
          9 'b111011100:
             casez_tmp =64'h0;
          9 'b111011101:
             casez_tmp =64'h0;
          9 'b111011110:
             casez_tmp =64'h0;
          9 'b111011111:
             casez_tmp =64'h0;
          9 'b111100000:
             casez_tmp =64'h0;
          9 'b111100001:
             casez_tmp =64'h0;
          9 'b111100010:
             casez_tmp =64'h0;
          9 'b111100011:
             casez_tmp =64'h0;
          9 'b111100100:
             casez_tmp =64'h0;
          9 'b111100101:
             casez_tmp =64'h0;
          9 'b111100110:
             casez_tmp =64'h0;
          9 'b111100111:
             casez_tmp =64'h0;
          9 'b111101000:
             casez_tmp =64'h0;
          9 'b111101001:
             casez_tmp =64'h0;
          9 'b111101010:
             casez_tmp =64'h0;
          9 'b111101011:
             casez_tmp =64'h0;
          9 'b111101100:
             casez_tmp =64'h0;
          9 'b111101101:
             casez_tmp =64'h0;
          9 'b111101110:
             casez_tmp =64'h0;
          9 'b111101111:
             casez_tmp =64'h0;
          9 'b111110000:
             casez_tmp =64'h0;
          9 'b111110001:
             casez_tmp =64'h0;
          9 'b111110010:
             casez_tmp =64'h0;
          9 'b111110011:
             casez_tmp =64'h0;
          9 'b111110100:
             casez_tmp =64'h0;
          9 'b111110101:
             casez_tmp =64'h0;
          9 'b111110110:
             casez_tmp =64'h0;
          9 'b111110111:
             casez_tmp =64'h0;
          9 'b111111000:
             casez_tmp =64'h0;
          9 'b111111001:
             casez_tmp =64'h0;
          9 'b111111010:
             casez_tmp =64'h0;
          9 'b111111011:
             casez_tmp =64'h0;
          9 'b111111100:
             casez_tmp =64'h0;
          9 'b111111101:
             casez_tmp =64'h0;
          9 'b111111110:
             casez_tmp =64'h0;
          default :
             casez_tmp =64'h0;
         endcase 
       end
  
  TLMonitor_35 monitor(.clock(clock),.reset(reset),.io_in_a_ready(auto_in_d_ready),.io_in_a_valid(auto_in_a_valid),.io_in_a_bits_opcode(auto_in_a_bits_opcode),.io_in_a_bits_param(auto_in_a_bits_param),.io_in_a_bits_size(auto_in_a_bits_size),.io_in_a_bits_source(auto_in_a_bits_source),.io_in_a_bits_address(auto_in_a_bits_address),.io_in_a_bits_mask(auto_in_a_bits_mask),.io_in_a_bits_corrupt(auto_in_a_bits_corrupt),.io_in_d_ready(auto_in_d_ready),.io_in_d_valid(auto_in_a_valid),.io_in_d_bits_size(auto_in_a_bits_size),.io_in_d_bits_source(auto_in_a_bits_source)); 
  assign auto_in_a_ready=auto_in_d_ready; 
  assign auto_in_d_valid=auto_in_a_valid; 
  assign auto_in_d_bits_size=auto_in_a_bits_size; 
  assign auto_in_d_bits_source=auto_in_a_bits_source; 
  assign auto_in_d_bits_data=(|(auto_in_a_bits_address[15:12])) ? 64'h0:casez_tmp; 
endmodule
 
module ClockSinkDomain_1 (
  output auto_bootrom_in_a_ready,
  input auto_bootrom_in_a_valid,
  input [2:0] auto_bootrom_in_a_bits_opcode,
  input [2:0] auto_bootrom_in_a_bits_param,
  input [1:0] auto_bootrom_in_a_bits_size,
  input [8:0] auto_bootrom_in_a_bits_source,
  input [16:0] auto_bootrom_in_a_bits_address,
  input [7:0] auto_bootrom_in_a_bits_mask,
  input auto_bootrom_in_a_bits_corrupt,
  input auto_bootrom_in_d_ready,
  output auto_bootrom_in_d_valid,
  output [1:0] auto_bootrom_in_d_bits_size,
  output [8:0] auto_bootrom_in_d_bits_source,
  output [63:0] auto_bootrom_in_d_bits_data,
  input auto_clock_in_clock,
  input auto_clock_in_reset) ; 
  TLROM bootrom(.clock(auto_clock_in_clock),.reset(auto_clock_in_reset),.auto_in_a_ready(auto_bootrom_in_a_ready),.auto_in_a_valid(auto_bootrom_in_a_valid),.auto_in_a_bits_opcode(auto_bootrom_in_a_bits_opcode),.auto_in_a_bits_param(auto_bootrom_in_a_bits_param),.auto_in_a_bits_size(auto_bootrom_in_a_bits_size),.auto_in_a_bits_source(auto_bootrom_in_a_bits_source),.auto_in_a_bits_address(auto_bootrom_in_a_bits_address),.auto_in_a_bits_mask(auto_bootrom_in_a_bits_mask),.auto_in_a_bits_corrupt(auto_bootrom_in_a_bits_corrupt),.auto_in_d_ready(auto_bootrom_in_d_ready),.auto_in_d_valid(auto_bootrom_in_d_valid),.auto_in_d_bits_size(auto_bootrom_in_d_bits_size),.auto_in_d_bits_source(auto_bootrom_in_d_bits_source),.auto_in_d_bits_data(auto_bootrom_in_d_bits_data)); 
endmodule
 
module ExampleRocketSystem (
  input clock,
  input reset,
  input resetctrl_hartIsInReset_0,
  input debug_clock,
  input debug_reset,
  output debug_clockeddmi_dmi_req_ready,
  input debug_clockeddmi_dmi_req_valid,
  input [6:0] debug_clockeddmi_dmi_req_bits_addr,
  input [31:0] debug_clockeddmi_dmi_req_bits_data,
  input [1:0] debug_clockeddmi_dmi_req_bits_op,
  input debug_clockeddmi_dmi_resp_ready,
  output debug_clockeddmi_dmi_resp_valid,
  output [31:0] debug_clockeddmi_dmi_resp_bits_data,
  output [1:0] debug_clockeddmi_dmi_resp_bits_resp,
  input debug_clockeddmi_dmiClock,
  input debug_clockeddmi_dmiReset,
  output debug_ndreset,
  output debug_dmactive,
  input debug_dmactiveAck,
  input mem_axi4_0_aw_ready,
  output mem_axi4_0_aw_valid,
  output [3:0] mem_axi4_0_aw_bits_id,
  output [31:0] mem_axi4_0_aw_bits_addr,
  output [7:0] mem_axi4_0_aw_bits_len,
  output [2:0] mem_axi4_0_aw_bits_size,
  output [1:0] mem_axi4_0_aw_bits_burst,
  output mem_axi4_0_aw_bits_lock,
  output [3:0] mem_axi4_0_aw_bits_cache,
  output [2:0] mem_axi4_0_aw_bits_prot,
  output [3:0] mem_axi4_0_aw_bits_qos,
  input mem_axi4_0_w_ready,
  output mem_axi4_0_w_valid,
  output [63:0] mem_axi4_0_w_bits_data,
  output [7:0] mem_axi4_0_w_bits_strb,
  output mem_axi4_0_w_bits_last,
  output mem_axi4_0_b_ready,
  input mem_axi4_0_b_valid,
  input [3:0] mem_axi4_0_b_bits_id,
  input [1:0] mem_axi4_0_b_bits_resp,
  input mem_axi4_0_ar_ready,
  output mem_axi4_0_ar_valid,
  output [3:0] mem_axi4_0_ar_bits_id,
  output [31:0] mem_axi4_0_ar_bits_addr,
  output [7:0] mem_axi4_0_ar_bits_len,
  output [2:0] mem_axi4_0_ar_bits_size,
  output [1:0] mem_axi4_0_ar_bits_burst,
  output mem_axi4_0_ar_bits_lock,
  output [3:0] mem_axi4_0_ar_bits_cache,
  output [2:0] mem_axi4_0_ar_bits_prot,
  output [3:0] mem_axi4_0_ar_bits_qos,
  output mem_axi4_0_r_ready,
  input mem_axi4_0_r_valid,
  input [3:0] mem_axi4_0_r_bits_id,
  input [63:0] mem_axi4_0_r_bits_data,
  input [1:0] mem_axi4_0_r_bits_resp,
  input mem_axi4_0_r_bits_last,
  input mmio_axi4_0_aw_ready,
  output mmio_axi4_0_aw_valid,
  output [3:0] mmio_axi4_0_aw_bits_id,
  output [30:0] mmio_axi4_0_aw_bits_addr,
  output [7:0] mmio_axi4_0_aw_bits_len,
  output [2:0] mmio_axi4_0_aw_bits_size,
  output [1:0] mmio_axi4_0_aw_bits_burst,
  output mmio_axi4_0_aw_bits_lock,
  output [3:0] mmio_axi4_0_aw_bits_cache,
  output [2:0] mmio_axi4_0_aw_bits_prot,
  output [3:0] mmio_axi4_0_aw_bits_qos,
  input mmio_axi4_0_w_ready,
  output mmio_axi4_0_w_valid,
  output [63:0] mmio_axi4_0_w_bits_data,
  output [7:0] mmio_axi4_0_w_bits_strb,
  output mmio_axi4_0_w_bits_last,
  output mmio_axi4_0_b_ready,
  input mmio_axi4_0_b_valid,
  input [3:0] mmio_axi4_0_b_bits_id,
  input [1:0] mmio_axi4_0_b_bits_resp,
  input mmio_axi4_0_ar_ready,
  output mmio_axi4_0_ar_valid,
  output [3:0] mmio_axi4_0_ar_bits_id,
  output [30:0] mmio_axi4_0_ar_bits_addr,
  output [7:0] mmio_axi4_0_ar_bits_len,
  output [2:0] mmio_axi4_0_ar_bits_size,
  output [1:0] mmio_axi4_0_ar_bits_burst,
  output mmio_axi4_0_ar_bits_lock,
  output [3:0] mmio_axi4_0_ar_bits_cache,
  output [2:0] mmio_axi4_0_ar_bits_prot,
  output [3:0] mmio_axi4_0_ar_bits_qos,
  output mmio_axi4_0_r_ready,
  input mmio_axi4_0_r_valid,
  input [3:0] mmio_axi4_0_r_bits_id,
  input [63:0] mmio_axi4_0_r_bits_data,
  input [1:0] mmio_axi4_0_r_bits_resp,
  input mmio_axi4_0_r_bits_last,
  output l2_frontend_bus_axi4_0_aw_ready,
  input l2_frontend_bus_axi4_0_aw_valid,
  input [7:0] l2_frontend_bus_axi4_0_aw_bits_id,
  input [31:0] l2_frontend_bus_axi4_0_aw_bits_addr,
  input [7:0] l2_frontend_bus_axi4_0_aw_bits_len,
  input [2:0] l2_frontend_bus_axi4_0_aw_bits_size,
  input [1:0] l2_frontend_bus_axi4_0_aw_bits_burst,
  input l2_frontend_bus_axi4_0_aw_bits_lock,
  input [3:0] l2_frontend_bus_axi4_0_aw_bits_cache,
  input [2:0] l2_frontend_bus_axi4_0_aw_bits_prot,
  input [3:0] l2_frontend_bus_axi4_0_aw_bits_qos,
  output l2_frontend_bus_axi4_0_w_ready,
  input l2_frontend_bus_axi4_0_w_valid,
  input [63:0] l2_frontend_bus_axi4_0_w_bits_data,
  input [7:0] l2_frontend_bus_axi4_0_w_bits_strb,
  input l2_frontend_bus_axi4_0_w_bits_last,
  input l2_frontend_bus_axi4_0_b_ready,
  output l2_frontend_bus_axi4_0_b_valid,
  output [7:0] l2_frontend_bus_axi4_0_b_bits_id,
  output [1:0] l2_frontend_bus_axi4_0_b_bits_resp,
  output l2_frontend_bus_axi4_0_ar_ready,
  input l2_frontend_bus_axi4_0_ar_valid,
  input [7:0] l2_frontend_bus_axi4_0_ar_bits_id,
  input [31:0] l2_frontend_bus_axi4_0_ar_bits_addr,
  input [7:0] l2_frontend_bus_axi4_0_ar_bits_len,
  input [2:0] l2_frontend_bus_axi4_0_ar_bits_size,
  input [1:0] l2_frontend_bus_axi4_0_ar_bits_burst,
  input l2_frontend_bus_axi4_0_ar_bits_lock,
  input [3:0] l2_frontend_bus_axi4_0_ar_bits_cache,
  input [2:0] l2_frontend_bus_axi4_0_ar_bits_prot,
  input [3:0] l2_frontend_bus_axi4_0_ar_bits_qos,
  input l2_frontend_bus_axi4_0_r_ready,
  output l2_frontend_bus_axi4_0_r_valid,
  output [7:0] l2_frontend_bus_axi4_0_r_bits_id,
  output [63:0] l2_frontend_bus_axi4_0_r_bits_data,
  output [1:0] l2_frontend_bus_axi4_0_r_bits_resp,
  output l2_frontend_bus_axi4_0_r_bits_last,
  input [1:0] interrupts) ; 
   wire _bootROMDomainWrapper_auto_bootrom_in_a_ready ;  
   wire _bootROMDomainWrapper_auto_bootrom_in_d_valid ;  
   wire [1:0] _bootROMDomainWrapper_auto_bootrom_in_d_bits_size ;  
   wire [8:0] _bootROMDomainWrapper_auto_bootrom_in_d_bits_source ;  
   wire [63:0] _bootROMDomainWrapper_auto_bootrom_in_d_bits_data ;  
   wire _intsource_2_auto_out_sync_0 ;  
   wire _intsource_2_auto_out_sync_1 ;  
   wire _intsource_1_auto_out_sync_0 ;  
   wire _intsource_auto_out_sync_0 ;  
   wire _intsource_auto_out_sync_1 ;  
   wire _tlDM_auto_dmInner_dmInner_tl_in_a_ready ;  
   wire _tlDM_auto_dmInner_dmInner_tl_in_d_valid ;  
   wire [2:0] _tlDM_auto_dmInner_dmInner_tl_in_d_bits_opcode ;  
   wire [1:0] _tlDM_auto_dmInner_dmInner_tl_in_d_bits_size ;  
   wire [8:0] _tlDM_auto_dmInner_dmInner_tl_in_d_bits_source ;  
   wire [63:0] _tlDM_auto_dmInner_dmInner_tl_in_d_bits_data ;  
   wire _tlDM_auto_dmOuter_intsource_out_sync_0 ;  
   wire _tileHartIdNexusNode_auto_out ;  
   wire _clint_auto_int_out_0 ;  
   wire _clint_auto_int_out_1 ;  
   wire _clint_auto_in_a_ready ;  
   wire _clint_auto_in_d_valid ;  
   wire [2:0] _clint_auto_in_d_bits_opcode ;  
   wire [1:0] _clint_auto_in_d_bits_size ;  
   wire [8:0] _clint_auto_in_d_bits_source ;  
   wire [63:0] _clint_auto_in_d_bits_data ;  
   wire _plicDomainWrapper_auto_plic_int_out_0 ;  
   wire _plicDomainWrapper_auto_plic_in_a_ready ;  
   wire _plicDomainWrapper_auto_plic_in_d_valid ;  
   wire [2:0] _plicDomainWrapper_auto_plic_in_d_bits_opcode ;  
   wire [1:0] _plicDomainWrapper_auto_plic_in_d_bits_size ;  
   wire [8:0] _plicDomainWrapper_auto_plic_in_d_bits_source ;  
   wire [63:0] _plicDomainWrapper_auto_plic_in_d_bits_data ;  
   wire _tile_prci_domain_auto_tl_master_clock_xing_out_a_valid ;  
   wire [2:0] _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode ;  
   wire [2:0] _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param ;  
   wire [3:0] _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size ;  
   wire [1:0] _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source ;  
   wire [31:0] _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address ;  
   wire [7:0] _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask ;  
   wire [63:0] _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data ;  
   wire _tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_corrupt ;  
   wire _tile_prci_domain_auto_tl_master_clock_xing_out_b_ready ;  
   wire _tile_prci_domain_auto_tl_master_clock_xing_out_c_valid ;  
   wire [2:0] _tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_opcode ;  
   wire [2:0] _tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_param ;  
   wire [3:0] _tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_size ;  
   wire [1:0] _tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_source ;  
   wire [31:0] _tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_address ;  
   wire [63:0] _tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_data ;  
   wire _tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_corrupt ;  
   wire _tile_prci_domain_auto_tl_master_clock_xing_out_d_ready ;  
   wire _tile_prci_domain_auto_tl_master_clock_xing_out_e_valid ;  
   wire [1:0] _tile_prci_domain_auto_tl_master_clock_xing_out_e_bits_sink ;  
   wire _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid ;  
   wire [2:0] _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode ;  
   wire [2:0] _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_param ;  
   wire [2:0] _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size ;  
   wire [6:0] _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source ;  
   wire [31:0] _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address ;  
   wire [7:0] _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask ;  
   wire [63:0] _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data ;  
   wire _subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready ;  
   wire _subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready ;  
   wire _subsystem_l2_wrapper_auto_coherent_jbar_in_b_valid ;  
   wire [1:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_param ;  
   wire [31:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_address ;  
   wire _subsystem_l2_wrapper_auto_coherent_jbar_in_c_ready ;  
   wire _subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid ;  
   wire [2:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode ;  
   wire [1:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_param ;  
   wire [2:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size ;  
   wire [4:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source ;  
   wire [1:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_sink ;  
   wire _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied ;  
   wire [63:0] _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data ;  
   wire _subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt ;  
   wire _subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock ;  
   wire _subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset ;  
   wire _subsystem_mbus_auto_bus_xing_in_a_ready ;  
   wire _subsystem_mbus_auto_bus_xing_in_d_valid ;  
   wire [2:0] _subsystem_mbus_auto_bus_xing_in_d_bits_opcode ;  
   wire [2:0] _subsystem_mbus_auto_bus_xing_in_d_bits_size ;  
   wire [6:0] _subsystem_mbus_auto_bus_xing_in_d_bits_source ;  
   wire _subsystem_mbus_auto_bus_xing_in_d_bits_denied ;  
   wire [63:0] _subsystem_mbus_auto_bus_xing_in_d_bits_data ;  
   wire _subsystem_mbus_auto_bus_xing_in_d_bits_corrupt ;  
   wire _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_param ;  
   wire [1:0] _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size ;  
   wire [8:0] _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source ;  
   wire [16:0] _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address ;  
   wire [7:0] _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_mask ;  
   wire _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt ;  
   wire _subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready ;  
   wire _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_valid ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_opcode ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_param ;  
   wire [1:0] _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_size ;  
   wire [8:0] _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_source ;  
   wire [11:0] _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_address ;  
   wire [7:0] _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_mask ;  
   wire [63:0] _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_data ;  
   wire _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_corrupt ;  
   wire _subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_ready ;  
   wire _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_param ;  
   wire [1:0] _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size ;  
   wire [8:0] _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source ;  
   wire [25:0] _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address ;  
   wire [7:0] _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask ;  
   wire [63:0] _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data ;  
   wire _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_corrupt ;  
   wire _subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready ;  
   wire _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode ;  
   wire [2:0] _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_param ;  
   wire [1:0] _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size ;  
   wire [8:0] _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source ;  
   wire [27:0] _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address ;  
   wire [7:0] _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask ;  
   wire [63:0] _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data ;  
   wire _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_corrupt ;  
   wire _subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready ;  
   wire _subsystem_cbus_auto_fixedClockNode_out_2_clock ;  
   wire _subsystem_cbus_auto_fixedClockNode_out_2_reset ;  
   wire _subsystem_cbus_auto_fixedClockNode_out_0_clock ;  
   wire _subsystem_cbus_auto_fixedClockNode_out_0_reset ;  
   wire _subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock ;  
   wire _subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset ;  
   wire _subsystem_cbus_auto_bus_xing_in_a_ready ;  
   wire _subsystem_cbus_auto_bus_xing_in_d_valid ;  
   wire [2:0] _subsystem_cbus_auto_bus_xing_in_d_bits_opcode ;  
   wire [1:0] _subsystem_cbus_auto_bus_xing_in_d_bits_param ;  
   wire [3:0] _subsystem_cbus_auto_bus_xing_in_d_bits_size ;  
   wire [4:0] _subsystem_cbus_auto_bus_xing_in_d_bits_source ;  
   wire _subsystem_cbus_auto_bus_xing_in_d_bits_sink ;  
   wire _subsystem_cbus_auto_bus_xing_in_d_bits_denied ;  
   wire [63:0] _subsystem_cbus_auto_bus_xing_in_d_bits_data ;  
   wire _subsystem_cbus_auto_bus_xing_in_d_bits_corrupt ;  
   wire _subsystem_cbus_clock ;  
   wire _subsystem_cbus_reset ;  
   wire _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_valid ;  
   wire [2:0] _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_opcode ;  
   wire [2:0] _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_param ;  
   wire [3:0] _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_size ;  
   wire [3:0] _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_source ;  
   wire [31:0] _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_address ;  
   wire [7:0] _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_mask ;  
   wire [63:0] _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_data ;  
   wire _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_corrupt ;  
   wire _subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_ready ;  
   wire _subsystem_fbus_buffer_auto_in_a_ready ;  
   wire _subsystem_fbus_buffer_auto_in_d_valid ;  
   wire [2:0] _subsystem_fbus_buffer_auto_in_d_bits_opcode ;  
   wire [1:0] _subsystem_fbus_buffer_auto_in_d_bits_param ;  
   wire [3:0] _subsystem_fbus_buffer_auto_in_d_bits_size ;  
   wire [3:0] _subsystem_fbus_buffer_auto_in_d_bits_source ;  
   wire [1:0] _subsystem_fbus_buffer_auto_in_d_bits_sink ;  
   wire _subsystem_fbus_buffer_auto_in_d_bits_denied ;  
   wire [63:0] _subsystem_fbus_buffer_auto_in_d_bits_data ;  
   wire _subsystem_fbus_buffer_auto_in_d_bits_corrupt ;  
   wire _subsystem_fbus_buffer_auto_out_a_valid ;  
   wire [2:0] _subsystem_fbus_buffer_auto_out_a_bits_opcode ;  
   wire [2:0] _subsystem_fbus_buffer_auto_out_a_bits_param ;  
   wire [3:0] _subsystem_fbus_buffer_auto_out_a_bits_size ;  
   wire [3:0] _subsystem_fbus_buffer_auto_out_a_bits_source ;  
   wire [31:0] _subsystem_fbus_buffer_auto_out_a_bits_address ;  
   wire [7:0] _subsystem_fbus_buffer_auto_out_a_bits_mask ;  
   wire [63:0] _subsystem_fbus_buffer_auto_out_a_bits_data ;  
   wire _subsystem_fbus_buffer_auto_out_a_bits_corrupt ;  
   wire _subsystem_fbus_buffer_auto_out_d_ready ;  
   wire _subsystem_pbus_clock ;  
   wire _subsystem_pbus_reset ;  
   wire _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready ;  
   wire _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_valid ;  
   wire [1:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param ;  
   wire [31:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address ;  
   wire _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_ready ;  
   wire _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid ;  
   wire [2:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode ;  
   wire [1:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param ;  
   wire [3:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size ;  
   wire [1:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source ;  
   wire [1:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink ;  
   wire _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied ;  
   wire [63:0] _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data ;  
   wire _subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size ;  
   wire [4:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source ;  
   wire [31:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address ;  
   wire [7:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask ;  
   wire [63:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_corrupt ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size ;  
   wire [4:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source ;  
   wire [31:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address ;  
   wire [63:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_corrupt ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid ;  
   wire [1:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink ;  
   wire _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready ;  
   wire _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid ;  
   wire [2:0] _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode ;  
   wire [1:0] _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param ;  
   wire [3:0] _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size ;  
   wire [3:0] _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source ;  
   wire [1:0] _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink ;  
   wire _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied ;  
   wire [63:0] _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data ;  
   wire _subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode ;  
   wire [2:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param ;  
   wire [3:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size ;  
   wire [4:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source ;  
   wire [27:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address ;  
   wire [7:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask ;  
   wire [63:0] _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt ;  
   wire _subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready ;  
   wire _subsystem_sbus_auto_fixedClockNode_out_1_clock ;  
   wire _subsystem_sbus_auto_fixedClockNode_out_1_reset ;  
   wire _subsystem_sbus_auto_fixedClockNode_out_0_clock ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock ;  
   wire _subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock ;  
   wire _dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset ;  
   wire _ibus_intsink_auto_out_0 ;  
   wire _ibus_intsink_auto_out_1 ;  
   wire _ibus_int_bus_auto_int_out_0 ;  
   wire _ibus_int_bus_auto_int_out_1 ;  
   reg [6:0] int_rtc_tick_c_value ;  
   wire int_rtc_tick=int_rtc_tick_c_value==7'h63 ;  
  always @( posedge _subsystem_pbus_clock)
       begin 
         if (_subsystem_pbus_reset)
            int_rtc_tick_c_value <=7'h0;
          else 
            if (int_rtc_tick)
               int_rtc_tick_c_value <=7'h0;
             else 
               int_rtc_tick_c_value <=int_rtc_tick_c_value+7'h1;
       end
  
  IntXbar ibus_int_bus(.auto_int_in_0(_ibus_intsink_auto_out_0),.auto_int_in_1(_ibus_intsink_auto_out_1),.auto_int_out_0(_ibus_int_bus_auto_int_out_0),.auto_int_out_1(_ibus_int_bus_auto_int_out_1)); 
  IntSyncAsyncCrossingSink ibus_intsink(.clock(_subsystem_sbus_auto_fixedClockNode_out_0_clock),.auto_in_sync_0(_intsource_2_auto_out_sync_0),.auto_in_sync_1(_intsource_2_auto_out_sync_1),.auto_out_0(_ibus_intsink_auto_out_0),.auto_out_1(_ibus_intsink_auto_out_1)); 
  SimpleClockGroupSource dummyClockGroupSourceNode(.clock(clock),.reset(reset),.auto_out_member_subsystem_sbus_5_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock),.auto_out_member_subsystem_sbus_5_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset),.auto_out_member_subsystem_sbus_4_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock),.auto_out_member_subsystem_sbus_4_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset),.auto_out_member_subsystem_sbus_3_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock),.auto_out_member_subsystem_sbus_3_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset),.auto_out_member_subsystem_sbus_2_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock),.auto_out_member_subsystem_sbus_2_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset),.auto_out_member_subsystem_sbus_1_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock),.auto_out_member_subsystem_sbus_1_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset),.auto_out_member_subsystem_sbus_0_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock),.auto_out_member_subsystem_sbus_0_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset)); 
  SystemBus subsystem_sbus(.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_ready(mmio_axi4_0_aw_ready),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_valid(mmio_axi4_0_aw_valid),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_id(mmio_axi4_0_aw_bits_id),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_addr(mmio_axi4_0_aw_bits_addr),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_len(mmio_axi4_0_aw_bits_len),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_size(mmio_axi4_0_aw_bits_size),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_burst(mmio_axi4_0_aw_bits_burst),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_lock(mmio_axi4_0_aw_bits_lock),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_cache(mmio_axi4_0_aw_bits_cache),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_prot(mmio_axi4_0_aw_bits_prot),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_aw_bits_qos(mmio_axi4_0_aw_bits_qos),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_ready(mmio_axi4_0_w_ready),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_valid(mmio_axi4_0_w_valid),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_data(mmio_axi4_0_w_bits_data),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_strb(mmio_axi4_0_w_bits_strb),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_w_bits_last(mmio_axi4_0_w_bits_last),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_ready(mmio_axi4_0_b_ready),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_valid(mmio_axi4_0_b_valid),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_bits_id(mmio_axi4_0_b_bits_id),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_b_bits_resp(mmio_axi4_0_b_bits_resp),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_ready(mmio_axi4_0_ar_ready),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_valid(mmio_axi4_0_ar_valid),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_id(mmio_axi4_0_ar_bits_id),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_addr(mmio_axi4_0_ar_bits_addr),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_len(mmio_axi4_0_ar_bits_len),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_size(mmio_axi4_0_ar_bits_size),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_burst(mmio_axi4_0_ar_bits_burst),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_lock(mmio_axi4_0_ar_bits_lock),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_cache(mmio_axi4_0_ar_bits_cache),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_prot(mmio_axi4_0_ar_bits_prot),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_ar_bits_qos(mmio_axi4_0_ar_bits_qos),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_ready(mmio_axi4_0_r_ready),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_valid(mmio_axi4_0_r_valid),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_id(mmio_axi4_0_r_bits_id),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_data(mmio_axi4_0_r_bits_data),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_resp(mmio_axi4_0_r_bits_resp),.auto_coupler_to_port_named_mmio_port_axi4_axi4buf_out_r_bits_last(mmio_axi4_0_r_bits_last),.auto_coupler_from_tile_tl_master_clock_xing_in_a_ready(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready),.auto_coupler_from_tile_tl_master_clock_xing_in_a_valid(_tile_prci_domain_auto_tl_master_clock_xing_out_a_valid),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_opcode(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_param(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_size(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_source(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_address(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_mask(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_data(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data),.auto_coupler_from_tile_tl_master_clock_xing_in_a_bits_corrupt(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_corrupt),.auto_coupler_from_tile_tl_master_clock_xing_in_b_ready(_tile_prci_domain_auto_tl_master_clock_xing_out_b_ready),.auto_coupler_from_tile_tl_master_clock_xing_in_b_valid(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_valid),.auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param),.auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address),.auto_coupler_from_tile_tl_master_clock_xing_in_c_ready(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_ready),.auto_coupler_from_tile_tl_master_clock_xing_in_c_valid(_tile_prci_domain_auto_tl_master_clock_xing_out_c_valid),.auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_opcode(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_opcode),.auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_param(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_param),.auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_size(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_size),.auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_source(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_source),.auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_address(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_address),.auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_data(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_data),.auto_coupler_from_tile_tl_master_clock_xing_in_c_bits_corrupt(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_corrupt),.auto_coupler_from_tile_tl_master_clock_xing_in_d_ready(_tile_prci_domain_auto_tl_master_clock_xing_out_d_ready),.auto_coupler_from_tile_tl_master_clock_xing_in_d_valid(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data),.auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt),.auto_coupler_from_tile_tl_master_clock_xing_in_e_valid(_tile_prci_domain_auto_tl_master_clock_xing_out_e_valid),.auto_coupler_from_tile_tl_master_clock_xing_in_e_bits_sink(_tile_prci_domain_auto_tl_master_clock_xing_out_e_bits_sink),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_ready(_subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data),.auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_corrupt(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_corrupt),.auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready),.auto_coupler_to_bus_named_subsystem_l2_widget_out_b_valid(_subsystem_l2_wrapper_auto_coherent_jbar_in_b_valid),.auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_param(_subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_param),.auto_coupler_to_bus_named_subsystem_l2_widget_out_b_bits_address(_subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_address),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_ready(_subsystem_l2_wrapper_auto_coherent_jbar_in_c_ready),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data),.auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_corrupt(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_corrupt),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_valid(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_opcode(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_param(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_param),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_size(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_source(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_sink(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_sink),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_denied(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_data(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data),.auto_coupler_to_bus_named_subsystem_l2_widget_out_d_bits_corrupt(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt),.auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid),.auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_valid(_subsystem_fbus_buffer_auto_out_a_valid),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_opcode(_subsystem_fbus_buffer_auto_out_a_bits_opcode),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_param(_subsystem_fbus_buffer_auto_out_a_bits_param),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_size(_subsystem_fbus_buffer_auto_out_a_bits_size),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_source(_subsystem_fbus_buffer_auto_out_a_bits_source),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_address(_subsystem_fbus_buffer_auto_out_a_bits_address),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_mask(_subsystem_fbus_buffer_auto_out_a_bits_mask),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_data(_subsystem_fbus_buffer_auto_out_a_bits_data),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_bits_corrupt(_subsystem_fbus_buffer_auto_out_a_bits_corrupt),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_ready(_subsystem_fbus_buffer_auto_out_d_ready),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data),.auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_ready(_subsystem_cbus_auto_bus_xing_in_a_ready),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_valid(_subsystem_cbus_auto_bus_xing_in_d_valid),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_opcode(_subsystem_cbus_auto_bus_xing_in_d_bits_opcode),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_param(_subsystem_cbus_auto_bus_xing_in_d_bits_param),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_size(_subsystem_cbus_auto_bus_xing_in_d_bits_size),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_source(_subsystem_cbus_auto_bus_xing_in_d_bits_source),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_sink(_subsystem_cbus_auto_bus_xing_in_d_bits_sink),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_denied(_subsystem_cbus_auto_bus_xing_in_d_bits_denied),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_data(_subsystem_cbus_auto_bus_xing_in_d_bits_data),.auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_bits_corrupt(_subsystem_cbus_auto_bus_xing_in_d_bits_corrupt),.auto_fixedClockNode_out_1_clock(_subsystem_sbus_auto_fixedClockNode_out_1_clock),.auto_fixedClockNode_out_1_reset(_subsystem_sbus_auto_fixedClockNode_out_1_reset),.auto_fixedClockNode_out_0_clock(_subsystem_sbus_auto_fixedClockNode_out_0_clock),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_clock),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_5_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_5_reset),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_clock),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_4_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_4_reset),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_clock),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_3_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_3_reset),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_clock),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_2_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_2_reset),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_clock),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_1_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_1_reset),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_clock(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_clock),.auto_subsystem_sbus_clock_groups_in_member_subsystem_sbus_0_reset(_dummyClockGroupSourceNode_auto_out_member_subsystem_sbus_0_reset),.auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock),.auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset),.auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock),.auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset),.auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock),.auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset),.auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock),.auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset),.auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock),.auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset)); 
  PeripheryBus subsystem_pbus(.auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_clock(_subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock),.auto_subsystem_pbus_clock_groups_in_member_subsystem_pbus_0_reset(_subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset),.clock(_subsystem_pbus_clock),.reset(_subsystem_pbus_reset)); 
  TLBuffer_2 subsystem_fbus_buffer(.clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock),.reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset),.auto_in_a_ready(_subsystem_fbus_buffer_auto_in_a_ready),.auto_in_a_valid(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_valid),.auto_in_a_bits_opcode(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_opcode),.auto_in_a_bits_param(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_param),.auto_in_a_bits_size(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_size),.auto_in_a_bits_source(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_source),.auto_in_a_bits_address(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_address),.auto_in_a_bits_mask(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_mask),.auto_in_a_bits_data(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_data),.auto_in_a_bits_corrupt(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_corrupt),.auto_in_d_ready(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_ready),.auto_in_d_valid(_subsystem_fbus_buffer_auto_in_d_valid),.auto_in_d_bits_opcode(_subsystem_fbus_buffer_auto_in_d_bits_opcode),.auto_in_d_bits_param(_subsystem_fbus_buffer_auto_in_d_bits_param),.auto_in_d_bits_size(_subsystem_fbus_buffer_auto_in_d_bits_size),.auto_in_d_bits_source(_subsystem_fbus_buffer_auto_in_d_bits_source),.auto_in_d_bits_sink(_subsystem_fbus_buffer_auto_in_d_bits_sink),.auto_in_d_bits_denied(_subsystem_fbus_buffer_auto_in_d_bits_denied),.auto_in_d_bits_data(_subsystem_fbus_buffer_auto_in_d_bits_data),.auto_in_d_bits_corrupt(_subsystem_fbus_buffer_auto_in_d_bits_corrupt),.auto_out_a_ready(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_a_ready),.auto_out_a_valid(_subsystem_fbus_buffer_auto_out_a_valid),.auto_out_a_bits_opcode(_subsystem_fbus_buffer_auto_out_a_bits_opcode),.auto_out_a_bits_param(_subsystem_fbus_buffer_auto_out_a_bits_param),.auto_out_a_bits_size(_subsystem_fbus_buffer_auto_out_a_bits_size),.auto_out_a_bits_source(_subsystem_fbus_buffer_auto_out_a_bits_source),.auto_out_a_bits_address(_subsystem_fbus_buffer_auto_out_a_bits_address),.auto_out_a_bits_mask(_subsystem_fbus_buffer_auto_out_a_bits_mask),.auto_out_a_bits_data(_subsystem_fbus_buffer_auto_out_a_bits_data),.auto_out_a_bits_corrupt(_subsystem_fbus_buffer_auto_out_a_bits_corrupt),.auto_out_d_ready(_subsystem_fbus_buffer_auto_out_d_ready),.auto_out_d_valid(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_valid),.auto_out_d_bits_opcode(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_opcode),.auto_out_d_bits_param(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_param),.auto_out_d_bits_size(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_size),.auto_out_d_bits_source(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_source),.auto_out_d_bits_sink(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_sink),.auto_out_d_bits_denied(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_denied),.auto_out_d_bits_data(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_data),.auto_out_d_bits_corrupt(_subsystem_sbus_auto_coupler_from_bus_named_subsystem_fbus_bus_xing_in_d_bits_corrupt)); 
  TLInterconnectCoupler_5 subsystem_fbus_coupler_from_port_named_slave_port_axi4(.clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_clock),.reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_1_member_subsystem_fbus_0_reset),.auto_axi4index_in_aw_ready(l2_frontend_bus_axi4_0_aw_ready),.auto_axi4index_in_aw_valid(l2_frontend_bus_axi4_0_aw_valid),.auto_axi4index_in_aw_bits_id(l2_frontend_bus_axi4_0_aw_bits_id),.auto_axi4index_in_aw_bits_addr(l2_frontend_bus_axi4_0_aw_bits_addr),.auto_axi4index_in_aw_bits_len(l2_frontend_bus_axi4_0_aw_bits_len),.auto_axi4index_in_aw_bits_size(l2_frontend_bus_axi4_0_aw_bits_size),.auto_axi4index_in_aw_bits_burst(l2_frontend_bus_axi4_0_aw_bits_burst),.auto_axi4index_in_w_ready(l2_frontend_bus_axi4_0_w_ready),.auto_axi4index_in_w_valid(l2_frontend_bus_axi4_0_w_valid),.auto_axi4index_in_w_bits_data(l2_frontend_bus_axi4_0_w_bits_data),.auto_axi4index_in_w_bits_strb(l2_frontend_bus_axi4_0_w_bits_strb),.auto_axi4index_in_w_bits_last(l2_frontend_bus_axi4_0_w_bits_last),.auto_axi4index_in_b_ready(l2_frontend_bus_axi4_0_b_ready),.auto_axi4index_in_b_valid(l2_frontend_bus_axi4_0_b_valid),.auto_axi4index_in_b_bits_id(l2_frontend_bus_axi4_0_b_bits_id),.auto_axi4index_in_b_bits_resp(l2_frontend_bus_axi4_0_b_bits_resp),.auto_axi4index_in_ar_ready(l2_frontend_bus_axi4_0_ar_ready),.auto_axi4index_in_ar_valid(l2_frontend_bus_axi4_0_ar_valid),.auto_axi4index_in_ar_bits_id(l2_frontend_bus_axi4_0_ar_bits_id),.auto_axi4index_in_ar_bits_addr(l2_frontend_bus_axi4_0_ar_bits_addr),.auto_axi4index_in_ar_bits_len(l2_frontend_bus_axi4_0_ar_bits_len),.auto_axi4index_in_ar_bits_size(l2_frontend_bus_axi4_0_ar_bits_size),.auto_axi4index_in_ar_bits_burst(l2_frontend_bus_axi4_0_ar_bits_burst),.auto_axi4index_in_r_ready(l2_frontend_bus_axi4_0_r_ready),.auto_axi4index_in_r_valid(l2_frontend_bus_axi4_0_r_valid),.auto_axi4index_in_r_bits_id(l2_frontend_bus_axi4_0_r_bits_id),.auto_axi4index_in_r_bits_data(l2_frontend_bus_axi4_0_r_bits_data),.auto_axi4index_in_r_bits_resp(l2_frontend_bus_axi4_0_r_bits_resp),.auto_axi4index_in_r_bits_last(l2_frontend_bus_axi4_0_r_bits_last),.auto_tl_out_a_ready(_subsystem_fbus_buffer_auto_in_a_ready),.auto_tl_out_a_valid(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_valid),.auto_tl_out_a_bits_opcode(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_opcode),.auto_tl_out_a_bits_param(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_param),.auto_tl_out_a_bits_size(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_size),.auto_tl_out_a_bits_source(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_source),.auto_tl_out_a_bits_address(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_address),.auto_tl_out_a_bits_mask(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_mask),.auto_tl_out_a_bits_data(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_data),.auto_tl_out_a_bits_corrupt(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_a_bits_corrupt),.auto_tl_out_d_ready(_subsystem_fbus_coupler_from_port_named_slave_port_axi4_auto_tl_out_d_ready),.auto_tl_out_d_valid(_subsystem_fbus_buffer_auto_in_d_valid),.auto_tl_out_d_bits_opcode(_subsystem_fbus_buffer_auto_in_d_bits_opcode),.auto_tl_out_d_bits_param(_subsystem_fbus_buffer_auto_in_d_bits_param),.auto_tl_out_d_bits_size(_subsystem_fbus_buffer_auto_in_d_bits_size),.auto_tl_out_d_bits_source(_subsystem_fbus_buffer_auto_in_d_bits_source),.auto_tl_out_d_bits_sink(_subsystem_fbus_buffer_auto_in_d_bits_sink),.auto_tl_out_d_bits_denied(_subsystem_fbus_buffer_auto_in_d_bits_denied),.auto_tl_out_d_bits_data(_subsystem_fbus_buffer_auto_in_d_bits_data),.auto_tl_out_d_bits_corrupt(_subsystem_fbus_buffer_auto_in_d_bits_corrupt)); 
  PeripheryBus_1 subsystem_cbus(.auto_coupler_to_bootrom_fragmenter_out_a_ready(_bootROMDomainWrapper_auto_bootrom_in_a_ready),.auto_coupler_to_bootrom_fragmenter_out_a_valid(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid),.auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode),.auto_coupler_to_bootrom_fragmenter_out_a_bits_param(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_param),.auto_coupler_to_bootrom_fragmenter_out_a_bits_size(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size),.auto_coupler_to_bootrom_fragmenter_out_a_bits_source(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source),.auto_coupler_to_bootrom_fragmenter_out_a_bits_address(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address),.auto_coupler_to_bootrom_fragmenter_out_a_bits_mask(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_mask),.auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt),.auto_coupler_to_bootrom_fragmenter_out_d_ready(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready),.auto_coupler_to_bootrom_fragmenter_out_d_valid(_bootROMDomainWrapper_auto_bootrom_in_d_valid),.auto_coupler_to_bootrom_fragmenter_out_d_bits_size(_bootROMDomainWrapper_auto_bootrom_in_d_bits_size),.auto_coupler_to_bootrom_fragmenter_out_d_bits_source(_bootROMDomainWrapper_auto_bootrom_in_d_bits_source),.auto_coupler_to_bootrom_fragmenter_out_d_bits_data(_bootROMDomainWrapper_auto_bootrom_in_d_bits_data),.auto_coupler_to_debug_fragmenter_out_a_ready(_tlDM_auto_dmInner_dmInner_tl_in_a_ready),.auto_coupler_to_debug_fragmenter_out_a_valid(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_valid),.auto_coupler_to_debug_fragmenter_out_a_bits_opcode(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_opcode),.auto_coupler_to_debug_fragmenter_out_a_bits_param(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_param),.auto_coupler_to_debug_fragmenter_out_a_bits_size(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_size),.auto_coupler_to_debug_fragmenter_out_a_bits_source(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_source),.auto_coupler_to_debug_fragmenter_out_a_bits_address(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_address),.auto_coupler_to_debug_fragmenter_out_a_bits_mask(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_mask),.auto_coupler_to_debug_fragmenter_out_a_bits_data(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_data),.auto_coupler_to_debug_fragmenter_out_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_corrupt),.auto_coupler_to_debug_fragmenter_out_d_ready(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_ready),.auto_coupler_to_debug_fragmenter_out_d_valid(_tlDM_auto_dmInner_dmInner_tl_in_d_valid),.auto_coupler_to_debug_fragmenter_out_d_bits_opcode(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_opcode),.auto_coupler_to_debug_fragmenter_out_d_bits_size(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_size),.auto_coupler_to_debug_fragmenter_out_d_bits_source(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_source),.auto_coupler_to_debug_fragmenter_out_d_bits_data(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_data),.auto_coupler_to_clint_fragmenter_out_a_ready(_clint_auto_in_a_ready),.auto_coupler_to_clint_fragmenter_out_a_valid(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid),.auto_coupler_to_clint_fragmenter_out_a_bits_opcode(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode),.auto_coupler_to_clint_fragmenter_out_a_bits_param(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_param),.auto_coupler_to_clint_fragmenter_out_a_bits_size(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size),.auto_coupler_to_clint_fragmenter_out_a_bits_source(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source),.auto_coupler_to_clint_fragmenter_out_a_bits_address(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address),.auto_coupler_to_clint_fragmenter_out_a_bits_mask(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask),.auto_coupler_to_clint_fragmenter_out_a_bits_data(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data),.auto_coupler_to_clint_fragmenter_out_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_corrupt),.auto_coupler_to_clint_fragmenter_out_d_ready(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready),.auto_coupler_to_clint_fragmenter_out_d_valid(_clint_auto_in_d_valid),.auto_coupler_to_clint_fragmenter_out_d_bits_opcode(_clint_auto_in_d_bits_opcode),.auto_coupler_to_clint_fragmenter_out_d_bits_size(_clint_auto_in_d_bits_size),.auto_coupler_to_clint_fragmenter_out_d_bits_source(_clint_auto_in_d_bits_source),.auto_coupler_to_clint_fragmenter_out_d_bits_data(_clint_auto_in_d_bits_data),.auto_coupler_to_plic_fragmenter_out_a_ready(_plicDomainWrapper_auto_plic_in_a_ready),.auto_coupler_to_plic_fragmenter_out_a_valid(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid),.auto_coupler_to_plic_fragmenter_out_a_bits_opcode(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode),.auto_coupler_to_plic_fragmenter_out_a_bits_param(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_param),.auto_coupler_to_plic_fragmenter_out_a_bits_size(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size),.auto_coupler_to_plic_fragmenter_out_a_bits_source(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source),.auto_coupler_to_plic_fragmenter_out_a_bits_address(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address),.auto_coupler_to_plic_fragmenter_out_a_bits_mask(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask),.auto_coupler_to_plic_fragmenter_out_a_bits_data(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data),.auto_coupler_to_plic_fragmenter_out_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_corrupt),.auto_coupler_to_plic_fragmenter_out_d_ready(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready),.auto_coupler_to_plic_fragmenter_out_d_valid(_plicDomainWrapper_auto_plic_in_d_valid),.auto_coupler_to_plic_fragmenter_out_d_bits_opcode(_plicDomainWrapper_auto_plic_in_d_bits_opcode),.auto_coupler_to_plic_fragmenter_out_d_bits_size(_plicDomainWrapper_auto_plic_in_d_bits_size),.auto_coupler_to_plic_fragmenter_out_d_bits_source(_plicDomainWrapper_auto_plic_in_d_bits_source),.auto_coupler_to_plic_fragmenter_out_d_bits_data(_plicDomainWrapper_auto_plic_in_d_bits_data),.auto_fixedClockNode_out_2_clock(_subsystem_cbus_auto_fixedClockNode_out_2_clock),.auto_fixedClockNode_out_2_reset(_subsystem_cbus_auto_fixedClockNode_out_2_reset),.auto_fixedClockNode_out_0_clock(_subsystem_cbus_auto_fixedClockNode_out_0_clock),.auto_fixedClockNode_out_0_reset(_subsystem_cbus_auto_fixedClockNode_out_0_reset),.auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_clock),.auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_1_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_1_reset),.auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_clock),.auto_subsystem_cbus_clock_groups_in_member_subsystem_cbus_0_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_0_member_subsystem_cbus_0_reset),.auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock(_subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_clock),.auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset(_subsystem_cbus_auto_subsystem_cbus_clock_groups_out_member_subsystem_pbus_0_reset),.auto_bus_xing_in_a_ready(_subsystem_cbus_auto_bus_xing_in_a_ready),.auto_bus_xing_in_a_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_valid),.auto_bus_xing_in_a_bits_opcode(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_opcode),.auto_bus_xing_in_a_bits_param(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_param),.auto_bus_xing_in_a_bits_size(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_size),.auto_bus_xing_in_a_bits_source(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_source),.auto_bus_xing_in_a_bits_address(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_address),.auto_bus_xing_in_a_bits_mask(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_mask),.auto_bus_xing_in_a_bits_data(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_data),.auto_bus_xing_in_a_bits_corrupt(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_a_bits_corrupt),.auto_bus_xing_in_d_ready(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_cbus_bus_xing_out_d_ready),.auto_bus_xing_in_d_valid(_subsystem_cbus_auto_bus_xing_in_d_valid),.auto_bus_xing_in_d_bits_opcode(_subsystem_cbus_auto_bus_xing_in_d_bits_opcode),.auto_bus_xing_in_d_bits_param(_subsystem_cbus_auto_bus_xing_in_d_bits_param),.auto_bus_xing_in_d_bits_size(_subsystem_cbus_auto_bus_xing_in_d_bits_size),.auto_bus_xing_in_d_bits_source(_subsystem_cbus_auto_bus_xing_in_d_bits_source),.auto_bus_xing_in_d_bits_sink(_subsystem_cbus_auto_bus_xing_in_d_bits_sink),.auto_bus_xing_in_d_bits_denied(_subsystem_cbus_auto_bus_xing_in_d_bits_denied),.auto_bus_xing_in_d_bits_data(_subsystem_cbus_auto_bus_xing_in_d_bits_data),.auto_bus_xing_in_d_bits_corrupt(_subsystem_cbus_auto_bus_xing_in_d_bits_corrupt),.clock(_subsystem_cbus_clock),.reset(_subsystem_cbus_reset)); 
  MemoryBus subsystem_mbus(.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_ready(mem_axi4_0_aw_ready),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_valid(mem_axi4_0_aw_valid),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_id(mem_axi4_0_aw_bits_id),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_addr(mem_axi4_0_aw_bits_addr),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_len(mem_axi4_0_aw_bits_len),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_aw_bits_size(mem_axi4_0_aw_bits_size),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_ready(mem_axi4_0_w_ready),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_valid(mem_axi4_0_w_valid),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_data(mem_axi4_0_w_bits_data),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_strb(mem_axi4_0_w_bits_strb),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_w_bits_last(mem_axi4_0_w_bits_last),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_ready(mem_axi4_0_b_ready),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_valid(mem_axi4_0_b_valid),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_id(mem_axi4_0_b_bits_id),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_b_bits_resp(mem_axi4_0_b_bits_resp),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_ready(mem_axi4_0_ar_ready),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_valid(mem_axi4_0_ar_valid),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_id(mem_axi4_0_ar_bits_id),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_addr(mem_axi4_0_ar_bits_addr),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_len(mem_axi4_0_ar_bits_len),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_ar_bits_size(mem_axi4_0_ar_bits_size),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_ready(mem_axi4_0_r_ready),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_valid(mem_axi4_0_r_valid),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_id(mem_axi4_0_r_bits_id),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_data(mem_axi4_0_r_bits_data),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_resp(mem_axi4_0_r_bits_resp),.auto_coupler_to_memory_controller_port_named_axi4_axi4yank_out_r_bits_last(mem_axi4_0_r_bits_last),.auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_clock(_subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock),.auto_subsystem_mbus_clock_groups_in_member_subsystem_mbus_0_reset(_subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset),.auto_bus_xing_in_a_ready(_subsystem_mbus_auto_bus_xing_in_a_ready),.auto_bus_xing_in_a_valid(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid),.auto_bus_xing_in_a_bits_opcode(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode),.auto_bus_xing_in_a_bits_param(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_param),.auto_bus_xing_in_a_bits_size(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size),.auto_bus_xing_in_a_bits_source(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source),.auto_bus_xing_in_a_bits_address(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address),.auto_bus_xing_in_a_bits_mask(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask),.auto_bus_xing_in_a_bits_data(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data),.auto_bus_xing_in_d_ready(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready),.auto_bus_xing_in_d_valid(_subsystem_mbus_auto_bus_xing_in_d_valid),.auto_bus_xing_in_d_bits_opcode(_subsystem_mbus_auto_bus_xing_in_d_bits_opcode),.auto_bus_xing_in_d_bits_size(_subsystem_mbus_auto_bus_xing_in_d_bits_size),.auto_bus_xing_in_d_bits_source(_subsystem_mbus_auto_bus_xing_in_d_bits_source),.auto_bus_xing_in_d_bits_denied(_subsystem_mbus_auto_bus_xing_in_d_bits_denied),.auto_bus_xing_in_d_bits_data(_subsystem_mbus_auto_bus_xing_in_d_bits_data),.auto_bus_xing_in_d_bits_corrupt(_subsystem_mbus_auto_bus_xing_in_d_bits_corrupt)); 
  CoherenceManagerWrapper subsystem_l2_wrapper(.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_ready(_subsystem_mbus_auto_bus_xing_in_a_ready),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_valid),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_opcode),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_param(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_param),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_size),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_source),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_address),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_mask),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_a_bits_data),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready(_subsystem_l2_wrapper_auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_ready),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_valid(_subsystem_mbus_auto_bus_xing_in_d_valid),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_opcode(_subsystem_mbus_auto_bus_xing_in_d_bits_opcode),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_size(_subsystem_mbus_auto_bus_xing_in_d_bits_size),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_source(_subsystem_mbus_auto_bus_xing_in_d_bits_source),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_denied(_subsystem_mbus_auto_bus_xing_in_d_bits_denied),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_data(_subsystem_mbus_auto_bus_xing_in_d_bits_data),.auto_coupler_to_bus_named_subsystem_mbus_bus_xing_out_d_bits_corrupt(_subsystem_mbus_auto_bus_xing_in_d_bits_corrupt),.auto_coherent_jbar_in_a_ready(_subsystem_l2_wrapper_auto_coherent_jbar_in_a_ready),.auto_coherent_jbar_in_a_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_valid),.auto_coherent_jbar_in_a_bits_opcode(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_opcode),.auto_coherent_jbar_in_a_bits_param(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_param),.auto_coherent_jbar_in_a_bits_size(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_size),.auto_coherent_jbar_in_a_bits_source(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_source),.auto_coherent_jbar_in_a_bits_address(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_address),.auto_coherent_jbar_in_a_bits_mask(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_mask),.auto_coherent_jbar_in_a_bits_data(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_data),.auto_coherent_jbar_in_a_bits_corrupt(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_a_bits_corrupt),.auto_coherent_jbar_in_b_ready(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_b_ready),.auto_coherent_jbar_in_b_valid(_subsystem_l2_wrapper_auto_coherent_jbar_in_b_valid),.auto_coherent_jbar_in_b_bits_param(_subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_param),.auto_coherent_jbar_in_b_bits_address(_subsystem_l2_wrapper_auto_coherent_jbar_in_b_bits_address),.auto_coherent_jbar_in_c_ready(_subsystem_l2_wrapper_auto_coherent_jbar_in_c_ready),.auto_coherent_jbar_in_c_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_valid),.auto_coherent_jbar_in_c_bits_opcode(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_opcode),.auto_coherent_jbar_in_c_bits_param(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_param),.auto_coherent_jbar_in_c_bits_size(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_size),.auto_coherent_jbar_in_c_bits_source(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_source),.auto_coherent_jbar_in_c_bits_address(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_address),.auto_coherent_jbar_in_c_bits_data(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_data),.auto_coherent_jbar_in_c_bits_corrupt(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_c_bits_corrupt),.auto_coherent_jbar_in_d_ready(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_d_ready),.auto_coherent_jbar_in_d_valid(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_valid),.auto_coherent_jbar_in_d_bits_opcode(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_opcode),.auto_coherent_jbar_in_d_bits_param(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_param),.auto_coherent_jbar_in_d_bits_size(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_size),.auto_coherent_jbar_in_d_bits_source(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_source),.auto_coherent_jbar_in_d_bits_sink(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_sink),.auto_coherent_jbar_in_d_bits_denied(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_denied),.auto_coherent_jbar_in_d_bits_data(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_data),.auto_coherent_jbar_in_d_bits_corrupt(_subsystem_l2_wrapper_auto_coherent_jbar_in_d_bits_corrupt),.auto_coherent_jbar_in_e_valid(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_valid),.auto_coherent_jbar_in_e_bits_sink(_subsystem_sbus_auto_coupler_to_bus_named_subsystem_l2_widget_out_e_bits_sink),.auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_clock),.auto_subsystem_l2_clock_groups_in_member_subsystem_l2_1_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_1_reset),.auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_clock(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_clock),.auto_subsystem_l2_clock_groups_in_member_subsystem_l2_0_reset(_subsystem_sbus_auto_subsystem_sbus_clock_groups_out_2_member_subsystem_l2_0_reset),.auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock(_subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_clock),.auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset(_subsystem_l2_wrapper_auto_subsystem_l2_clock_groups_out_member_subsystem_mbus_0_reset)); 
  TilePRCIDomain tile_prci_domain(.auto_intsink_in_sync_0(_tlDM_auto_dmOuter_intsource_out_sync_0),.auto_tile_reset_domain_tile_hartid_in(_tileHartIdNexusNode_auto_out),.auto_int_in_clock_xing_in_1_sync_0(_intsource_1_auto_out_sync_0),.auto_int_in_clock_xing_in_0_sync_0(_intsource_auto_out_sync_0),.auto_int_in_clock_xing_in_0_sync_1(_intsource_auto_out_sync_1),.auto_tl_master_clock_xing_out_a_ready(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_a_ready),.auto_tl_master_clock_xing_out_a_valid(_tile_prci_domain_auto_tl_master_clock_xing_out_a_valid),.auto_tl_master_clock_xing_out_a_bits_opcode(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_opcode),.auto_tl_master_clock_xing_out_a_bits_param(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_param),.auto_tl_master_clock_xing_out_a_bits_size(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_size),.auto_tl_master_clock_xing_out_a_bits_source(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_source),.auto_tl_master_clock_xing_out_a_bits_address(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_address),.auto_tl_master_clock_xing_out_a_bits_mask(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_mask),.auto_tl_master_clock_xing_out_a_bits_data(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_data),.auto_tl_master_clock_xing_out_a_bits_corrupt(_tile_prci_domain_auto_tl_master_clock_xing_out_a_bits_corrupt),.auto_tl_master_clock_xing_out_b_ready(_tile_prci_domain_auto_tl_master_clock_xing_out_b_ready),.auto_tl_master_clock_xing_out_b_valid(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_valid),.auto_tl_master_clock_xing_out_b_bits_param(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_param),.auto_tl_master_clock_xing_out_b_bits_address(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_b_bits_address),.auto_tl_master_clock_xing_out_c_ready(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_c_ready),.auto_tl_master_clock_xing_out_c_valid(_tile_prci_domain_auto_tl_master_clock_xing_out_c_valid),.auto_tl_master_clock_xing_out_c_bits_opcode(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_opcode),.auto_tl_master_clock_xing_out_c_bits_param(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_param),.auto_tl_master_clock_xing_out_c_bits_size(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_size),.auto_tl_master_clock_xing_out_c_bits_source(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_source),.auto_tl_master_clock_xing_out_c_bits_address(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_address),.auto_tl_master_clock_xing_out_c_bits_data(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_data),.auto_tl_master_clock_xing_out_c_bits_corrupt(_tile_prci_domain_auto_tl_master_clock_xing_out_c_bits_corrupt),.auto_tl_master_clock_xing_out_d_ready(_tile_prci_domain_auto_tl_master_clock_xing_out_d_ready),.auto_tl_master_clock_xing_out_d_valid(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_valid),.auto_tl_master_clock_xing_out_d_bits_opcode(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_opcode),.auto_tl_master_clock_xing_out_d_bits_param(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_param),.auto_tl_master_clock_xing_out_d_bits_size(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_size),.auto_tl_master_clock_xing_out_d_bits_source(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_source),.auto_tl_master_clock_xing_out_d_bits_sink(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_sink),.auto_tl_master_clock_xing_out_d_bits_denied(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_denied),.auto_tl_master_clock_xing_out_d_bits_data(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_data),.auto_tl_master_clock_xing_out_d_bits_corrupt(_subsystem_sbus_auto_coupler_from_tile_tl_master_clock_xing_in_d_bits_corrupt),.auto_tl_master_clock_xing_out_e_valid(_tile_prci_domain_auto_tl_master_clock_xing_out_e_valid),.auto_tl_master_clock_xing_out_e_bits_sink(_tile_prci_domain_auto_tl_master_clock_xing_out_e_bits_sink),.auto_tap_clock_in_clock(_subsystem_sbus_auto_fixedClockNode_out_1_clock),.auto_tap_clock_in_reset(_subsystem_sbus_auto_fixedClockNode_out_1_reset)); 
  ClockSinkDomain plicDomainWrapper(.auto_plic_int_in_0(_ibus_int_bus_auto_int_out_0),.auto_plic_int_in_1(_ibus_int_bus_auto_int_out_1),.auto_plic_int_out_0(_plicDomainWrapper_auto_plic_int_out_0),.auto_plic_in_a_ready(_plicDomainWrapper_auto_plic_in_a_ready),.auto_plic_in_a_valid(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_valid),.auto_plic_in_a_bits_opcode(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_opcode),.auto_plic_in_a_bits_param(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_param),.auto_plic_in_a_bits_size(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_size),.auto_plic_in_a_bits_source(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_source),.auto_plic_in_a_bits_address(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_address),.auto_plic_in_a_bits_mask(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_mask),.auto_plic_in_a_bits_data(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_data),.auto_plic_in_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_a_bits_corrupt),.auto_plic_in_d_ready(_subsystem_cbus_auto_coupler_to_plic_fragmenter_out_d_ready),.auto_plic_in_d_valid(_plicDomainWrapper_auto_plic_in_d_valid),.auto_plic_in_d_bits_opcode(_plicDomainWrapper_auto_plic_in_d_bits_opcode),.auto_plic_in_d_bits_size(_plicDomainWrapper_auto_plic_in_d_bits_size),.auto_plic_in_d_bits_source(_plicDomainWrapper_auto_plic_in_d_bits_source),.auto_plic_in_d_bits_data(_plicDomainWrapper_auto_plic_in_d_bits_data),.auto_clock_in_clock(_subsystem_cbus_auto_fixedClockNode_out_0_clock),.auto_clock_in_reset(_subsystem_cbus_auto_fixedClockNode_out_0_reset)); 
  CLINT clint(.clock(_subsystem_cbus_clock),.reset(_subsystem_cbus_reset),.auto_int_out_0(_clint_auto_int_out_0),.auto_int_out_1(_clint_auto_int_out_1),.auto_in_a_ready(_clint_auto_in_a_ready),.auto_in_a_valid(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_valid),.auto_in_a_bits_opcode(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_opcode),.auto_in_a_bits_param(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_param),.auto_in_a_bits_size(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_size),.auto_in_a_bits_source(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_source),.auto_in_a_bits_address(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_address),.auto_in_a_bits_mask(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_mask),.auto_in_a_bits_data(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_data),.auto_in_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_a_bits_corrupt),.auto_in_d_ready(_subsystem_cbus_auto_coupler_to_clint_fragmenter_out_d_ready),.auto_in_d_valid(_clint_auto_in_d_valid),.auto_in_d_bits_opcode(_clint_auto_in_d_bits_opcode),.auto_in_d_bits_size(_clint_auto_in_d_bits_size),.auto_in_d_bits_source(_clint_auto_in_d_bits_source),.auto_in_d_bits_data(_clint_auto_in_d_bits_data),.io_rtcTick(int_rtc_tick)); 
  BundleBridgeNexus_15 tileHartIdNexusNode(.auto_out(_tileHartIdNexusNode_auto_out)); 
  TLDebugModule tlDM(.auto_dmInner_dmInner_tl_in_a_ready(_tlDM_auto_dmInner_dmInner_tl_in_a_ready),.auto_dmInner_dmInner_tl_in_a_valid(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_valid),.auto_dmInner_dmInner_tl_in_a_bits_opcode(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_opcode),.auto_dmInner_dmInner_tl_in_a_bits_param(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_param),.auto_dmInner_dmInner_tl_in_a_bits_size(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_size),.auto_dmInner_dmInner_tl_in_a_bits_source(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_source),.auto_dmInner_dmInner_tl_in_a_bits_address(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_address),.auto_dmInner_dmInner_tl_in_a_bits_mask(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_mask),.auto_dmInner_dmInner_tl_in_a_bits_data(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_data),.auto_dmInner_dmInner_tl_in_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_a_bits_corrupt),.auto_dmInner_dmInner_tl_in_d_ready(_subsystem_cbus_auto_coupler_to_debug_fragmenter_out_d_ready),.auto_dmInner_dmInner_tl_in_d_valid(_tlDM_auto_dmInner_dmInner_tl_in_d_valid),.auto_dmInner_dmInner_tl_in_d_bits_opcode(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_opcode),.auto_dmInner_dmInner_tl_in_d_bits_size(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_size),.auto_dmInner_dmInner_tl_in_d_bits_source(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_source),.auto_dmInner_dmInner_tl_in_d_bits_data(_tlDM_auto_dmInner_dmInner_tl_in_d_bits_data),.auto_dmOuter_intsource_out_sync_0(_tlDM_auto_dmOuter_intsource_out_sync_0),.io_debug_clock(debug_clock),.io_debug_reset(debug_reset),.io_ctrl_ndreset(debug_ndreset),.io_ctrl_dmactive(debug_dmactive),.io_ctrl_dmactiveAck(debug_dmactiveAck),.io_dmi_dmi_req_ready(debug_clockeddmi_dmi_req_ready),.io_dmi_dmi_req_valid(debug_clockeddmi_dmi_req_valid),.io_dmi_dmi_req_bits_addr(debug_clockeddmi_dmi_req_bits_addr),.io_dmi_dmi_req_bits_data(debug_clockeddmi_dmi_req_bits_data),.io_dmi_dmi_req_bits_op(debug_clockeddmi_dmi_req_bits_op),.io_dmi_dmi_resp_ready(debug_clockeddmi_dmi_resp_ready),.io_dmi_dmi_resp_valid(debug_clockeddmi_dmi_resp_valid),.io_dmi_dmi_resp_bits_data(debug_clockeddmi_dmi_resp_bits_data),.io_dmi_dmi_resp_bits_resp(debug_clockeddmi_dmi_resp_bits_resp),.io_dmi_dmiClock(debug_clockeddmi_dmiClock),.io_dmi_dmiReset(debug_clockeddmi_dmiReset),.io_hartIsInReset_0(resetctrl_hartIsInReset_0)); 
  IntSyncCrossingSource_5 intsource(.clock(clock),.reset(reset),.auto_in_0(_clint_auto_int_out_0),.auto_in_1(_clint_auto_int_out_1),.auto_out_sync_0(_intsource_auto_out_sync_0),.auto_out_sync_1(_intsource_auto_out_sync_1)); 
  IntSyncCrossingSource_1 intsource_1(.clock(clock),.reset(reset),.auto_in_0(_plicDomainWrapper_auto_plic_int_out_0),.auto_out_sync_0(_intsource_1_auto_out_sync_0)); 
  IntSyncCrossingSource_5 intsource_2(.clock(clock),.reset(reset),.auto_in_0(interrupts[0]),.auto_in_1(interrupts[1]),.auto_out_sync_0(_intsource_2_auto_out_sync_0),.auto_out_sync_1(_intsource_2_auto_out_sync_1)); 
  ClockSinkDomain_1 bootROMDomainWrapper(.auto_bootrom_in_a_ready(_bootROMDomainWrapper_auto_bootrom_in_a_ready),.auto_bootrom_in_a_valid(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_valid),.auto_bootrom_in_a_bits_opcode(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_opcode),.auto_bootrom_in_a_bits_param(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_param),.auto_bootrom_in_a_bits_size(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_size),.auto_bootrom_in_a_bits_source(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_source),.auto_bootrom_in_a_bits_address(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_address),.auto_bootrom_in_a_bits_mask(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_mask),.auto_bootrom_in_a_bits_corrupt(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_a_bits_corrupt),.auto_bootrom_in_d_ready(_subsystem_cbus_auto_coupler_to_bootrom_fragmenter_out_d_ready),.auto_bootrom_in_d_valid(_bootROMDomainWrapper_auto_bootrom_in_d_valid),.auto_bootrom_in_d_bits_size(_bootROMDomainWrapper_auto_bootrom_in_d_bits_size),.auto_bootrom_in_d_bits_source(_bootROMDomainWrapper_auto_bootrom_in_d_bits_source),.auto_bootrom_in_d_bits_data(_bootROMDomainWrapper_auto_bootrom_in_d_bits_data),.auto_clock_in_clock(_subsystem_cbus_auto_fixedClockNode_out_2_clock),.auto_clock_in_reset(_subsystem_cbus_auto_fixedClockNode_out_2_reset)); 
  assign mem_axi4_0_aw_bits_burst=2'h1; 
  assign mem_axi4_0_aw_bits_lock=1'h0; 
  assign mem_axi4_0_aw_bits_cache=4'h0; 
  assign mem_axi4_0_aw_bits_prot=3'h2; 
  assign mem_axi4_0_aw_bits_qos=4'h0; 
  assign mem_axi4_0_ar_bits_burst=2'h1; 
  assign mem_axi4_0_ar_bits_lock=1'h0; 
  assign mem_axi4_0_ar_bits_cache=4'h0; 
  assign mem_axi4_0_ar_bits_prot=3'h2; 
  assign mem_axi4_0_ar_bits_qos=4'h0; 
endmodule
 
module mem_33554432x64 (
  input [24:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [63:0] R0_data,
  input [24:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [63:0] W0_data,
  input [7:0] W0_mask) ; 
   reg [63:0] Memory[0:33554431] ;  
   reg _R0_en_d0 ;  
   reg [24:0] _R0_addr_d0 ;  
  always @( posedge R0_clk)
       begin 
         _R0_en_d0 <=R0_en;
         _R0_addr_d0 <=R0_addr;
       end
  
  always @( posedge W0_clk)
       begin 
         if (W0_en&W0_mask[0])
            Memory [W0_addr][32'h0+:8]<=W0_data[7:0];
         if (W0_en&W0_mask[1])
            Memory [W0_addr][32'h8+:8]<=W0_data[15:8];
         if (W0_en&W0_mask[2])
            Memory [W0_addr][32'h10+:8]<=W0_data[23:16];
         if (W0_en&W0_mask[3])
            Memory [W0_addr][32'h18+:8]<=W0_data[31:24];
         if (W0_en&W0_mask[4])
            Memory [W0_addr][32'h20+:8]<=W0_data[39:32];
         if (W0_en&W0_mask[5])
            Memory [W0_addr][32'h28+:8]<=W0_data[47:40];
         if (W0_en&W0_mask[6])
            Memory [W0_addr][32'h30+:8]<=W0_data[55:48];
         if (W0_en&W0_mask[7])
            Memory [W0_addr][32'h38+:8]<=W0_data[63:56];
       end
  
  assign R0_data=_R0_en_d0 ? Memory[_R0_addr_d0]:64'bx; 
endmodule
 
module AXI4RAM (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input auto_in_aw_bits_echo_real_last,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_b_bits_echo_real_last,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input auto_in_ar_bits_echo_real_last,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_echo_real_last) ; 
   wire nodeIn_ar_ready ;  
   wire nodeIn_aw_ready ;  
   wire [63:0] _mem_ext_R0_data ;  
   wire w_sel0=auto_in_aw_bits_addr[31:28]==4'h8 ;  
   reg w_full ;  
   reg [3:0] w_id ;  
   reg w_echo_real_last ;  
   reg r_sel1 ;  
   reg w_sel1 ;  
   wire _GEN=nodeIn_aw_ready&auto_in_aw_valid ;  
  assign nodeIn_aw_ready=auto_in_w_valid&(auto_in_b_ready|~w_full); 
   reg r_full ;  
   reg [3:0] r_id ;  
   reg r_echo_real_last ;  
   wire ren=nodeIn_ar_ready&auto_in_ar_valid ;  
   reg rdata_REG ;  
   reg [7:0] rdata_r_0 ;  
   reg [7:0] rdata_r_1 ;  
   reg [7:0] rdata_r_2 ;  
   reg [7:0] rdata_r_3 ;  
   reg [7:0] rdata_r_4 ;  
   reg [7:0] rdata_r_5 ;  
   reg [7:0] rdata_r_6 ;  
   reg [7:0] rdata_r_7 ;  
  assign nodeIn_ar_ready=auto_in_r_ready|~r_full; 
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              w_full <=1'h0;
              r_full <=1'h0;
            end 
          else 
            begin 
              w_full <=_GEN|~(auto_in_b_ready&w_full)&w_full;
              r_full <=ren|~(auto_in_r_ready&r_full)&r_full;
            end 
         if (_GEN)
            begin 
              w_id <=auto_in_aw_bits_id;
              w_echo_real_last <=auto_in_aw_bits_echo_real_last;
            end 
         r_sel1 <=auto_in_ar_bits_addr[31:28]==4'h8;
         w_sel1 <=w_sel0;
         if (ren)
            begin 
              r_id <=auto_in_ar_bits_id;
              r_echo_real_last <=auto_in_ar_bits_echo_real_last;
            end 
         rdata_REG <=ren;
         if (rdata_REG)
            begin 
              rdata_r_0 <=_mem_ext_R0_data[7:0];
              rdata_r_1 <=_mem_ext_R0_data[15:8];
              rdata_r_2 <=_mem_ext_R0_data[23:16];
              rdata_r_3 <=_mem_ext_R0_data[31:24];
              rdata_r_4 <=_mem_ext_R0_data[39:32];
              rdata_r_5 <=_mem_ext_R0_data[47:40];
              rdata_r_6 <=_mem_ext_R0_data[55:48];
              rdata_r_7 <=_mem_ext_R0_data[63:56];
            end 
       end
  
  mem_33554432x64 mem_ext(.R0_addr(auto_in_ar_bits_addr[27:3]),.R0_en(ren),.R0_clk(clock),.R0_data(_mem_ext_R0_data),.W0_addr(auto_in_aw_bits_addr[27:3]),.W0_en(_GEN&w_sel0),.W0_clk(clock),.W0_data(auto_in_w_bits_data),.W0_mask(auto_in_w_bits_strb)); 
  assign auto_in_aw_ready=nodeIn_aw_ready; 
  assign auto_in_w_ready=auto_in_aw_valid&(auto_in_b_ready|~w_full); 
  assign auto_in_b_valid=w_full; 
  assign auto_in_b_bits_id=w_id; 
  assign auto_in_b_bits_resp=w_sel1 ? 2'h0:2'h3; 
  assign auto_in_b_bits_echo_real_last=w_echo_real_last; 
  assign auto_in_ar_ready=nodeIn_ar_ready; 
  assign auto_in_r_valid=r_full; 
  assign auto_in_r_bits_id=r_id; 
  assign auto_in_r_bits_data={rdata_REG ? _mem_ext_R0_data[63:56]:rdata_r_7,rdata_REG ? _mem_ext_R0_data[55:48]:rdata_r_6,rdata_REG ? _mem_ext_R0_data[47:40]:rdata_r_5,rdata_REG ? _mem_ext_R0_data[39:32]:rdata_r_4,rdata_REG ? _mem_ext_R0_data[31:24]:rdata_r_3,rdata_REG ? _mem_ext_R0_data[23:16]:rdata_r_2,rdata_REG ? _mem_ext_R0_data[15:8]:rdata_r_1,rdata_REG ? _mem_ext_R0_data[7:0]:rdata_r_0}; 
  assign auto_in_r_bits_resp=r_sel1 ? 2'h0:2'h3; 
  assign auto_in_r_bits_echo_real_last=r_echo_real_last; 
endmodule
 
module AXI4Xbar (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [1:0] auto_in_aw_bits_burst,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [1:0] auto_in_ar_bits_burst,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [1:0] auto_out_aw_bits_burst,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [1:0] auto_out_ar_bits_burst,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_last) ; 
  assign auto_in_aw_ready=auto_out_aw_ready; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_ar_ready=auto_out_ar_ready; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_aw_bits_burst=auto_in_aw_bits_burst; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_ar_bits_burst=auto_in_ar_bits_burst; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module Queue_86 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [31:0] io_enq_bits_addr,
  input io_enq_bits_echo_real_last,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output io_deq_bits_echo_real_last) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x4 ram_id_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_addr_2x32 ram_addr_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_addr),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_addr)); 
  ram_2x1 ram_echo_real_last_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_echo_real_last),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_echo_real_last)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_88 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [1:0] io_enq_bits_resp,
  input io_enq_bits_echo_real_last,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp,
  output io_deq_bits_echo_real_last) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x4 ram_id_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_2x2 ram_resp_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_resp),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_resp)); 
  ram_2x1 ram_echo_real_last_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_echo_real_last),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_echo_real_last)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module Queue_90 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [63:0] io_enq_bits_data,
  input [1:0] io_enq_bits_resp,
  input io_enq_bits_echo_real_last,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0] io_deq_bits_resp,
  output io_deq_bits_echo_real_last,
  output io_deq_bits_last) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x4 ram_id_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_data_2x64 ram_data_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_data),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_data)); 
  ram_2x2 ram_resp_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_resp),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_resp)); 
  ram_2x1 ram_echo_real_last_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_echo_real_last),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_echo_real_last)); 
  ram_2x1 ram_last_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_last),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(1'h1)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module AXI4Buffer_1 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input auto_in_aw_bits_echo_real_last,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_b_bits_echo_real_last,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input auto_in_ar_bits_echo_real_last,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_echo_real_last,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output auto_out_aw_bits_echo_real_last,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_b_bits_echo_real_last,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output auto_out_ar_bits_echo_real_last,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_echo_real_last) ; 
  Queue_86 nodeOut_aw_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_aw_ready),.io_enq_valid(auto_in_aw_valid),.io_enq_bits_id(auto_in_aw_bits_id),.io_enq_bits_addr(auto_in_aw_bits_addr),.io_enq_bits_echo_real_last(auto_in_aw_bits_echo_real_last),.io_deq_ready(auto_out_aw_ready),.io_deq_valid(auto_out_aw_valid),.io_deq_bits_id(auto_out_aw_bits_id),.io_deq_bits_addr(auto_out_aw_bits_addr),.io_deq_bits_echo_real_last(auto_out_aw_bits_echo_real_last)); 
  Queue_1 nodeOut_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_w_ready),.io_enq_valid(auto_in_w_valid),.io_enq_bits_data(auto_in_w_bits_data),.io_enq_bits_strb(auto_in_w_bits_strb),.io_enq_bits_last(auto_in_w_bits_last),.io_deq_ready(auto_out_w_ready),.io_deq_valid(auto_out_w_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last()); 
  Queue_88 nodeIn_b_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_b_ready),.io_enq_valid(auto_out_b_valid),.io_enq_bits_id(auto_out_b_bits_id),.io_enq_bits_resp(auto_out_b_bits_resp),.io_enq_bits_echo_real_last(auto_out_b_bits_echo_real_last),.io_deq_ready(auto_in_b_ready),.io_deq_valid(auto_in_b_valid),.io_deq_bits_id(auto_in_b_bits_id),.io_deq_bits_resp(auto_in_b_bits_resp),.io_deq_bits_echo_real_last(auto_in_b_bits_echo_real_last)); 
  Queue_86 nodeOut_ar_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_ar_ready),.io_enq_valid(auto_in_ar_valid),.io_enq_bits_id(auto_in_ar_bits_id),.io_enq_bits_addr(auto_in_ar_bits_addr),.io_enq_bits_echo_real_last(auto_in_ar_bits_echo_real_last),.io_deq_ready(auto_out_ar_ready),.io_deq_valid(auto_out_ar_valid),.io_deq_bits_id(auto_out_ar_bits_id),.io_deq_bits_addr(auto_out_ar_bits_addr),.io_deq_bits_echo_real_last(auto_out_ar_bits_echo_real_last)); 
  Queue_90 nodeIn_r_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_r_ready),.io_enq_valid(auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_echo_real_last(auto_out_r_bits_echo_real_last),.io_deq_ready(auto_in_r_ready),.io_deq_valid(auto_in_r_valid),.io_deq_bits_id(auto_in_r_bits_id),.io_deq_bits_data(auto_in_r_bits_data),.io_deq_bits_resp(auto_in_r_bits_resp),.io_deq_bits_echo_real_last(auto_in_r_bits_echo_real_last),.io_deq_bits_last(auto_in_r_bits_last)); 
endmodule
 
module Queue_91 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [31:0] io_enq_bits_addr,
  input [7:0] io_enq_bits_len,
  input [2:0] io_enq_bits_size,
  input [1:0] io_enq_bits_burst,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst) ; 
   reg [1:0] ram_burst ;  
   reg [2:0] ram_size ;  
   reg [7:0] ram_len ;  
   reg [31:0] ram_addr ;  
   reg [3:0] ram_id ;  
   reg full ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire do_enq=~(~full&io_deq_ready)&~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_burst <=io_enq_bits_burst;
              ram_size <=io_enq_bits_size;
              ram_len <=io_enq_bits_len;
              ram_addr <=io_enq_bits_addr;
              ram_id <=io_enq_bits_id;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(full&io_deq_ready&io_deq_valid_0)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_id=full ? ram_id:io_enq_bits_id; 
  assign io_deq_bits_addr=full ? ram_addr:io_enq_bits_addr; 
  assign io_deq_bits_len=full ? ram_len:io_enq_bits_len; 
  assign io_deq_bits_size=full ? ram_size:io_enq_bits_size; 
  assign io_deq_bits_burst=full ? ram_burst:io_enq_bits_burst; 
endmodule
 
module AXI4Fragmenter_1 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [31:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [1:0] auto_in_aw_bits_burst,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [31:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [1:0] auto_in_ar_bits_burst,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output auto_out_aw_bits_echo_real_last,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_b_bits_echo_real_last,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output auto_out_ar_bits_echo_real_last,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_echo_real_last,
  input auto_out_r_bits_last) ; 
   wire nodeOut_w_valid ;  
   wire w_idle ;  
   wire in_aw_ready ;  
   wire _in_w_deq_q_io_deq_valid ;  
   wire _in_w_deq_q_io_deq_bits_last ;  
   wire _deq_q_1_io_deq_valid ;  
   wire [31:0] _deq_q_1_io_deq_bits_addr ;  
   wire [7:0] _deq_q_1_io_deq_bits_len ;  
   wire [2:0] _deq_q_1_io_deq_bits_size ;  
   wire [1:0] _deq_q_1_io_deq_bits_burst ;  
   wire _deq_q_io_deq_valid ;  
   wire [31:0] _deq_q_io_deq_bits_addr ;  
   wire [7:0] _deq_q_io_deq_bits_len ;  
   wire [2:0] _deq_q_io_deq_bits_size ;  
   wire [1:0] _deq_q_io_deq_bits_burst ;  
   reg busy ;  
   reg [31:0] r_addr ;  
   reg [7:0] r_len ;  
   wire [7:0] len=busy ? r_len:_deq_q_io_deq_bits_len ;  
   wire [31:0] addr=busy ? r_addr:_deq_q_io_deq_bits_addr ;  
   wire [31:0] _out_bits_addr_T=~addr ;  
   wire [9:0] _out_bits_addr_T_2=10'h7<<_deq_q_io_deq_bits_size ;  
   reg busy_1 ;  
   reg [31:0] r_addr_1 ;  
   reg [7:0] r_len_1 ;  
   wire [7:0] len_1=busy_1 ? r_len_1:_deq_q_1_io_deq_bits_len ;  
   wire [31:0] addr_1=busy_1 ? r_addr_1:_deq_q_1_io_deq_bits_addr ;  
   wire [31:0] _out_bits_addr_T_7=~addr_1 ;  
   wire [9:0] _out_bits_addr_T_9=10'h7<<_deq_q_1_io_deq_bits_size ;  
   reg wbeats_latched ;  
   wire _in_aw_ready_T=w_idle|wbeats_latched ;  
   wire nodeOut_aw_valid=_deq_q_1_io_deq_valid&_in_aw_ready_T ;  
  assign in_aw_ready=auto_out_aw_ready&_in_aw_ready_T; 
   wire wbeats_valid=_deq_q_1_io_deq_valid&~wbeats_latched ;  
   reg [8:0] w_counter ;  
  assign w_idle=w_counter==9'h0; 
   wire [8:0] w_todo=w_idle ? {8'h0,wbeats_valid}:w_counter ;  
   wire w_last=w_todo==9'h1 ;  
   wire _w_counter_T=auto_out_w_ready&nodeOut_w_valid ;  
  assign nodeOut_w_valid=_in_w_deq_q_io_deq_valid&(~w_idle|wbeats_valid); 
  always @( posedge clock)
       begin 
         if (~reset&~(~_w_counter_T|(|w_todo)))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:177 assert (!out.w.fire || w_todo =/= 0.U) // underflow impossible\n");
              if (1)$display("");
            end 
         if (~reset&~(~nodeOut_w_valid|~_in_w_deq_q_io_deq_bits_last|w_last))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:186 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
              if (1)$display("");
            end 
       end
  
   wire nodeOut_b_ready=auto_in_b_ready|~auto_out_b_bits_echo_real_last ;  
   reg [1:0] error_0 ;  
   reg [1:0] error_1 ;  
   reg [1:0] error_2 ;  
   reg [1:0] error_3 ;  
   reg [1:0] error_4 ;  
   reg [1:0] error_5 ;  
   reg [1:0] error_6 ;  
   reg [1:0] error_7 ;  
   reg [1:0] error_8 ;  
   reg [1:0] error_9 ;  
   reg [1:0] error_10 ;  
   reg [1:0] error_11 ;  
   reg [1:0] error_12 ;  
   reg [1:0] error_13 ;  
   reg [1:0] error_14 ;  
   reg [1:0] error_15 ;  
   reg [1:0] casez_tmp ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp =error_0;
          4 'b0001:
             casez_tmp =error_1;
          4 'b0010:
             casez_tmp =error_2;
          4 'b0011:
             casez_tmp =error_3;
          4 'b0100:
             casez_tmp =error_4;
          4 'b0101:
             casez_tmp =error_5;
          4 'b0110:
             casez_tmp =error_6;
          4 'b0111:
             casez_tmp =error_7;
          4 'b1000:
             casez_tmp =error_8;
          4 'b1001:
             casez_tmp =error_9;
          4 'b1010:
             casez_tmp =error_10;
          4 'b1011:
             casez_tmp =error_11;
          4 'b1100:
             casez_tmp =error_12;
          4 'b1101:
             casez_tmp =error_13;
          4 'b1110:
             casez_tmp =error_14;
          default :
             casez_tmp =error_15;
         endcase 
       end
  
   wire _GEN=nodeOut_b_ready&auto_out_b_valid ;  
   wire [22:0] _wrapMask_T_1={7'h0,_deq_q_io_deq_bits_len,8'hFF}<<_deq_q_io_deq_bits_size ;  
   wire [31:0] _mux_addr_T_1=~_deq_q_io_deq_bits_addr ;  
   wire [31:0] _inc_addr_T_1=addr+{16'h0,16'h1<<_deq_q_io_deq_bits_size} ;  
   wire [22:0] _wrapMask_T_3={7'h0,_deq_q_1_io_deq_bits_len,8'hFF}<<_deq_q_1_io_deq_bits_size ;  
   wire [31:0] _mux_addr_T_6=~_deq_q_1_io_deq_bits_addr ;  
   wire [31:0] _inc_addr_T_3=addr_1+{16'h0,16'h1<<_deq_q_1_io_deq_bits_size} ;  
   wire _GEN_0=auto_out_ar_ready&_deq_q_io_deq_valid ;  
   wire _GEN_1=in_aw_ready&_deq_q_1_io_deq_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              busy <=1'h0;
              busy_1 <=1'h0;
              wbeats_latched <=1'h0;
              w_counter <=9'h0;
              error_0 <=2'h0;
              error_1 <=2'h0;
              error_2 <=2'h0;
              error_3 <=2'h0;
              error_4 <=2'h0;
              error_5 <=2'h0;
              error_6 <=2'h0;
              error_7 <=2'h0;
              error_8 <=2'h0;
              error_9 <=2'h0;
              error_10 <=2'h0;
              error_11 <=2'h0;
              error_12 <=2'h0;
              error_13 <=2'h0;
              error_14 <=2'h0;
              error_15 <=2'h0;
            end 
          else 
            begin 
              if (_GEN_0)
                 busy <=|len;
              if (_GEN_1)
                 busy_1 <=|len_1;
              wbeats_latched <=~(auto_out_aw_ready&nodeOut_aw_valid)&(wbeats_valid&w_idle|wbeats_latched);
              w_counter <=w_todo-{8'h0,_w_counter_T};
              if (auto_out_b_bits_id==4'h0&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_0 <=2'h0;
                    else 
                      error_0 <=error_0|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h1&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_1 <=2'h0;
                    else 
                      error_1 <=error_1|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h2&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_2 <=2'h0;
                    else 
                      error_2 <=error_2|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h3&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_3 <=2'h0;
                    else 
                      error_3 <=error_3|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h4&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_4 <=2'h0;
                    else 
                      error_4 <=error_4|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h5&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_5 <=2'h0;
                    else 
                      error_5 <=error_5|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h6&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_6 <=2'h0;
                    else 
                      error_6 <=error_6|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h7&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_7 <=2'h0;
                    else 
                      error_7 <=error_7|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h8&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_8 <=2'h0;
                    else 
                      error_8 <=error_8|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h9&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_9 <=2'h0;
                    else 
                      error_9 <=error_9|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hA&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_10 <=2'h0;
                    else 
                      error_10 <=error_10|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hB&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_11 <=2'h0;
                    else 
                      error_11 <=error_11|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hC&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_12 <=2'h0;
                    else 
                      error_12 <=error_12|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hD&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_13 <=2'h0;
                    else 
                      error_13 <=error_13|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hE&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_14 <=2'h0;
                    else 
                      error_14 <=error_14|auto_out_b_bits_resp;
                 end 
              if ((&auto_out_b_bits_id)&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_15 <=2'h0;
                    else 
                      error_15 <=error_15|auto_out_b_bits_resp;
                 end 
            end 
         if (_GEN_0)
            begin 
              if (_deq_q_io_deq_bits_burst==2'h0)
                 r_addr <=_deq_q_io_deq_bits_addr;
               else 
                 if (_deq_q_io_deq_bits_burst==2'h2)
                    r_addr <={17'h0,_inc_addr_T_1[14:0]&_wrapMask_T_1[22:8]}|~{_mux_addr_T_1[31:15],_mux_addr_T_1[14:0]|_wrapMask_T_1[22:8]};
                  else 
                    r_addr <=_inc_addr_T_1;
              r_len <=len-8'h1;
            end 
         if (_GEN_1)
            begin 
              if (_deq_q_1_io_deq_bits_burst==2'h0)
                 r_addr_1 <=_deq_q_1_io_deq_bits_addr;
               else 
                 if (_deq_q_1_io_deq_bits_burst==2'h2)
                    r_addr_1 <={17'h0,_inc_addr_T_3[14:0]&_wrapMask_T_3[22:8]}|~{_mux_addr_T_6[31:15],_mux_addr_T_6[14:0]|_wrapMask_T_3[22:8]};
                  else 
                    r_addr_1 <=_inc_addr_T_3;
              r_len_1 <=len_1-8'h1;
            end 
       end
  
  Queue_91 deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_ar_ready),.io_enq_valid(auto_in_ar_valid),.io_enq_bits_id(auto_in_ar_bits_id),.io_enq_bits_addr(auto_in_ar_bits_addr),.io_enq_bits_len(auto_in_ar_bits_len),.io_enq_bits_size(auto_in_ar_bits_size),.io_enq_bits_burst(auto_in_ar_bits_burst),.io_deq_ready(auto_out_ar_ready&~(|len)),.io_deq_valid(_deq_q_io_deq_valid),.io_deq_bits_id(auto_out_ar_bits_id),.io_deq_bits_addr(_deq_q_io_deq_bits_addr),.io_deq_bits_len(_deq_q_io_deq_bits_len),.io_deq_bits_size(_deq_q_io_deq_bits_size),.io_deq_bits_burst(_deq_q_io_deq_bits_burst)); 
  Queue_91 deq_q_1(.clock(clock),.reset(reset),.io_enq_ready(auto_in_aw_ready),.io_enq_valid(auto_in_aw_valid),.io_enq_bits_id(auto_in_aw_bits_id),.io_enq_bits_addr(auto_in_aw_bits_addr),.io_enq_bits_len(auto_in_aw_bits_len),.io_enq_bits_size(auto_in_aw_bits_size),.io_enq_bits_burst(auto_in_aw_bits_burst),.io_deq_ready(in_aw_ready&~(|len_1)),.io_deq_valid(_deq_q_1_io_deq_valid),.io_deq_bits_id(auto_out_aw_bits_id),.io_deq_bits_addr(_deq_q_1_io_deq_bits_addr),.io_deq_bits_len(_deq_q_1_io_deq_bits_len),.io_deq_bits_size(_deq_q_1_io_deq_bits_size),.io_deq_bits_burst(_deq_q_1_io_deq_bits_burst)); 
  Queue_34 in_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_w_ready),.io_enq_valid(auto_in_w_valid),.io_enq_bits_data(auto_in_w_bits_data),.io_enq_bits_strb(auto_in_w_bits_strb),.io_enq_bits_last(auto_in_w_bits_last),.io_deq_ready(auto_out_w_ready&(~w_idle|wbeats_valid)),.io_deq_valid(_in_w_deq_q_io_deq_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last(_in_w_deq_q_io_deq_bits_last)); 
  assign auto_in_b_valid=auto_out_b_valid&auto_out_b_bits_echo_real_last; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp|casez_tmp; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_last=auto_out_r_bits_last&auto_out_r_bits_echo_real_last; 
  assign auto_out_aw_valid=nodeOut_aw_valid; 
  assign auto_out_aw_bits_addr=~{_out_bits_addr_T_7[31:3],_out_bits_addr_T_7[2:0]|~(_out_bits_addr_T_9[2:0])}; 
  assign auto_out_aw_bits_echo_real_last=~(|len_1); 
  assign auto_out_w_valid=nodeOut_w_valid; 
  assign auto_out_w_bits_last=w_last; 
  assign auto_out_b_ready=nodeOut_b_ready; 
  assign auto_out_ar_valid=_deq_q_io_deq_valid; 
  assign auto_out_ar_bits_addr=~{_out_bits_addr_T[31:3],_out_bits_addr_T[2:0]|~(_out_bits_addr_T_2[2:0])}; 
  assign auto_out_ar_bits_echo_real_last=~(|len); 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module SimAXIMem (
  input clock,
  input reset,
  output io_axi4_0_aw_ready,
  input io_axi4_0_aw_valid,
  input [3:0] io_axi4_0_aw_bits_id,
  input [31:0] io_axi4_0_aw_bits_addr,
  input [7:0] io_axi4_0_aw_bits_len,
  input [2:0] io_axi4_0_aw_bits_size,
  input [1:0] io_axi4_0_aw_bits_burst,
  output io_axi4_0_w_ready,
  input io_axi4_0_w_valid,
  input [63:0] io_axi4_0_w_bits_data,
  input [7:0] io_axi4_0_w_bits_strb,
  input io_axi4_0_w_bits_last,
  input io_axi4_0_b_ready,
  output io_axi4_0_b_valid,
  output [3:0] io_axi4_0_b_bits_id,
  output [1:0] io_axi4_0_b_bits_resp,
  output io_axi4_0_ar_ready,
  input io_axi4_0_ar_valid,
  input [3:0] io_axi4_0_ar_bits_id,
  input [31:0] io_axi4_0_ar_bits_addr,
  input [7:0] io_axi4_0_ar_bits_len,
  input [2:0] io_axi4_0_ar_bits_size,
  input [1:0] io_axi4_0_ar_bits_burst,
  input io_axi4_0_r_ready,
  output io_axi4_0_r_valid,
  output [3:0] io_axi4_0_r_bits_id,
  output [63:0] io_axi4_0_r_bits_data,
  output [1:0] io_axi4_0_r_bits_resp,
  output io_axi4_0_r_bits_last) ; 
   wire _axi4frag_auto_in_aw_ready ;  
   wire _axi4frag_auto_in_w_ready ;  
   wire _axi4frag_auto_in_b_valid ;  
   wire [3:0] _axi4frag_auto_in_b_bits_id ;  
   wire [1:0] _axi4frag_auto_in_b_bits_resp ;  
   wire _axi4frag_auto_in_ar_ready ;  
   wire _axi4frag_auto_in_r_valid ;  
   wire [3:0] _axi4frag_auto_in_r_bits_id ;  
   wire [63:0] _axi4frag_auto_in_r_bits_data ;  
   wire [1:0] _axi4frag_auto_in_r_bits_resp ;  
   wire _axi4frag_auto_in_r_bits_last ;  
   wire _axi4frag_auto_out_aw_valid ;  
   wire [3:0] _axi4frag_auto_out_aw_bits_id ;  
   wire [31:0] _axi4frag_auto_out_aw_bits_addr ;  
   wire _axi4frag_auto_out_aw_bits_echo_real_last ;  
   wire _axi4frag_auto_out_w_valid ;  
   wire [63:0] _axi4frag_auto_out_w_bits_data ;  
   wire [7:0] _axi4frag_auto_out_w_bits_strb ;  
   wire _axi4frag_auto_out_w_bits_last ;  
   wire _axi4frag_auto_out_b_ready ;  
   wire _axi4frag_auto_out_ar_valid ;  
   wire [3:0] _axi4frag_auto_out_ar_bits_id ;  
   wire [31:0] _axi4frag_auto_out_ar_bits_addr ;  
   wire _axi4frag_auto_out_ar_bits_echo_real_last ;  
   wire _axi4frag_auto_out_r_ready ;  
   wire _axi4buf_auto_in_aw_ready ;  
   wire _axi4buf_auto_in_w_ready ;  
   wire _axi4buf_auto_in_b_valid ;  
   wire [3:0] _axi4buf_auto_in_b_bits_id ;  
   wire [1:0] _axi4buf_auto_in_b_bits_resp ;  
   wire _axi4buf_auto_in_b_bits_echo_real_last ;  
   wire _axi4buf_auto_in_ar_ready ;  
   wire _axi4buf_auto_in_r_valid ;  
   wire [3:0] _axi4buf_auto_in_r_bits_id ;  
   wire [63:0] _axi4buf_auto_in_r_bits_data ;  
   wire [1:0] _axi4buf_auto_in_r_bits_resp ;  
   wire _axi4buf_auto_in_r_bits_echo_real_last ;  
   wire _axi4buf_auto_in_r_bits_last ;  
   wire _axi4buf_auto_out_aw_valid ;  
   wire [3:0] _axi4buf_auto_out_aw_bits_id ;  
   wire [31:0] _axi4buf_auto_out_aw_bits_addr ;  
   wire _axi4buf_auto_out_aw_bits_echo_real_last ;  
   wire _axi4buf_auto_out_w_valid ;  
   wire [63:0] _axi4buf_auto_out_w_bits_data ;  
   wire [7:0] _axi4buf_auto_out_w_bits_strb ;  
   wire _axi4buf_auto_out_b_ready ;  
   wire _axi4buf_auto_out_ar_valid ;  
   wire [3:0] _axi4buf_auto_out_ar_bits_id ;  
   wire [31:0] _axi4buf_auto_out_ar_bits_addr ;  
   wire _axi4buf_auto_out_ar_bits_echo_real_last ;  
   wire _axi4buf_auto_out_r_ready ;  
   wire _axi4xbar_auto_out_aw_valid ;  
   wire [3:0] _axi4xbar_auto_out_aw_bits_id ;  
   wire [31:0] _axi4xbar_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4xbar_auto_out_aw_bits_len ;  
   wire [2:0] _axi4xbar_auto_out_aw_bits_size ;  
   wire [1:0] _axi4xbar_auto_out_aw_bits_burst ;  
   wire _axi4xbar_auto_out_w_valid ;  
   wire [63:0] _axi4xbar_auto_out_w_bits_data ;  
   wire [7:0] _axi4xbar_auto_out_w_bits_strb ;  
   wire _axi4xbar_auto_out_w_bits_last ;  
   wire _axi4xbar_auto_out_b_ready ;  
   wire _axi4xbar_auto_out_ar_valid ;  
   wire [3:0] _axi4xbar_auto_out_ar_bits_id ;  
   wire [31:0] _axi4xbar_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4xbar_auto_out_ar_bits_len ;  
   wire [2:0] _axi4xbar_auto_out_ar_bits_size ;  
   wire [1:0] _axi4xbar_auto_out_ar_bits_burst ;  
   wire _axi4xbar_auto_out_r_ready ;  
   wire _srams_auto_in_aw_ready ;  
   wire _srams_auto_in_w_ready ;  
   wire _srams_auto_in_b_valid ;  
   wire [3:0] _srams_auto_in_b_bits_id ;  
   wire [1:0] _srams_auto_in_b_bits_resp ;  
   wire _srams_auto_in_b_bits_echo_real_last ;  
   wire _srams_auto_in_ar_ready ;  
   wire _srams_auto_in_r_valid ;  
   wire [3:0] _srams_auto_in_r_bits_id ;  
   wire [63:0] _srams_auto_in_r_bits_data ;  
   wire [1:0] _srams_auto_in_r_bits_resp ;  
   wire _srams_auto_in_r_bits_echo_real_last ;  
  AXI4RAM srams(.clock(clock),.reset(reset),.auto_in_aw_ready(_srams_auto_in_aw_ready),.auto_in_aw_valid(_axi4buf_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4buf_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4buf_auto_out_aw_bits_addr),.auto_in_aw_bits_echo_real_last(_axi4buf_auto_out_aw_bits_echo_real_last),.auto_in_w_ready(_srams_auto_in_w_ready),.auto_in_w_valid(_axi4buf_auto_out_w_valid),.auto_in_w_bits_data(_axi4buf_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4buf_auto_out_w_bits_strb),.auto_in_b_ready(_axi4buf_auto_out_b_ready),.auto_in_b_valid(_srams_auto_in_b_valid),.auto_in_b_bits_id(_srams_auto_in_b_bits_id),.auto_in_b_bits_resp(_srams_auto_in_b_bits_resp),.auto_in_b_bits_echo_real_last(_srams_auto_in_b_bits_echo_real_last),.auto_in_ar_ready(_srams_auto_in_ar_ready),.auto_in_ar_valid(_axi4buf_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4buf_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4buf_auto_out_ar_bits_addr),.auto_in_ar_bits_echo_real_last(_axi4buf_auto_out_ar_bits_echo_real_last),.auto_in_r_ready(_axi4buf_auto_out_r_ready),.auto_in_r_valid(_srams_auto_in_r_valid),.auto_in_r_bits_id(_srams_auto_in_r_bits_id),.auto_in_r_bits_data(_srams_auto_in_r_bits_data),.auto_in_r_bits_resp(_srams_auto_in_r_bits_resp),.auto_in_r_bits_echo_real_last(_srams_auto_in_r_bits_echo_real_last)); 
  AXI4Xbar axi4xbar(.clock(clock),.reset(reset),.auto_in_aw_ready(io_axi4_0_aw_ready),.auto_in_aw_valid(io_axi4_0_aw_valid),.auto_in_aw_bits_id(io_axi4_0_aw_bits_id),.auto_in_aw_bits_addr(io_axi4_0_aw_bits_addr),.auto_in_aw_bits_len(io_axi4_0_aw_bits_len),.auto_in_aw_bits_size(io_axi4_0_aw_bits_size),.auto_in_aw_bits_burst(io_axi4_0_aw_bits_burst),.auto_in_w_ready(io_axi4_0_w_ready),.auto_in_w_valid(io_axi4_0_w_valid),.auto_in_w_bits_data(io_axi4_0_w_bits_data),.auto_in_w_bits_strb(io_axi4_0_w_bits_strb),.auto_in_w_bits_last(io_axi4_0_w_bits_last),.auto_in_b_ready(io_axi4_0_b_ready),.auto_in_b_valid(io_axi4_0_b_valid),.auto_in_b_bits_id(io_axi4_0_b_bits_id),.auto_in_b_bits_resp(io_axi4_0_b_bits_resp),.auto_in_ar_ready(io_axi4_0_ar_ready),.auto_in_ar_valid(io_axi4_0_ar_valid),.auto_in_ar_bits_id(io_axi4_0_ar_bits_id),.auto_in_ar_bits_addr(io_axi4_0_ar_bits_addr),.auto_in_ar_bits_len(io_axi4_0_ar_bits_len),.auto_in_ar_bits_size(io_axi4_0_ar_bits_size),.auto_in_ar_bits_burst(io_axi4_0_ar_bits_burst),.auto_in_r_ready(io_axi4_0_r_ready),.auto_in_r_valid(io_axi4_0_r_valid),.auto_in_r_bits_id(io_axi4_0_r_bits_id),.auto_in_r_bits_data(io_axi4_0_r_bits_data),.auto_in_r_bits_resp(io_axi4_0_r_bits_resp),.auto_in_r_bits_last(io_axi4_0_r_bits_last),.auto_out_aw_ready(_axi4frag_auto_in_aw_ready),.auto_out_aw_valid(_axi4xbar_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4xbar_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4xbar_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4xbar_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4xbar_auto_out_aw_bits_size),.auto_out_aw_bits_burst(_axi4xbar_auto_out_aw_bits_burst),.auto_out_w_ready(_axi4frag_auto_in_w_ready),.auto_out_w_valid(_axi4xbar_auto_out_w_valid),.auto_out_w_bits_data(_axi4xbar_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4xbar_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4xbar_auto_out_w_bits_last),.auto_out_b_ready(_axi4xbar_auto_out_b_ready),.auto_out_b_valid(_axi4frag_auto_in_b_valid),.auto_out_b_bits_id(_axi4frag_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4frag_auto_in_b_bits_resp),.auto_out_ar_ready(_axi4frag_auto_in_ar_ready),.auto_out_ar_valid(_axi4xbar_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4xbar_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4xbar_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4xbar_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4xbar_auto_out_ar_bits_size),.auto_out_ar_bits_burst(_axi4xbar_auto_out_ar_bits_burst),.auto_out_r_ready(_axi4xbar_auto_out_r_ready),.auto_out_r_valid(_axi4frag_auto_in_r_valid),.auto_out_r_bits_id(_axi4frag_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4frag_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4frag_auto_in_r_bits_resp),.auto_out_r_bits_last(_axi4frag_auto_in_r_bits_last)); 
  AXI4Buffer_1 axi4buf(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4buf_auto_in_aw_ready),.auto_in_aw_valid(_axi4frag_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4frag_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),.auto_in_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),.auto_in_w_ready(_axi4buf_auto_in_w_ready),.auto_in_w_valid(_axi4frag_auto_out_w_valid),.auto_in_w_bits_data(_axi4frag_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4frag_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4frag_auto_out_w_bits_last),.auto_in_b_ready(_axi4frag_auto_out_b_ready),.auto_in_b_valid(_axi4buf_auto_in_b_valid),.auto_in_b_bits_id(_axi4buf_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4buf_auto_in_b_bits_resp),.auto_in_b_bits_echo_real_last(_axi4buf_auto_in_b_bits_echo_real_last),.auto_in_ar_ready(_axi4buf_auto_in_ar_ready),.auto_in_ar_valid(_axi4frag_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4frag_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),.auto_in_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),.auto_in_r_ready(_axi4frag_auto_out_r_ready),.auto_in_r_valid(_axi4buf_auto_in_r_valid),.auto_in_r_bits_id(_axi4buf_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4buf_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4buf_auto_in_r_bits_resp),.auto_in_r_bits_echo_real_last(_axi4buf_auto_in_r_bits_echo_real_last),.auto_in_r_bits_last(_axi4buf_auto_in_r_bits_last),.auto_out_aw_ready(_srams_auto_in_aw_ready),.auto_out_aw_valid(_axi4buf_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4buf_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4buf_auto_out_aw_bits_addr),.auto_out_aw_bits_echo_real_last(_axi4buf_auto_out_aw_bits_echo_real_last),.auto_out_w_ready(_srams_auto_in_w_ready),.auto_out_w_valid(_axi4buf_auto_out_w_valid),.auto_out_w_bits_data(_axi4buf_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4buf_auto_out_w_bits_strb),.auto_out_b_ready(_axi4buf_auto_out_b_ready),.auto_out_b_valid(_srams_auto_in_b_valid),.auto_out_b_bits_id(_srams_auto_in_b_bits_id),.auto_out_b_bits_resp(_srams_auto_in_b_bits_resp),.auto_out_b_bits_echo_real_last(_srams_auto_in_b_bits_echo_real_last),.auto_out_ar_ready(_srams_auto_in_ar_ready),.auto_out_ar_valid(_axi4buf_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4buf_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4buf_auto_out_ar_bits_addr),.auto_out_ar_bits_echo_real_last(_axi4buf_auto_out_ar_bits_echo_real_last),.auto_out_r_ready(_axi4buf_auto_out_r_ready),.auto_out_r_valid(_srams_auto_in_r_valid),.auto_out_r_bits_id(_srams_auto_in_r_bits_id),.auto_out_r_bits_data(_srams_auto_in_r_bits_data),.auto_out_r_bits_resp(_srams_auto_in_r_bits_resp),.auto_out_r_bits_echo_real_last(_srams_auto_in_r_bits_echo_real_last)); 
  AXI4Fragmenter_1 axi4frag(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4frag_auto_in_aw_ready),.auto_in_aw_valid(_axi4xbar_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4xbar_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4xbar_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4xbar_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4xbar_auto_out_aw_bits_size),.auto_in_aw_bits_burst(_axi4xbar_auto_out_aw_bits_burst),.auto_in_w_ready(_axi4frag_auto_in_w_ready),.auto_in_w_valid(_axi4xbar_auto_out_w_valid),.auto_in_w_bits_data(_axi4xbar_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4xbar_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4xbar_auto_out_w_bits_last),.auto_in_b_ready(_axi4xbar_auto_out_b_ready),.auto_in_b_valid(_axi4frag_auto_in_b_valid),.auto_in_b_bits_id(_axi4frag_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4frag_auto_in_b_bits_resp),.auto_in_ar_ready(_axi4frag_auto_in_ar_ready),.auto_in_ar_valid(_axi4xbar_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4xbar_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4xbar_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4xbar_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4xbar_auto_out_ar_bits_size),.auto_in_ar_bits_burst(_axi4xbar_auto_out_ar_bits_burst),.auto_in_r_ready(_axi4xbar_auto_out_r_ready),.auto_in_r_valid(_axi4frag_auto_in_r_valid),.auto_in_r_bits_id(_axi4frag_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4frag_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4frag_auto_in_r_bits_resp),.auto_in_r_bits_last(_axi4frag_auto_in_r_bits_last),.auto_out_aw_ready(_axi4buf_auto_in_aw_ready),.auto_out_aw_valid(_axi4frag_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4frag_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),.auto_out_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),.auto_out_w_ready(_axi4buf_auto_in_w_ready),.auto_out_w_valid(_axi4frag_auto_out_w_valid),.auto_out_w_bits_data(_axi4frag_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4frag_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4frag_auto_out_w_bits_last),.auto_out_b_ready(_axi4frag_auto_out_b_ready),.auto_out_b_valid(_axi4buf_auto_in_b_valid),.auto_out_b_bits_id(_axi4buf_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4buf_auto_in_b_bits_resp),.auto_out_b_bits_echo_real_last(_axi4buf_auto_in_b_bits_echo_real_last),.auto_out_ar_ready(_axi4buf_auto_in_ar_ready),.auto_out_ar_valid(_axi4frag_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4frag_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),.auto_out_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),.auto_out_r_ready(_axi4frag_auto_out_r_ready),.auto_out_r_valid(_axi4buf_auto_in_r_valid),.auto_out_r_bits_id(_axi4buf_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4buf_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4buf_auto_in_r_bits_resp),.auto_out_r_bits_echo_real_last(_axi4buf_auto_in_r_bits_echo_real_last),.auto_out_r_bits_last(_axi4buf_auto_in_r_bits_last)); 
endmodule
 
module mem_512x64 (
  input [8:0] R0_addr,
  input R0_en,
  input R0_clk,
  output [63:0] R0_data,
  input [8:0] W0_addr,
  input W0_en,
  input W0_clk,
  input [63:0] W0_data,
  input [7:0] W0_mask) ; 
   reg [63:0] Memory[0:511] ;  
   reg _R0_en_d0 ;  
   reg [8:0] _R0_addr_d0 ;  
  always @( posedge R0_clk)
       begin 
         _R0_en_d0 <=R0_en;
         _R0_addr_d0 <=R0_addr;
       end
  
  always @( posedge W0_clk)
       begin 
         if (W0_en&W0_mask[0])
            Memory [W0_addr][32'h0+:8]<=W0_data[7:0];
         if (W0_en&W0_mask[1])
            Memory [W0_addr][32'h8+:8]<=W0_data[15:8];
         if (W0_en&W0_mask[2])
            Memory [W0_addr][32'h10+:8]<=W0_data[23:16];
         if (W0_en&W0_mask[3])
            Memory [W0_addr][32'h18+:8]<=W0_data[31:24];
         if (W0_en&W0_mask[4])
            Memory [W0_addr][32'h20+:8]<=W0_data[39:32];
         if (W0_en&W0_mask[5])
            Memory [W0_addr][32'h28+:8]<=W0_data[47:40];
         if (W0_en&W0_mask[6])
            Memory [W0_addr][32'h30+:8]<=W0_data[55:48];
         if (W0_en&W0_mask[7])
            Memory [W0_addr][32'h38+:8]<=W0_data[63:56];
       end
  
  assign R0_data=_R0_en_d0 ? Memory[_R0_addr_d0]:64'bx; 
endmodule
 
module AXI4RAM_1 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input auto_in_aw_bits_echo_real_last,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_b_bits_echo_real_last,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input auto_in_ar_bits_echo_real_last,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_echo_real_last) ; 
   wire nodeIn_ar_ready ;  
   wire nodeIn_aw_ready ;  
   wire [63:0] _mem_ext_R0_data ;  
   wire w_sel0=auto_in_aw_bits_addr[30:12]==19'h60000 ;  
   reg w_full ;  
   reg [3:0] w_id ;  
   reg w_echo_real_last ;  
   reg r_sel1 ;  
   reg w_sel1 ;  
   wire _GEN=nodeIn_aw_ready&auto_in_aw_valid ;  
  assign nodeIn_aw_ready=auto_in_w_valid&(auto_in_b_ready|~w_full); 
   reg r_full ;  
   reg [3:0] r_id ;  
   reg r_echo_real_last ;  
   wire ren=nodeIn_ar_ready&auto_in_ar_valid ;  
   reg rdata_REG ;  
   reg [7:0] rdata_r_0 ;  
   reg [7:0] rdata_r_1 ;  
   reg [7:0] rdata_r_2 ;  
   reg [7:0] rdata_r_3 ;  
   reg [7:0] rdata_r_4 ;  
   reg [7:0] rdata_r_5 ;  
   reg [7:0] rdata_r_6 ;  
   reg [7:0] rdata_r_7 ;  
  assign nodeIn_ar_ready=auto_in_r_ready|~r_full; 
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              w_full <=1'h0;
              r_full <=1'h0;
            end 
          else 
            begin 
              w_full <=_GEN|~(auto_in_b_ready&w_full)&w_full;
              r_full <=ren|~(auto_in_r_ready&r_full)&r_full;
            end 
         if (_GEN)
            begin 
              w_id <=auto_in_aw_bits_id;
              w_echo_real_last <=auto_in_aw_bits_echo_real_last;
            end 
         r_sel1 <=auto_in_ar_bits_addr[30:12]==19'h60000;
         w_sel1 <=w_sel0;
         if (ren)
            begin 
              r_id <=auto_in_ar_bits_id;
              r_echo_real_last <=auto_in_ar_bits_echo_real_last;
            end 
         rdata_REG <=ren;
         if (rdata_REG)
            begin 
              rdata_r_0 <=_mem_ext_R0_data[7:0];
              rdata_r_1 <=_mem_ext_R0_data[15:8];
              rdata_r_2 <=_mem_ext_R0_data[23:16];
              rdata_r_3 <=_mem_ext_R0_data[31:24];
              rdata_r_4 <=_mem_ext_R0_data[39:32];
              rdata_r_5 <=_mem_ext_R0_data[47:40];
              rdata_r_6 <=_mem_ext_R0_data[55:48];
              rdata_r_7 <=_mem_ext_R0_data[63:56];
            end 
       end
  
  mem_512x64 mem_ext(.R0_addr(auto_in_ar_bits_addr[11:3]),.R0_en(ren),.R0_clk(clock),.R0_data(_mem_ext_R0_data),.W0_addr(auto_in_aw_bits_addr[11:3]),.W0_en(_GEN&w_sel0),.W0_clk(clock),.W0_data(auto_in_w_bits_data),.W0_mask(auto_in_w_bits_strb)); 
  assign auto_in_aw_ready=nodeIn_aw_ready; 
  assign auto_in_w_ready=auto_in_aw_valid&(auto_in_b_ready|~w_full); 
  assign auto_in_b_valid=w_full; 
  assign auto_in_b_bits_id=w_id; 
  assign auto_in_b_bits_resp=w_sel1 ? 2'h0:2'h3; 
  assign auto_in_b_bits_echo_real_last=w_echo_real_last; 
  assign auto_in_ar_ready=nodeIn_ar_ready; 
  assign auto_in_r_valid=r_full; 
  assign auto_in_r_bits_id=r_id; 
  assign auto_in_r_bits_data={rdata_REG ? _mem_ext_R0_data[63:56]:rdata_r_7,rdata_REG ? _mem_ext_R0_data[55:48]:rdata_r_6,rdata_REG ? _mem_ext_R0_data[47:40]:rdata_r_5,rdata_REG ? _mem_ext_R0_data[39:32]:rdata_r_4,rdata_REG ? _mem_ext_R0_data[31:24]:rdata_r_3,rdata_REG ? _mem_ext_R0_data[23:16]:rdata_r_2,rdata_REG ? _mem_ext_R0_data[15:8]:rdata_r_1,rdata_REG ? _mem_ext_R0_data[7:0]:rdata_r_0}; 
  assign auto_in_r_bits_resp=r_sel1 ? 2'h0:2'h3; 
  assign auto_in_r_bits_echo_real_last=r_echo_real_last; 
endmodule
 
module AXI4Xbar_1 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [1:0] auto_in_aw_bits_burst,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [1:0] auto_in_ar_bits_burst,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output [7:0] auto_out_aw_bits_len,
  output [2:0] auto_out_aw_bits_size,
  output [1:0] auto_out_aw_bits_burst,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output [7:0] auto_out_ar_bits_len,
  output [2:0] auto_out_ar_bits_size,
  output [1:0] auto_out_ar_bits_burst,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_last) ; 
  assign auto_in_aw_ready=auto_out_aw_ready; 
  assign auto_in_w_ready=auto_out_w_ready; 
  assign auto_in_b_valid=auto_out_b_valid; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp; 
  assign auto_in_ar_ready=auto_out_ar_ready; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_last=auto_out_r_bits_last; 
  assign auto_out_aw_valid=auto_in_aw_valid; 
  assign auto_out_aw_bits_id=auto_in_aw_bits_id; 
  assign auto_out_aw_bits_addr=auto_in_aw_bits_addr; 
  assign auto_out_aw_bits_len=auto_in_aw_bits_len; 
  assign auto_out_aw_bits_size=auto_in_aw_bits_size; 
  assign auto_out_aw_bits_burst=auto_in_aw_bits_burst; 
  assign auto_out_w_valid=auto_in_w_valid; 
  assign auto_out_w_bits_data=auto_in_w_bits_data; 
  assign auto_out_w_bits_strb=auto_in_w_bits_strb; 
  assign auto_out_w_bits_last=auto_in_w_bits_last; 
  assign auto_out_b_ready=auto_in_b_ready; 
  assign auto_out_ar_valid=auto_in_ar_valid; 
  assign auto_out_ar_bits_id=auto_in_ar_bits_id; 
  assign auto_out_ar_bits_addr=auto_in_ar_bits_addr; 
  assign auto_out_ar_bits_len=auto_in_ar_bits_len; 
  assign auto_out_ar_bits_size=auto_in_ar_bits_size; 
  assign auto_out_ar_bits_burst=auto_in_ar_bits_burst; 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module Queue_96 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [30:0] io_enq_bits_addr,
  input io_enq_bits_echo_real_last,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output io_deq_bits_echo_real_last) ; 
   reg wrap ;  
   reg wrap_1 ;  
   reg maybe_full ;  
   wire ptr_match=wrap==wrap_1 ;  
   wire empty=ptr_match&~maybe_full ;  
   wire full=ptr_match&maybe_full ;  
   wire do_enq=~full&io_enq_valid ;  
   wire do_deq=io_deq_ready&~empty ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              wrap <=1'h0;
              wrap_1 <=1'h0;
              maybe_full <=1'h0;
            end 
          else 
            begin 
              if (do_enq)
                 wrap <=wrap-1'h1;
              if (do_deq)
                 wrap_1 <=wrap_1-1'h1;
              if (~(do_enq==do_deq))
                 maybe_full <=do_enq;
            end 
       end
  
  ram_2x4 ram_id_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_id),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_id)); 
  ram_addr_2x31 ram_addr_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_addr),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_addr)); 
  ram_2x1 ram_echo_real_last_ext(.R0_addr(wrap_1),.R0_en(1'h1),.R0_clk(clock),.R0_data(io_deq_bits_echo_real_last),.W0_addr(wrap),.W0_en(do_enq),.W0_clk(clock),.W0_data(io_enq_bits_echo_real_last)); 
  assign io_enq_ready=~full; 
  assign io_deq_valid=~empty; 
endmodule
 
module AXI4Buffer_2 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input auto_in_aw_bits_echo_real_last,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_b_bits_echo_real_last,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input auto_in_ar_bits_echo_real_last,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_echo_real_last,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output auto_out_aw_bits_echo_real_last,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_b_bits_echo_real_last,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output auto_out_ar_bits_echo_real_last,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_echo_real_last) ; 
  Queue_96 nodeOut_aw_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_aw_ready),.io_enq_valid(auto_in_aw_valid),.io_enq_bits_id(auto_in_aw_bits_id),.io_enq_bits_addr(auto_in_aw_bits_addr),.io_enq_bits_echo_real_last(auto_in_aw_bits_echo_real_last),.io_deq_ready(auto_out_aw_ready),.io_deq_valid(auto_out_aw_valid),.io_deq_bits_id(auto_out_aw_bits_id),.io_deq_bits_addr(auto_out_aw_bits_addr),.io_deq_bits_echo_real_last(auto_out_aw_bits_echo_real_last)); 
  Queue_1 nodeOut_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_w_ready),.io_enq_valid(auto_in_w_valid),.io_enq_bits_data(auto_in_w_bits_data),.io_enq_bits_strb(auto_in_w_bits_strb),.io_enq_bits_last(auto_in_w_bits_last),.io_deq_ready(auto_out_w_ready),.io_deq_valid(auto_out_w_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last()); 
  Queue_88 nodeIn_b_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_b_ready),.io_enq_valid(auto_out_b_valid),.io_enq_bits_id(auto_out_b_bits_id),.io_enq_bits_resp(auto_out_b_bits_resp),.io_enq_bits_echo_real_last(auto_out_b_bits_echo_real_last),.io_deq_ready(auto_in_b_ready),.io_deq_valid(auto_in_b_valid),.io_deq_bits_id(auto_in_b_bits_id),.io_deq_bits_resp(auto_in_b_bits_resp),.io_deq_bits_echo_real_last(auto_in_b_bits_echo_real_last)); 
  Queue_96 nodeOut_ar_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_ar_ready),.io_enq_valid(auto_in_ar_valid),.io_enq_bits_id(auto_in_ar_bits_id),.io_enq_bits_addr(auto_in_ar_bits_addr),.io_enq_bits_echo_real_last(auto_in_ar_bits_echo_real_last),.io_deq_ready(auto_out_ar_ready),.io_deq_valid(auto_out_ar_valid),.io_deq_bits_id(auto_out_ar_bits_id),.io_deq_bits_addr(auto_out_ar_bits_addr),.io_deq_bits_echo_real_last(auto_out_ar_bits_echo_real_last)); 
  Queue_90 nodeIn_r_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_out_r_ready),.io_enq_valid(auto_out_r_valid),.io_enq_bits_id(auto_out_r_bits_id),.io_enq_bits_data(auto_out_r_bits_data),.io_enq_bits_resp(auto_out_r_bits_resp),.io_enq_bits_echo_real_last(auto_out_r_bits_echo_real_last),.io_deq_ready(auto_in_r_ready),.io_deq_valid(auto_in_r_valid),.io_deq_bits_id(auto_in_r_bits_id),.io_deq_bits_data(auto_in_r_bits_data),.io_deq_bits_resp(auto_in_r_bits_resp),.io_deq_bits_echo_real_last(auto_in_r_bits_echo_real_last),.io_deq_bits_last(auto_in_r_bits_last)); 
endmodule
 
module Queue_101 (
  input clock,
  input reset,
  output io_enq_ready,
  input io_enq_valid,
  input [3:0] io_enq_bits_id,
  input [30:0] io_enq_bits_addr,
  input [7:0] io_enq_bits_len,
  input [2:0] io_enq_bits_size,
  input [1:0] io_enq_bits_burst,
  input io_deq_ready,
  output io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst) ; 
   reg [1:0] ram_burst ;  
   reg [2:0] ram_size ;  
   reg [7:0] ram_len ;  
   reg [30:0] ram_addr ;  
   reg [3:0] ram_id ;  
   reg full ;  
   wire io_deq_valid_0=io_enq_valid|full ;  
   wire do_enq=~(~full&io_deq_ready)&~full&io_enq_valid ;  
  always @( posedge clock)
       begin 
         if (do_enq)
            begin 
              ram_burst <=io_enq_bits_burst;
              ram_size <=io_enq_bits_size;
              ram_len <=io_enq_bits_len;
              ram_addr <=io_enq_bits_addr;
              ram_id <=io_enq_bits_id;
            end 
         if (reset)
            full <=1'h0;
          else 
            if (~(do_enq==(full&io_deq_ready&io_deq_valid_0)))
               full <=do_enq;
       end
  
  assign io_enq_ready=~full; 
  assign io_deq_valid=io_deq_valid_0; 
  assign io_deq_bits_id=full ? ram_id:io_enq_bits_id; 
  assign io_deq_bits_addr=full ? ram_addr:io_enq_bits_addr; 
  assign io_deq_bits_len=full ? ram_len:io_enq_bits_len; 
  assign io_deq_bits_size=full ? ram_size:io_enq_bits_size; 
  assign io_deq_bits_burst=full ? ram_burst:io_enq_bits_burst; 
endmodule
 
module AXI4Fragmenter_2 (
  input clock,
  input reset,
  output auto_in_aw_ready,
  input auto_in_aw_valid,
  input [3:0] auto_in_aw_bits_id,
  input [30:0] auto_in_aw_bits_addr,
  input [7:0] auto_in_aw_bits_len,
  input [2:0] auto_in_aw_bits_size,
  input [1:0] auto_in_aw_bits_burst,
  output auto_in_w_ready,
  input auto_in_w_valid,
  input [63:0] auto_in_w_bits_data,
  input [7:0] auto_in_w_bits_strb,
  input auto_in_w_bits_last,
  input auto_in_b_ready,
  output auto_in_b_valid,
  output [3:0] auto_in_b_bits_id,
  output [1:0] auto_in_b_bits_resp,
  output auto_in_ar_ready,
  input auto_in_ar_valid,
  input [3:0] auto_in_ar_bits_id,
  input [30:0] auto_in_ar_bits_addr,
  input [7:0] auto_in_ar_bits_len,
  input [2:0] auto_in_ar_bits_size,
  input [1:0] auto_in_ar_bits_burst,
  input auto_in_r_ready,
  output auto_in_r_valid,
  output [3:0] auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0] auto_in_r_bits_resp,
  output auto_in_r_bits_last,
  input auto_out_aw_ready,
  output auto_out_aw_valid,
  output [3:0] auto_out_aw_bits_id,
  output [30:0] auto_out_aw_bits_addr,
  output auto_out_aw_bits_echo_real_last,
  input auto_out_w_ready,
  output auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0] auto_out_w_bits_strb,
  output auto_out_w_bits_last,
  output auto_out_b_ready,
  input auto_out_b_valid,
  input [3:0] auto_out_b_bits_id,
  input [1:0] auto_out_b_bits_resp,
  input auto_out_b_bits_echo_real_last,
  input auto_out_ar_ready,
  output auto_out_ar_valid,
  output [3:0] auto_out_ar_bits_id,
  output [30:0] auto_out_ar_bits_addr,
  output auto_out_ar_bits_echo_real_last,
  output auto_out_r_ready,
  input auto_out_r_valid,
  input [3:0] auto_out_r_bits_id,
  input [63:0] auto_out_r_bits_data,
  input [1:0] auto_out_r_bits_resp,
  input auto_out_r_bits_echo_real_last,
  input auto_out_r_bits_last) ; 
   wire nodeOut_w_valid ;  
   wire w_idle ;  
   wire in_aw_ready ;  
   wire _in_w_deq_q_io_deq_valid ;  
   wire _in_w_deq_q_io_deq_bits_last ;  
   wire _deq_q_1_io_deq_valid ;  
   wire [30:0] _deq_q_1_io_deq_bits_addr ;  
   wire [7:0] _deq_q_1_io_deq_bits_len ;  
   wire [2:0] _deq_q_1_io_deq_bits_size ;  
   wire [1:0] _deq_q_1_io_deq_bits_burst ;  
   wire _deq_q_io_deq_valid ;  
   wire [30:0] _deq_q_io_deq_bits_addr ;  
   wire [7:0] _deq_q_io_deq_bits_len ;  
   wire [2:0] _deq_q_io_deq_bits_size ;  
   wire [1:0] _deq_q_io_deq_bits_burst ;  
   reg busy ;  
   reg [30:0] r_addr ;  
   reg [7:0] r_len ;  
   wire [7:0] len=busy ? r_len:_deq_q_io_deq_bits_len ;  
   wire [30:0] addr=busy ? r_addr:_deq_q_io_deq_bits_addr ;  
   wire [30:0] _out_bits_addr_T=~addr ;  
   wire [9:0] _out_bits_addr_T_2=10'h7<<_deq_q_io_deq_bits_size ;  
   reg busy_1 ;  
   reg [30:0] r_addr_1 ;  
   reg [7:0] r_len_1 ;  
   wire [7:0] len_1=busy_1 ? r_len_1:_deq_q_1_io_deq_bits_len ;  
   wire [30:0] addr_1=busy_1 ? r_addr_1:_deq_q_1_io_deq_bits_addr ;  
   wire [30:0] _out_bits_addr_T_7=~addr_1 ;  
   wire [9:0] _out_bits_addr_T_9=10'h7<<_deq_q_1_io_deq_bits_size ;  
   reg wbeats_latched ;  
   wire _in_aw_ready_T=w_idle|wbeats_latched ;  
   wire nodeOut_aw_valid=_deq_q_1_io_deq_valid&_in_aw_ready_T ;  
  assign in_aw_ready=auto_out_aw_ready&_in_aw_ready_T; 
   wire wbeats_valid=_deq_q_1_io_deq_valid&~wbeats_latched ;  
   reg [8:0] w_counter ;  
  assign w_idle=w_counter==9'h0; 
   wire [8:0] w_todo=w_idle ? {8'h0,wbeats_valid}:w_counter ;  
   wire w_last=w_todo==9'h1 ;  
   wire _w_counter_T=auto_out_w_ready&nodeOut_w_valid ;  
  assign nodeOut_w_valid=_in_w_deq_q_io_deq_valid&(~w_idle|wbeats_valid); 
  always @( posedge clock)
       begin 
         if (~reset&~(~_w_counter_T|(|w_todo)))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:177 assert (!out.w.fire || w_todo =/= 0.U) // underflow impossible\n");
              if (1)$display("");
            end 
         if (~reset&~(~nodeOut_w_valid|~_in_w_deq_q_io_deq_bits_last|w_last))
            begin 
              if (1)$display("Assertion failed\n    at Fragmenter.scala:186 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
              if (1)$display("");
            end 
       end
  
   wire nodeOut_b_ready=auto_in_b_ready|~auto_out_b_bits_echo_real_last ;  
   reg [1:0] error_0 ;  
   reg [1:0] error_1 ;  
   reg [1:0] error_2 ;  
   reg [1:0] error_3 ;  
   reg [1:0] error_4 ;  
   reg [1:0] error_5 ;  
   reg [1:0] error_6 ;  
   reg [1:0] error_7 ;  
   reg [1:0] error_8 ;  
   reg [1:0] error_9 ;  
   reg [1:0] error_10 ;  
   reg [1:0] error_11 ;  
   reg [1:0] error_12 ;  
   reg [1:0] error_13 ;  
   reg [1:0] error_14 ;  
   reg [1:0] error_15 ;  
   reg [1:0] casez_tmp ;  
  always @(*)
       begin 
         casez (auto_out_b_bits_id)
          4 'b0000:
             casez_tmp =error_0;
          4 'b0001:
             casez_tmp =error_1;
          4 'b0010:
             casez_tmp =error_2;
          4 'b0011:
             casez_tmp =error_3;
          4 'b0100:
             casez_tmp =error_4;
          4 'b0101:
             casez_tmp =error_5;
          4 'b0110:
             casez_tmp =error_6;
          4 'b0111:
             casez_tmp =error_7;
          4 'b1000:
             casez_tmp =error_8;
          4 'b1001:
             casez_tmp =error_9;
          4 'b1010:
             casez_tmp =error_10;
          4 'b1011:
             casez_tmp =error_11;
          4 'b1100:
             casez_tmp =error_12;
          4 'b1101:
             casez_tmp =error_13;
          4 'b1110:
             casez_tmp =error_14;
          default :
             casez_tmp =error_15;
         endcase 
       end
  
   wire _GEN=nodeOut_b_ready&auto_out_b_valid ;  
   wire [22:0] _wrapMask_T_1={7'h0,_deq_q_io_deq_bits_len,8'hFF}<<_deq_q_io_deq_bits_size ;  
   wire [30:0] _mux_addr_T_1=~_deq_q_io_deq_bits_addr ;  
   wire [30:0] _inc_addr_T_1=addr+{15'h0,16'h1<<_deq_q_io_deq_bits_size} ;  
   wire [22:0] _wrapMask_T_3={7'h0,_deq_q_1_io_deq_bits_len,8'hFF}<<_deq_q_1_io_deq_bits_size ;  
   wire [30:0] _mux_addr_T_6=~_deq_q_1_io_deq_bits_addr ;  
   wire [30:0] _inc_addr_T_3=addr_1+{15'h0,16'h1<<_deq_q_1_io_deq_bits_size} ;  
   wire _GEN_0=auto_out_ar_ready&_deq_q_io_deq_valid ;  
   wire _GEN_1=in_aw_ready&_deq_q_1_io_deq_valid ;  
  always @( posedge clock)
       begin 
         if (reset)
            begin 
              busy <=1'h0;
              busy_1 <=1'h0;
              wbeats_latched <=1'h0;
              w_counter <=9'h0;
              error_0 <=2'h0;
              error_1 <=2'h0;
              error_2 <=2'h0;
              error_3 <=2'h0;
              error_4 <=2'h0;
              error_5 <=2'h0;
              error_6 <=2'h0;
              error_7 <=2'h0;
              error_8 <=2'h0;
              error_9 <=2'h0;
              error_10 <=2'h0;
              error_11 <=2'h0;
              error_12 <=2'h0;
              error_13 <=2'h0;
              error_14 <=2'h0;
              error_15 <=2'h0;
            end 
          else 
            begin 
              if (_GEN_0)
                 busy <=|len;
              if (_GEN_1)
                 busy_1 <=|len_1;
              wbeats_latched <=~(auto_out_aw_ready&nodeOut_aw_valid)&(wbeats_valid&w_idle|wbeats_latched);
              w_counter <=w_todo-{8'h0,_w_counter_T};
              if (auto_out_b_bits_id==4'h0&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_0 <=2'h0;
                    else 
                      error_0 <=error_0|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h1&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_1 <=2'h0;
                    else 
                      error_1 <=error_1|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h2&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_2 <=2'h0;
                    else 
                      error_2 <=error_2|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h3&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_3 <=2'h0;
                    else 
                      error_3 <=error_3|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h4&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_4 <=2'h0;
                    else 
                      error_4 <=error_4|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h5&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_5 <=2'h0;
                    else 
                      error_5 <=error_5|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h6&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_6 <=2'h0;
                    else 
                      error_6 <=error_6|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h7&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_7 <=2'h0;
                    else 
                      error_7 <=error_7|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h8&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_8 <=2'h0;
                    else 
                      error_8 <=error_8|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'h9&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_9 <=2'h0;
                    else 
                      error_9 <=error_9|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hA&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_10 <=2'h0;
                    else 
                      error_10 <=error_10|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hB&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_11 <=2'h0;
                    else 
                      error_11 <=error_11|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hC&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_12 <=2'h0;
                    else 
                      error_12 <=error_12|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hD&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_13 <=2'h0;
                    else 
                      error_13 <=error_13|auto_out_b_bits_resp;
                 end 
              if (auto_out_b_bits_id==4'hE&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_14 <=2'h0;
                    else 
                      error_14 <=error_14|auto_out_b_bits_resp;
                 end 
              if ((&auto_out_b_bits_id)&_GEN)
                 begin 
                   if (auto_out_b_bits_echo_real_last)
                      error_15 <=2'h0;
                    else 
                      error_15 <=error_15|auto_out_b_bits_resp;
                 end 
            end 
         if (_GEN_0)
            begin 
              if (_deq_q_io_deq_bits_burst==2'h0)
                 r_addr <=_deq_q_io_deq_bits_addr;
               else 
                 if (_deq_q_io_deq_bits_burst==2'h2)
                    r_addr <={16'h0,_inc_addr_T_1[14:0]&_wrapMask_T_1[22:8]}|~{_mux_addr_T_1[30:15],_mux_addr_T_1[14:0]|_wrapMask_T_1[22:8]};
                  else 
                    r_addr <=_inc_addr_T_1;
              r_len <=len-8'h1;
            end 
         if (_GEN_1)
            begin 
              if (_deq_q_1_io_deq_bits_burst==2'h0)
                 r_addr_1 <=_deq_q_1_io_deq_bits_addr;
               else 
                 if (_deq_q_1_io_deq_bits_burst==2'h2)
                    r_addr_1 <={16'h0,_inc_addr_T_3[14:0]&_wrapMask_T_3[22:8]}|~{_mux_addr_T_6[30:15],_mux_addr_T_6[14:0]|_wrapMask_T_3[22:8]};
                  else 
                    r_addr_1 <=_inc_addr_T_3;
              r_len_1 <=len_1-8'h1;
            end 
       end
  
  Queue_101 deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_ar_ready),.io_enq_valid(auto_in_ar_valid),.io_enq_bits_id(auto_in_ar_bits_id),.io_enq_bits_addr(auto_in_ar_bits_addr),.io_enq_bits_len(auto_in_ar_bits_len),.io_enq_bits_size(auto_in_ar_bits_size),.io_enq_bits_burst(auto_in_ar_bits_burst),.io_deq_ready(auto_out_ar_ready&~(|len)),.io_deq_valid(_deq_q_io_deq_valid),.io_deq_bits_id(auto_out_ar_bits_id),.io_deq_bits_addr(_deq_q_io_deq_bits_addr),.io_deq_bits_len(_deq_q_io_deq_bits_len),.io_deq_bits_size(_deq_q_io_deq_bits_size),.io_deq_bits_burst(_deq_q_io_deq_bits_burst)); 
  Queue_101 deq_q_1(.clock(clock),.reset(reset),.io_enq_ready(auto_in_aw_ready),.io_enq_valid(auto_in_aw_valid),.io_enq_bits_id(auto_in_aw_bits_id),.io_enq_bits_addr(auto_in_aw_bits_addr),.io_enq_bits_len(auto_in_aw_bits_len),.io_enq_bits_size(auto_in_aw_bits_size),.io_enq_bits_burst(auto_in_aw_bits_burst),.io_deq_ready(in_aw_ready&~(|len_1)),.io_deq_valid(_deq_q_1_io_deq_valid),.io_deq_bits_id(auto_out_aw_bits_id),.io_deq_bits_addr(_deq_q_1_io_deq_bits_addr),.io_deq_bits_len(_deq_q_1_io_deq_bits_len),.io_deq_bits_size(_deq_q_1_io_deq_bits_size),.io_deq_bits_burst(_deq_q_1_io_deq_bits_burst)); 
  Queue_34 in_w_deq_q(.clock(clock),.reset(reset),.io_enq_ready(auto_in_w_ready),.io_enq_valid(auto_in_w_valid),.io_enq_bits_data(auto_in_w_bits_data),.io_enq_bits_strb(auto_in_w_bits_strb),.io_enq_bits_last(auto_in_w_bits_last),.io_deq_ready(auto_out_w_ready&(~w_idle|wbeats_valid)),.io_deq_valid(_in_w_deq_q_io_deq_valid),.io_deq_bits_data(auto_out_w_bits_data),.io_deq_bits_strb(auto_out_w_bits_strb),.io_deq_bits_last(_in_w_deq_q_io_deq_bits_last)); 
  assign auto_in_b_valid=auto_out_b_valid&auto_out_b_bits_echo_real_last; 
  assign auto_in_b_bits_id=auto_out_b_bits_id; 
  assign auto_in_b_bits_resp=auto_out_b_bits_resp|casez_tmp; 
  assign auto_in_r_valid=auto_out_r_valid; 
  assign auto_in_r_bits_id=auto_out_r_bits_id; 
  assign auto_in_r_bits_data=auto_out_r_bits_data; 
  assign auto_in_r_bits_resp=auto_out_r_bits_resp; 
  assign auto_in_r_bits_last=auto_out_r_bits_last&auto_out_r_bits_echo_real_last; 
  assign auto_out_aw_valid=nodeOut_aw_valid; 
  assign auto_out_aw_bits_addr=~{_out_bits_addr_T_7[30:3],_out_bits_addr_T_7[2:0]|~(_out_bits_addr_T_9[2:0])}; 
  assign auto_out_aw_bits_echo_real_last=~(|len_1); 
  assign auto_out_w_valid=nodeOut_w_valid; 
  assign auto_out_w_bits_last=w_last; 
  assign auto_out_b_ready=nodeOut_b_ready; 
  assign auto_out_ar_valid=_deq_q_io_deq_valid; 
  assign auto_out_ar_bits_addr=~{_out_bits_addr_T[30:3],_out_bits_addr_T[2:0]|~(_out_bits_addr_T_2[2:0])}; 
  assign auto_out_ar_bits_echo_real_last=~(|len); 
  assign auto_out_r_ready=auto_in_r_ready; 
endmodule
 
module SimAXIMem_1 (
  input clock,
  input reset,
  output io_axi4_0_aw_ready,
  input io_axi4_0_aw_valid,
  input [3:0] io_axi4_0_aw_bits_id,
  input [30:0] io_axi4_0_aw_bits_addr,
  input [7:0] io_axi4_0_aw_bits_len,
  input [2:0] io_axi4_0_aw_bits_size,
  input [1:0] io_axi4_0_aw_bits_burst,
  output io_axi4_0_w_ready,
  input io_axi4_0_w_valid,
  input [63:0] io_axi4_0_w_bits_data,
  input [7:0] io_axi4_0_w_bits_strb,
  input io_axi4_0_w_bits_last,
  input io_axi4_0_b_ready,
  output io_axi4_0_b_valid,
  output [3:0] io_axi4_0_b_bits_id,
  output [1:0] io_axi4_0_b_bits_resp,
  output io_axi4_0_ar_ready,
  input io_axi4_0_ar_valid,
  input [3:0] io_axi4_0_ar_bits_id,
  input [30:0] io_axi4_0_ar_bits_addr,
  input [7:0] io_axi4_0_ar_bits_len,
  input [2:0] io_axi4_0_ar_bits_size,
  input [1:0] io_axi4_0_ar_bits_burst,
  input io_axi4_0_r_ready,
  output io_axi4_0_r_valid,
  output [3:0] io_axi4_0_r_bits_id,
  output [63:0] io_axi4_0_r_bits_data,
  output [1:0] io_axi4_0_r_bits_resp,
  output io_axi4_0_r_bits_last) ; 
   wire _axi4frag_auto_in_aw_ready ;  
   wire _axi4frag_auto_in_w_ready ;  
   wire _axi4frag_auto_in_b_valid ;  
   wire [3:0] _axi4frag_auto_in_b_bits_id ;  
   wire [1:0] _axi4frag_auto_in_b_bits_resp ;  
   wire _axi4frag_auto_in_ar_ready ;  
   wire _axi4frag_auto_in_r_valid ;  
   wire [3:0] _axi4frag_auto_in_r_bits_id ;  
   wire [63:0] _axi4frag_auto_in_r_bits_data ;  
   wire [1:0] _axi4frag_auto_in_r_bits_resp ;  
   wire _axi4frag_auto_in_r_bits_last ;  
   wire _axi4frag_auto_out_aw_valid ;  
   wire [3:0] _axi4frag_auto_out_aw_bits_id ;  
   wire [30:0] _axi4frag_auto_out_aw_bits_addr ;  
   wire _axi4frag_auto_out_aw_bits_echo_real_last ;  
   wire _axi4frag_auto_out_w_valid ;  
   wire [63:0] _axi4frag_auto_out_w_bits_data ;  
   wire [7:0] _axi4frag_auto_out_w_bits_strb ;  
   wire _axi4frag_auto_out_w_bits_last ;  
   wire _axi4frag_auto_out_b_ready ;  
   wire _axi4frag_auto_out_ar_valid ;  
   wire [3:0] _axi4frag_auto_out_ar_bits_id ;  
   wire [30:0] _axi4frag_auto_out_ar_bits_addr ;  
   wire _axi4frag_auto_out_ar_bits_echo_real_last ;  
   wire _axi4frag_auto_out_r_ready ;  
   wire _axi4buf_auto_in_aw_ready ;  
   wire _axi4buf_auto_in_w_ready ;  
   wire _axi4buf_auto_in_b_valid ;  
   wire [3:0] _axi4buf_auto_in_b_bits_id ;  
   wire [1:0] _axi4buf_auto_in_b_bits_resp ;  
   wire _axi4buf_auto_in_b_bits_echo_real_last ;  
   wire _axi4buf_auto_in_ar_ready ;  
   wire _axi4buf_auto_in_r_valid ;  
   wire [3:0] _axi4buf_auto_in_r_bits_id ;  
   wire [63:0] _axi4buf_auto_in_r_bits_data ;  
   wire [1:0] _axi4buf_auto_in_r_bits_resp ;  
   wire _axi4buf_auto_in_r_bits_echo_real_last ;  
   wire _axi4buf_auto_in_r_bits_last ;  
   wire _axi4buf_auto_out_aw_valid ;  
   wire [3:0] _axi4buf_auto_out_aw_bits_id ;  
   wire [30:0] _axi4buf_auto_out_aw_bits_addr ;  
   wire _axi4buf_auto_out_aw_bits_echo_real_last ;  
   wire _axi4buf_auto_out_w_valid ;  
   wire [63:0] _axi4buf_auto_out_w_bits_data ;  
   wire [7:0] _axi4buf_auto_out_w_bits_strb ;  
   wire _axi4buf_auto_out_b_ready ;  
   wire _axi4buf_auto_out_ar_valid ;  
   wire [3:0] _axi4buf_auto_out_ar_bits_id ;  
   wire [30:0] _axi4buf_auto_out_ar_bits_addr ;  
   wire _axi4buf_auto_out_ar_bits_echo_real_last ;  
   wire _axi4buf_auto_out_r_ready ;  
   wire _axi4xbar_auto_out_aw_valid ;  
   wire [3:0] _axi4xbar_auto_out_aw_bits_id ;  
   wire [30:0] _axi4xbar_auto_out_aw_bits_addr ;  
   wire [7:0] _axi4xbar_auto_out_aw_bits_len ;  
   wire [2:0] _axi4xbar_auto_out_aw_bits_size ;  
   wire [1:0] _axi4xbar_auto_out_aw_bits_burst ;  
   wire _axi4xbar_auto_out_w_valid ;  
   wire [63:0] _axi4xbar_auto_out_w_bits_data ;  
   wire [7:0] _axi4xbar_auto_out_w_bits_strb ;  
   wire _axi4xbar_auto_out_w_bits_last ;  
   wire _axi4xbar_auto_out_b_ready ;  
   wire _axi4xbar_auto_out_ar_valid ;  
   wire [3:0] _axi4xbar_auto_out_ar_bits_id ;  
   wire [30:0] _axi4xbar_auto_out_ar_bits_addr ;  
   wire [7:0] _axi4xbar_auto_out_ar_bits_len ;  
   wire [2:0] _axi4xbar_auto_out_ar_bits_size ;  
   wire [1:0] _axi4xbar_auto_out_ar_bits_burst ;  
   wire _axi4xbar_auto_out_r_ready ;  
   wire _srams_auto_in_aw_ready ;  
   wire _srams_auto_in_w_ready ;  
   wire _srams_auto_in_b_valid ;  
   wire [3:0] _srams_auto_in_b_bits_id ;  
   wire [1:0] _srams_auto_in_b_bits_resp ;  
   wire _srams_auto_in_b_bits_echo_real_last ;  
   wire _srams_auto_in_ar_ready ;  
   wire _srams_auto_in_r_valid ;  
   wire [3:0] _srams_auto_in_r_bits_id ;  
   wire [63:0] _srams_auto_in_r_bits_data ;  
   wire [1:0] _srams_auto_in_r_bits_resp ;  
   wire _srams_auto_in_r_bits_echo_real_last ;  
  AXI4RAM_1 srams(.clock(clock),.reset(reset),.auto_in_aw_ready(_srams_auto_in_aw_ready),.auto_in_aw_valid(_axi4buf_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4buf_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4buf_auto_out_aw_bits_addr),.auto_in_aw_bits_echo_real_last(_axi4buf_auto_out_aw_bits_echo_real_last),.auto_in_w_ready(_srams_auto_in_w_ready),.auto_in_w_valid(_axi4buf_auto_out_w_valid),.auto_in_w_bits_data(_axi4buf_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4buf_auto_out_w_bits_strb),.auto_in_b_ready(_axi4buf_auto_out_b_ready),.auto_in_b_valid(_srams_auto_in_b_valid),.auto_in_b_bits_id(_srams_auto_in_b_bits_id),.auto_in_b_bits_resp(_srams_auto_in_b_bits_resp),.auto_in_b_bits_echo_real_last(_srams_auto_in_b_bits_echo_real_last),.auto_in_ar_ready(_srams_auto_in_ar_ready),.auto_in_ar_valid(_axi4buf_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4buf_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4buf_auto_out_ar_bits_addr),.auto_in_ar_bits_echo_real_last(_axi4buf_auto_out_ar_bits_echo_real_last),.auto_in_r_ready(_axi4buf_auto_out_r_ready),.auto_in_r_valid(_srams_auto_in_r_valid),.auto_in_r_bits_id(_srams_auto_in_r_bits_id),.auto_in_r_bits_data(_srams_auto_in_r_bits_data),.auto_in_r_bits_resp(_srams_auto_in_r_bits_resp),.auto_in_r_bits_echo_real_last(_srams_auto_in_r_bits_echo_real_last)); 
  AXI4Xbar_1 axi4xbar(.clock(clock),.reset(reset),.auto_in_aw_ready(io_axi4_0_aw_ready),.auto_in_aw_valid(io_axi4_0_aw_valid),.auto_in_aw_bits_id(io_axi4_0_aw_bits_id),.auto_in_aw_bits_addr(io_axi4_0_aw_bits_addr),.auto_in_aw_bits_len(io_axi4_0_aw_bits_len),.auto_in_aw_bits_size(io_axi4_0_aw_bits_size),.auto_in_aw_bits_burst(io_axi4_0_aw_bits_burst),.auto_in_w_ready(io_axi4_0_w_ready),.auto_in_w_valid(io_axi4_0_w_valid),.auto_in_w_bits_data(io_axi4_0_w_bits_data),.auto_in_w_bits_strb(io_axi4_0_w_bits_strb),.auto_in_w_bits_last(io_axi4_0_w_bits_last),.auto_in_b_ready(io_axi4_0_b_ready),.auto_in_b_valid(io_axi4_0_b_valid),.auto_in_b_bits_id(io_axi4_0_b_bits_id),.auto_in_b_bits_resp(io_axi4_0_b_bits_resp),.auto_in_ar_ready(io_axi4_0_ar_ready),.auto_in_ar_valid(io_axi4_0_ar_valid),.auto_in_ar_bits_id(io_axi4_0_ar_bits_id),.auto_in_ar_bits_addr(io_axi4_0_ar_bits_addr),.auto_in_ar_bits_len(io_axi4_0_ar_bits_len),.auto_in_ar_bits_size(io_axi4_0_ar_bits_size),.auto_in_ar_bits_burst(io_axi4_0_ar_bits_burst),.auto_in_r_ready(io_axi4_0_r_ready),.auto_in_r_valid(io_axi4_0_r_valid),.auto_in_r_bits_id(io_axi4_0_r_bits_id),.auto_in_r_bits_data(io_axi4_0_r_bits_data),.auto_in_r_bits_resp(io_axi4_0_r_bits_resp),.auto_in_r_bits_last(io_axi4_0_r_bits_last),.auto_out_aw_ready(_axi4frag_auto_in_aw_ready),.auto_out_aw_valid(_axi4xbar_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4xbar_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4xbar_auto_out_aw_bits_addr),.auto_out_aw_bits_len(_axi4xbar_auto_out_aw_bits_len),.auto_out_aw_bits_size(_axi4xbar_auto_out_aw_bits_size),.auto_out_aw_bits_burst(_axi4xbar_auto_out_aw_bits_burst),.auto_out_w_ready(_axi4frag_auto_in_w_ready),.auto_out_w_valid(_axi4xbar_auto_out_w_valid),.auto_out_w_bits_data(_axi4xbar_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4xbar_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4xbar_auto_out_w_bits_last),.auto_out_b_ready(_axi4xbar_auto_out_b_ready),.auto_out_b_valid(_axi4frag_auto_in_b_valid),.auto_out_b_bits_id(_axi4frag_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4frag_auto_in_b_bits_resp),.auto_out_ar_ready(_axi4frag_auto_in_ar_ready),.auto_out_ar_valid(_axi4xbar_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4xbar_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4xbar_auto_out_ar_bits_addr),.auto_out_ar_bits_len(_axi4xbar_auto_out_ar_bits_len),.auto_out_ar_bits_size(_axi4xbar_auto_out_ar_bits_size),.auto_out_ar_bits_burst(_axi4xbar_auto_out_ar_bits_burst),.auto_out_r_ready(_axi4xbar_auto_out_r_ready),.auto_out_r_valid(_axi4frag_auto_in_r_valid),.auto_out_r_bits_id(_axi4frag_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4frag_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4frag_auto_in_r_bits_resp),.auto_out_r_bits_last(_axi4frag_auto_in_r_bits_last)); 
  AXI4Buffer_2 axi4buf(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4buf_auto_in_aw_ready),.auto_in_aw_valid(_axi4frag_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4frag_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),.auto_in_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),.auto_in_w_ready(_axi4buf_auto_in_w_ready),.auto_in_w_valid(_axi4frag_auto_out_w_valid),.auto_in_w_bits_data(_axi4frag_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4frag_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4frag_auto_out_w_bits_last),.auto_in_b_ready(_axi4frag_auto_out_b_ready),.auto_in_b_valid(_axi4buf_auto_in_b_valid),.auto_in_b_bits_id(_axi4buf_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4buf_auto_in_b_bits_resp),.auto_in_b_bits_echo_real_last(_axi4buf_auto_in_b_bits_echo_real_last),.auto_in_ar_ready(_axi4buf_auto_in_ar_ready),.auto_in_ar_valid(_axi4frag_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4frag_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),.auto_in_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),.auto_in_r_ready(_axi4frag_auto_out_r_ready),.auto_in_r_valid(_axi4buf_auto_in_r_valid),.auto_in_r_bits_id(_axi4buf_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4buf_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4buf_auto_in_r_bits_resp),.auto_in_r_bits_echo_real_last(_axi4buf_auto_in_r_bits_echo_real_last),.auto_in_r_bits_last(_axi4buf_auto_in_r_bits_last),.auto_out_aw_ready(_srams_auto_in_aw_ready),.auto_out_aw_valid(_axi4buf_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4buf_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4buf_auto_out_aw_bits_addr),.auto_out_aw_bits_echo_real_last(_axi4buf_auto_out_aw_bits_echo_real_last),.auto_out_w_ready(_srams_auto_in_w_ready),.auto_out_w_valid(_axi4buf_auto_out_w_valid),.auto_out_w_bits_data(_axi4buf_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4buf_auto_out_w_bits_strb),.auto_out_b_ready(_axi4buf_auto_out_b_ready),.auto_out_b_valid(_srams_auto_in_b_valid),.auto_out_b_bits_id(_srams_auto_in_b_bits_id),.auto_out_b_bits_resp(_srams_auto_in_b_bits_resp),.auto_out_b_bits_echo_real_last(_srams_auto_in_b_bits_echo_real_last),.auto_out_ar_ready(_srams_auto_in_ar_ready),.auto_out_ar_valid(_axi4buf_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4buf_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4buf_auto_out_ar_bits_addr),.auto_out_ar_bits_echo_real_last(_axi4buf_auto_out_ar_bits_echo_real_last),.auto_out_r_ready(_axi4buf_auto_out_r_ready),.auto_out_r_valid(_srams_auto_in_r_valid),.auto_out_r_bits_id(_srams_auto_in_r_bits_id),.auto_out_r_bits_data(_srams_auto_in_r_bits_data),.auto_out_r_bits_resp(_srams_auto_in_r_bits_resp),.auto_out_r_bits_echo_real_last(_srams_auto_in_r_bits_echo_real_last)); 
  AXI4Fragmenter_2 axi4frag(.clock(clock),.reset(reset),.auto_in_aw_ready(_axi4frag_auto_in_aw_ready),.auto_in_aw_valid(_axi4xbar_auto_out_aw_valid),.auto_in_aw_bits_id(_axi4xbar_auto_out_aw_bits_id),.auto_in_aw_bits_addr(_axi4xbar_auto_out_aw_bits_addr),.auto_in_aw_bits_len(_axi4xbar_auto_out_aw_bits_len),.auto_in_aw_bits_size(_axi4xbar_auto_out_aw_bits_size),.auto_in_aw_bits_burst(_axi4xbar_auto_out_aw_bits_burst),.auto_in_w_ready(_axi4frag_auto_in_w_ready),.auto_in_w_valid(_axi4xbar_auto_out_w_valid),.auto_in_w_bits_data(_axi4xbar_auto_out_w_bits_data),.auto_in_w_bits_strb(_axi4xbar_auto_out_w_bits_strb),.auto_in_w_bits_last(_axi4xbar_auto_out_w_bits_last),.auto_in_b_ready(_axi4xbar_auto_out_b_ready),.auto_in_b_valid(_axi4frag_auto_in_b_valid),.auto_in_b_bits_id(_axi4frag_auto_in_b_bits_id),.auto_in_b_bits_resp(_axi4frag_auto_in_b_bits_resp),.auto_in_ar_ready(_axi4frag_auto_in_ar_ready),.auto_in_ar_valid(_axi4xbar_auto_out_ar_valid),.auto_in_ar_bits_id(_axi4xbar_auto_out_ar_bits_id),.auto_in_ar_bits_addr(_axi4xbar_auto_out_ar_bits_addr),.auto_in_ar_bits_len(_axi4xbar_auto_out_ar_bits_len),.auto_in_ar_bits_size(_axi4xbar_auto_out_ar_bits_size),.auto_in_ar_bits_burst(_axi4xbar_auto_out_ar_bits_burst),.auto_in_r_ready(_axi4xbar_auto_out_r_ready),.auto_in_r_valid(_axi4frag_auto_in_r_valid),.auto_in_r_bits_id(_axi4frag_auto_in_r_bits_id),.auto_in_r_bits_data(_axi4frag_auto_in_r_bits_data),.auto_in_r_bits_resp(_axi4frag_auto_in_r_bits_resp),.auto_in_r_bits_last(_axi4frag_auto_in_r_bits_last),.auto_out_aw_ready(_axi4buf_auto_in_aw_ready),.auto_out_aw_valid(_axi4frag_auto_out_aw_valid),.auto_out_aw_bits_id(_axi4frag_auto_out_aw_bits_id),.auto_out_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),.auto_out_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),.auto_out_w_ready(_axi4buf_auto_in_w_ready),.auto_out_w_valid(_axi4frag_auto_out_w_valid),.auto_out_w_bits_data(_axi4frag_auto_out_w_bits_data),.auto_out_w_bits_strb(_axi4frag_auto_out_w_bits_strb),.auto_out_w_bits_last(_axi4frag_auto_out_w_bits_last),.auto_out_b_ready(_axi4frag_auto_out_b_ready),.auto_out_b_valid(_axi4buf_auto_in_b_valid),.auto_out_b_bits_id(_axi4buf_auto_in_b_bits_id),.auto_out_b_bits_resp(_axi4buf_auto_in_b_bits_resp),.auto_out_b_bits_echo_real_last(_axi4buf_auto_in_b_bits_echo_real_last),.auto_out_ar_ready(_axi4buf_auto_in_ar_ready),.auto_out_ar_valid(_axi4frag_auto_out_ar_valid),.auto_out_ar_bits_id(_axi4frag_auto_out_ar_bits_id),.auto_out_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),.auto_out_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),.auto_out_r_ready(_axi4frag_auto_out_r_ready),.auto_out_r_valid(_axi4buf_auto_in_r_valid),.auto_out_r_bits_id(_axi4buf_auto_in_r_bits_id),.auto_out_r_bits_data(_axi4buf_auto_in_r_bits_data),.auto_out_r_bits_resp(_axi4buf_auto_in_r_bits_resp),.auto_out_r_bits_echo_real_last(_axi4buf_auto_in_r_bits_echo_real_last),.auto_out_r_bits_last(_axi4buf_auto_in_r_bits_last)); 
endmodule
 
module ResetSynchronizerShiftReg_w1_d3_i0 (
  input clock,
  input reset,
  input io_d,
  output io_q) ; 
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain(.clock(clock),.reset(reset),.io_d(io_d),.io_q(io_q)); 
endmodule
 
module TestHarness (
  input clock,
  input reset,
  output io_success) ; 
   wire _SimDTM_debug_req_valid ;  
   wire [6:0] _SimDTM_debug_req_bits_addr ;  
   wire [31:0] _SimDTM_debug_req_bits_data ;  
   wire [1:0] _SimDTM_debug_req_bits_op ;  
   wire _SimDTM_debug_resp_ready ;  
   wire [31:0] _SimDTM_exit ;  
   wire _gated_clock_debug_clock_gate_out ;  
   wire _dmactiveAck_dmactiveAck_io_q ;  
   wire _debug_reset_syncd_debug_reset_sync_io_q ;  
   wire _mmio_mem_io_axi4_0_aw_ready ;  
   wire _mmio_mem_io_axi4_0_w_ready ;  
   wire _mmio_mem_io_axi4_0_b_valid ;  
   wire [3:0] _mmio_mem_io_axi4_0_b_bits_id ;  
   wire [1:0] _mmio_mem_io_axi4_0_b_bits_resp ;  
   wire _mmio_mem_io_axi4_0_ar_ready ;  
   wire _mmio_mem_io_axi4_0_r_valid ;  
   wire [3:0] _mmio_mem_io_axi4_0_r_bits_id ;  
   wire [63:0] _mmio_mem_io_axi4_0_r_bits_data ;  
   wire [1:0] _mmio_mem_io_axi4_0_r_bits_resp ;  
   wire _mmio_mem_io_axi4_0_r_bits_last ;  
   wire _mem_io_axi4_0_aw_ready ;  
   wire _mem_io_axi4_0_w_ready ;  
   wire _mem_io_axi4_0_b_valid ;  
   wire [3:0] _mem_io_axi4_0_b_bits_id ;  
   wire [1:0] _mem_io_axi4_0_b_bits_resp ;  
   wire _mem_io_axi4_0_ar_ready ;  
   wire _mem_io_axi4_0_r_valid ;  
   wire [3:0] _mem_io_axi4_0_r_bits_id ;  
   wire [63:0] _mem_io_axi4_0_r_bits_data ;  
   wire [1:0] _mem_io_axi4_0_r_bits_resp ;  
   wire _mem_io_axi4_0_r_bits_last ;  
   wire _ldut_reset_reg_io_q ;  
   wire _ldut_debug_clockeddmi_dmi_req_ready ;  
   wire _ldut_debug_clockeddmi_dmi_resp_valid ;  
   wire [31:0] _ldut_debug_clockeddmi_dmi_resp_bits_data ;  
   wire [1:0] _ldut_debug_clockeddmi_dmi_resp_bits_resp ;  
   wire _ldut_debug_ndreset ;  
   wire _ldut_debug_dmactive ;  
   wire _ldut_mem_axi4_0_aw_valid ;  
   wire [3:0] _ldut_mem_axi4_0_aw_bits_id ;  
   wire [31:0] _ldut_mem_axi4_0_aw_bits_addr ;  
   wire [7:0] _ldut_mem_axi4_0_aw_bits_len ;  
   wire [2:0] _ldut_mem_axi4_0_aw_bits_size ;  
   wire [1:0] _ldut_mem_axi4_0_aw_bits_burst ;  
   wire _ldut_mem_axi4_0_w_valid ;  
   wire [63:0] _ldut_mem_axi4_0_w_bits_data ;  
   wire [7:0] _ldut_mem_axi4_0_w_bits_strb ;  
   wire _ldut_mem_axi4_0_w_bits_last ;  
   wire _ldut_mem_axi4_0_b_ready ;  
   wire _ldut_mem_axi4_0_ar_valid ;  
   wire [3:0] _ldut_mem_axi4_0_ar_bits_id ;  
   wire [31:0] _ldut_mem_axi4_0_ar_bits_addr ;  
   wire [7:0] _ldut_mem_axi4_0_ar_bits_len ;  
   wire [2:0] _ldut_mem_axi4_0_ar_bits_size ;  
   wire [1:0] _ldut_mem_axi4_0_ar_bits_burst ;  
   wire _ldut_mem_axi4_0_r_ready ;  
   wire _ldut_mmio_axi4_0_aw_valid ;  
   wire [3:0] _ldut_mmio_axi4_0_aw_bits_id ;  
   wire [30:0] _ldut_mmio_axi4_0_aw_bits_addr ;  
   wire [7:0] _ldut_mmio_axi4_0_aw_bits_len ;  
   wire [2:0] _ldut_mmio_axi4_0_aw_bits_size ;  
   wire [1:0] _ldut_mmio_axi4_0_aw_bits_burst ;  
   wire _ldut_mmio_axi4_0_w_valid ;  
   wire [63:0] _ldut_mmio_axi4_0_w_bits_data ;  
   wire [7:0] _ldut_mmio_axi4_0_w_bits_strb ;  
   wire _ldut_mmio_axi4_0_w_bits_last ;  
   wire _ldut_mmio_axi4_0_b_ready ;  
   wire _ldut_mmio_axi4_0_ar_valid ;  
   wire [3:0] _ldut_mmio_axi4_0_ar_bits_id ;  
   wire [30:0] _ldut_mmio_axi4_0_ar_bits_addr ;  
   wire [7:0] _ldut_mmio_axi4_0_ar_bits_len ;  
   wire [2:0] _ldut_mmio_axi4_0_ar_bits_size ;  
   wire [1:0] _ldut_mmio_axi4_0_ar_bits_burst ;  
   wire _ldut_mmio_axi4_0_r_ready ;  
   wire debug_reset=~_debug_reset_syncd_debug_reset_sync_io_q ;  
   reg clock_en ;  
  always @( posedge clock)
       begin 
         if (~reset&(|(_SimDTM_exit[31:1])))
            begin 
              if (1)$display("Assertion failed: *** FAILED *** (exit code = %d)\n\n    at Periphery.scala:200 assert(io.exit < 2.U, \"*** FAILED *** (exit code = %%%%d)\\n\", io.exit >> 1.U)\n",{1'h0,_SimDTM_exit[31:1]});
              if (1)$display("");
            end 
       end
  
  always @(  posedge clock or  posedge debug_reset)
       begin 
         if (debug_reset)
            clock_en <=1'h1;
          else 
            clock_en <=_dmactiveAck_dmactiveAck_io_q;
       end
  initial
    begin #1ns;$readmemh("./hello_64bits.hex",TestHarness.mem.srams.mem_ext.Memory);
    end  initial
    begin #100ns;wait(TestHarness.ldut.mmio_axi4_0_aw_ready&TestHarness.ldut.mmio_axi4_0_aw_valid);wait(TestHarness.ldut.mmio_axi4_0_aw_bits_addr[30:0]==31'h7070_7070);wait(TestHarness.ldut.mmio_axi4_0_w_ready&TestHarness.ldut.mmio_axi4_0_w_valid);wait(TestHarness.ldut.mmio_axi4_0_w_bits_data[31:0]==32'hdead_beef);$display("**************************************************");$display("**************************************************");$display("****** PAT NAME : helloworld, PASS SUCCESSED********");$display("**************************************************");$display("**************************************************");
    end  
  ExampleRocketSystem ldut(.clock(clock),.reset(reset|_ldut_reset_reg_io_q),.resetctrl_hartIsInReset_0(reset),.debug_clock(_gated_clock_debug_clock_gate_out),.debug_reset(debug_reset),.debug_clockeddmi_dmi_req_ready(_ldut_debug_clockeddmi_dmi_req_ready),.debug_clockeddmi_dmi_req_valid(_SimDTM_debug_req_valid),.debug_clockeddmi_dmi_req_bits_addr(_SimDTM_debug_req_bits_addr),.debug_clockeddmi_dmi_req_bits_data(_SimDTM_debug_req_bits_data),.debug_clockeddmi_dmi_req_bits_op(_SimDTM_debug_req_bits_op),.debug_clockeddmi_dmi_resp_ready(_SimDTM_debug_resp_ready),.debug_clockeddmi_dmi_resp_valid(_ldut_debug_clockeddmi_dmi_resp_valid),.debug_clockeddmi_dmi_resp_bits_data(_ldut_debug_clockeddmi_dmi_resp_bits_data),.debug_clockeddmi_dmi_resp_bits_resp(_ldut_debug_clockeddmi_dmi_resp_bits_resp),.debug_clockeddmi_dmiClock(clock),.debug_clockeddmi_dmiReset(reset),.debug_ndreset(_ldut_debug_ndreset),.debug_dmactive(_ldut_debug_dmactive),.debug_dmactiveAck(_dmactiveAck_dmactiveAck_io_q),.mem_axi4_0_aw_ready(_mem_io_axi4_0_aw_ready),.mem_axi4_0_aw_valid(_ldut_mem_axi4_0_aw_valid),.mem_axi4_0_aw_bits_id(_ldut_mem_axi4_0_aw_bits_id),.mem_axi4_0_aw_bits_addr(_ldut_mem_axi4_0_aw_bits_addr),.mem_axi4_0_aw_bits_len(_ldut_mem_axi4_0_aw_bits_len),.mem_axi4_0_aw_bits_size(_ldut_mem_axi4_0_aw_bits_size),.mem_axi4_0_aw_bits_burst(_ldut_mem_axi4_0_aw_bits_burst),.mem_axi4_0_aw_bits_lock(),.mem_axi4_0_aw_bits_cache(),.mem_axi4_0_aw_bits_prot(),.mem_axi4_0_aw_bits_qos(),.mem_axi4_0_w_ready(_mem_io_axi4_0_w_ready),.mem_axi4_0_w_valid(_ldut_mem_axi4_0_w_valid),.mem_axi4_0_w_bits_data(_ldut_mem_axi4_0_w_bits_data),.mem_axi4_0_w_bits_strb(_ldut_mem_axi4_0_w_bits_strb),.mem_axi4_0_w_bits_last(_ldut_mem_axi4_0_w_bits_last),.mem_axi4_0_b_ready(_ldut_mem_axi4_0_b_ready),.mem_axi4_0_b_valid(_mem_io_axi4_0_b_valid),.mem_axi4_0_b_bits_id(_mem_io_axi4_0_b_bits_id),.mem_axi4_0_b_bits_resp(_mem_io_axi4_0_b_bits_resp),.mem_axi4_0_ar_ready(_mem_io_axi4_0_ar_ready),.mem_axi4_0_ar_valid(_ldut_mem_axi4_0_ar_valid),.mem_axi4_0_ar_bits_id(_ldut_mem_axi4_0_ar_bits_id),.mem_axi4_0_ar_bits_addr(_ldut_mem_axi4_0_ar_bits_addr),.mem_axi4_0_ar_bits_len(_ldut_mem_axi4_0_ar_bits_len),.mem_axi4_0_ar_bits_size(_ldut_mem_axi4_0_ar_bits_size),.mem_axi4_0_ar_bits_burst(_ldut_mem_axi4_0_ar_bits_burst),.mem_axi4_0_ar_bits_lock(),.mem_axi4_0_ar_bits_cache(),.mem_axi4_0_ar_bits_prot(),.mem_axi4_0_ar_bits_qos(),.mem_axi4_0_r_ready(_ldut_mem_axi4_0_r_ready),.mem_axi4_0_r_valid(_mem_io_axi4_0_r_valid),.mem_axi4_0_r_bits_id(_mem_io_axi4_0_r_bits_id),.mem_axi4_0_r_bits_data(_mem_io_axi4_0_r_bits_data),.mem_axi4_0_r_bits_resp(_mem_io_axi4_0_r_bits_resp),.mem_axi4_0_r_bits_last(_mem_io_axi4_0_r_bits_last),.mmio_axi4_0_aw_ready(_mmio_mem_io_axi4_0_aw_ready),.mmio_axi4_0_aw_valid(_ldut_mmio_axi4_0_aw_valid),.mmio_axi4_0_aw_bits_id(_ldut_mmio_axi4_0_aw_bits_id),.mmio_axi4_0_aw_bits_addr(_ldut_mmio_axi4_0_aw_bits_addr),.mmio_axi4_0_aw_bits_len(_ldut_mmio_axi4_0_aw_bits_len),.mmio_axi4_0_aw_bits_size(_ldut_mmio_axi4_0_aw_bits_size),.mmio_axi4_0_aw_bits_burst(_ldut_mmio_axi4_0_aw_bits_burst),.mmio_axi4_0_aw_bits_lock(),.mmio_axi4_0_aw_bits_cache(),.mmio_axi4_0_aw_bits_prot(),.mmio_axi4_0_aw_bits_qos(),.mmio_axi4_0_w_ready(_mmio_mem_io_axi4_0_w_ready),.mmio_axi4_0_w_valid(_ldut_mmio_axi4_0_w_valid),.mmio_axi4_0_w_bits_data(_ldut_mmio_axi4_0_w_bits_data),.mmio_axi4_0_w_bits_strb(_ldut_mmio_axi4_0_w_bits_strb),.mmio_axi4_0_w_bits_last(_ldut_mmio_axi4_0_w_bits_last),.mmio_axi4_0_b_ready(_ldut_mmio_axi4_0_b_ready),.mmio_axi4_0_b_valid(_mmio_mem_io_axi4_0_b_valid),.mmio_axi4_0_b_bits_id(_mmio_mem_io_axi4_0_b_bits_id),.mmio_axi4_0_b_bits_resp(_mmio_mem_io_axi4_0_b_bits_resp),.mmio_axi4_0_ar_ready(_mmio_mem_io_axi4_0_ar_ready),.mmio_axi4_0_ar_valid(_ldut_mmio_axi4_0_ar_valid),.mmio_axi4_0_ar_bits_id(_ldut_mmio_axi4_0_ar_bits_id),.mmio_axi4_0_ar_bits_addr(_ldut_mmio_axi4_0_ar_bits_addr),.mmio_axi4_0_ar_bits_len(_ldut_mmio_axi4_0_ar_bits_len),.mmio_axi4_0_ar_bits_size(_ldut_mmio_axi4_0_ar_bits_size),.mmio_axi4_0_ar_bits_burst(_ldut_mmio_axi4_0_ar_bits_burst),.mmio_axi4_0_ar_bits_lock(),.mmio_axi4_0_ar_bits_cache(),.mmio_axi4_0_ar_bits_prot(),.mmio_axi4_0_ar_bits_qos(),.mmio_axi4_0_r_ready(_ldut_mmio_axi4_0_r_ready),.mmio_axi4_0_r_valid(_mmio_mem_io_axi4_0_r_valid),.mmio_axi4_0_r_bits_id(_mmio_mem_io_axi4_0_r_bits_id),.mmio_axi4_0_r_bits_data(_mmio_mem_io_axi4_0_r_bits_data),.mmio_axi4_0_r_bits_resp(_mmio_mem_io_axi4_0_r_bits_resp),.mmio_axi4_0_r_bits_last(_mmio_mem_io_axi4_0_r_bits_last),.l2_frontend_bus_axi4_0_aw_ready(),.l2_frontend_bus_axi4_0_aw_valid(1'h0),.l2_frontend_bus_axi4_0_aw_bits_id(8'h0),.l2_frontend_bus_axi4_0_aw_bits_addr(32'h0),.l2_frontend_bus_axi4_0_aw_bits_len(8'h0),.l2_frontend_bus_axi4_0_aw_bits_size(3'h0),.l2_frontend_bus_axi4_0_aw_bits_burst(2'h0),.l2_frontend_bus_axi4_0_aw_bits_lock(1'h0),.l2_frontend_bus_axi4_0_aw_bits_cache(4'h0),.l2_frontend_bus_axi4_0_aw_bits_prot(3'h0),.l2_frontend_bus_axi4_0_aw_bits_qos(4'h0),.l2_frontend_bus_axi4_0_w_ready(),.l2_frontend_bus_axi4_0_w_valid(1'h0),.l2_frontend_bus_axi4_0_w_bits_data(64'h0),.l2_frontend_bus_axi4_0_w_bits_strb(8'h0),.l2_frontend_bus_axi4_0_w_bits_last(1'h0),.l2_frontend_bus_axi4_0_b_ready(1'h0),.l2_frontend_bus_axi4_0_b_valid(),.l2_frontend_bus_axi4_0_b_bits_id(),.l2_frontend_bus_axi4_0_b_bits_resp(),.l2_frontend_bus_axi4_0_ar_ready(),.l2_frontend_bus_axi4_0_ar_valid(1'h0),.l2_frontend_bus_axi4_0_ar_bits_id(8'h0),.l2_frontend_bus_axi4_0_ar_bits_addr(32'h0),.l2_frontend_bus_axi4_0_ar_bits_len(8'h0),.l2_frontend_bus_axi4_0_ar_bits_size(3'h0),.l2_frontend_bus_axi4_0_ar_bits_burst(2'h0),.l2_frontend_bus_axi4_0_ar_bits_lock(1'h0),.l2_frontend_bus_axi4_0_ar_bits_cache(4'h0),.l2_frontend_bus_axi4_0_ar_bits_prot(3'h0),.l2_frontend_bus_axi4_0_ar_bits_qos(4'h0),.l2_frontend_bus_axi4_0_r_ready(1'h0),.l2_frontend_bus_axi4_0_r_valid(),.l2_frontend_bus_axi4_0_r_bits_id(),.l2_frontend_bus_axi4_0_r_bits_data(),.l2_frontend_bus_axi4_0_r_bits_resp(),.l2_frontend_bus_axi4_0_r_bits_last(),.interrupts(2'h0)); 
  AsyncResetRegVec_w1_i0 ldut_reset_reg(.clock(clock),.reset(reset),.io_d(_ldut_debug_ndreset),.io_q(_ldut_reset_reg_io_q)); 
  SimAXIMem mem(.clock(clock),.reset(reset),.io_axi4_0_aw_ready(_mem_io_axi4_0_aw_ready),.io_axi4_0_aw_valid(_ldut_mem_axi4_0_aw_valid),.io_axi4_0_aw_bits_id(_ldut_mem_axi4_0_aw_bits_id),.io_axi4_0_aw_bits_addr(_ldut_mem_axi4_0_aw_bits_addr),.io_axi4_0_aw_bits_len(_ldut_mem_axi4_0_aw_bits_len),.io_axi4_0_aw_bits_size(_ldut_mem_axi4_0_aw_bits_size),.io_axi4_0_aw_bits_burst(_ldut_mem_axi4_0_aw_bits_burst),.io_axi4_0_w_ready(_mem_io_axi4_0_w_ready),.io_axi4_0_w_valid(_ldut_mem_axi4_0_w_valid),.io_axi4_0_w_bits_data(_ldut_mem_axi4_0_w_bits_data),.io_axi4_0_w_bits_strb(_ldut_mem_axi4_0_w_bits_strb),.io_axi4_0_w_bits_last(_ldut_mem_axi4_0_w_bits_last),.io_axi4_0_b_ready(_ldut_mem_axi4_0_b_ready),.io_axi4_0_b_valid(_mem_io_axi4_0_b_valid),.io_axi4_0_b_bits_id(_mem_io_axi4_0_b_bits_id),.io_axi4_0_b_bits_resp(_mem_io_axi4_0_b_bits_resp),.io_axi4_0_ar_ready(_mem_io_axi4_0_ar_ready),.io_axi4_0_ar_valid(_ldut_mem_axi4_0_ar_valid),.io_axi4_0_ar_bits_id(_ldut_mem_axi4_0_ar_bits_id),.io_axi4_0_ar_bits_addr(_ldut_mem_axi4_0_ar_bits_addr),.io_axi4_0_ar_bits_len(_ldut_mem_axi4_0_ar_bits_len),.io_axi4_0_ar_bits_size(_ldut_mem_axi4_0_ar_bits_size),.io_axi4_0_ar_bits_burst(_ldut_mem_axi4_0_ar_bits_burst),.io_axi4_0_r_ready(_ldut_mem_axi4_0_r_ready),.io_axi4_0_r_valid(_mem_io_axi4_0_r_valid),.io_axi4_0_r_bits_id(_mem_io_axi4_0_r_bits_id),.io_axi4_0_r_bits_data(_mem_io_axi4_0_r_bits_data),.io_axi4_0_r_bits_resp(_mem_io_axi4_0_r_bits_resp),.io_axi4_0_r_bits_last(_mem_io_axi4_0_r_bits_last)); 
  SimAXIMem_1 mmio_mem(.clock(clock),.reset(reset),.io_axi4_0_aw_ready(_mmio_mem_io_axi4_0_aw_ready),.io_axi4_0_aw_valid(_ldut_mmio_axi4_0_aw_valid),.io_axi4_0_aw_bits_id(_ldut_mmio_axi4_0_aw_bits_id),.io_axi4_0_aw_bits_addr(_ldut_mmio_axi4_0_aw_bits_addr),.io_axi4_0_aw_bits_len(_ldut_mmio_axi4_0_aw_bits_len),.io_axi4_0_aw_bits_size(_ldut_mmio_axi4_0_aw_bits_size),.io_axi4_0_aw_bits_burst(_ldut_mmio_axi4_0_aw_bits_burst),.io_axi4_0_w_ready(_mmio_mem_io_axi4_0_w_ready),.io_axi4_0_w_valid(_ldut_mmio_axi4_0_w_valid),.io_axi4_0_w_bits_data(_ldut_mmio_axi4_0_w_bits_data),.io_axi4_0_w_bits_strb(_ldut_mmio_axi4_0_w_bits_strb),.io_axi4_0_w_bits_last(_ldut_mmio_axi4_0_w_bits_last),.io_axi4_0_b_ready(_ldut_mmio_axi4_0_b_ready),.io_axi4_0_b_valid(_mmio_mem_io_axi4_0_b_valid),.io_axi4_0_b_bits_id(_mmio_mem_io_axi4_0_b_bits_id),.io_axi4_0_b_bits_resp(_mmio_mem_io_axi4_0_b_bits_resp),.io_axi4_0_ar_ready(_mmio_mem_io_axi4_0_ar_ready),.io_axi4_0_ar_valid(_ldut_mmio_axi4_0_ar_valid),.io_axi4_0_ar_bits_id(_ldut_mmio_axi4_0_ar_bits_id),.io_axi4_0_ar_bits_addr(_ldut_mmio_axi4_0_ar_bits_addr),.io_axi4_0_ar_bits_len(_ldut_mmio_axi4_0_ar_bits_len),.io_axi4_0_ar_bits_size(_ldut_mmio_axi4_0_ar_bits_size),.io_axi4_0_ar_bits_burst(_ldut_mmio_axi4_0_ar_bits_burst),.io_axi4_0_r_ready(_ldut_mmio_axi4_0_r_ready),.io_axi4_0_r_valid(_mmio_mem_io_axi4_0_r_valid),.io_axi4_0_r_bits_id(_mmio_mem_io_axi4_0_r_bits_id),.io_axi4_0_r_bits_data(_mmio_mem_io_axi4_0_r_bits_data),.io_axi4_0_r_bits_resp(_mmio_mem_io_axi4_0_r_bits_resp),.io_axi4_0_r_bits_last(_mmio_mem_io_axi4_0_r_bits_last)); 
  AsyncResetSynchronizerShiftReg_w1_d3_i0 debug_reset_syncd_debug_reset_sync(.clock(clock),.reset(reset),.io_d(1'h1),.io_q(_debug_reset_syncd_debug_reset_sync_io_q)); 
  ResetSynchronizerShiftReg_w1_d3_i0 dmactiveAck_dmactiveAck(.clock(clock),.reset(debug_reset),.io_d(_ldut_debug_dmactive),.io_q(_dmactiveAck_dmactiveAck_io_q)); 
endmodule
 
module plusarg_reader #(
 parameter FORMAT ="borked=%d",
 parameter WIDTH =1,
 parameter[WIDTH-1:0] DEFAULT =0) (
  output [WIDTH-1:0] out) ; 
   reg [WIDTH-1:0] myplus ;  
  assign out=myplus; initial
    begin 
      if (!$value$plusargs(FORMAT,myplus))
         myplus =DEFAULT;
    end  
endmodule
 

























